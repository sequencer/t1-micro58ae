
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module T1(
  input          indexedLoadStorePort_aw_ready,
  output         indexedLoadStorePort_aw_valid,
  output [1:0]   indexedLoadStorePort_aw_bits_id,
  output [31:0]  indexedLoadStorePort_aw_bits_addr,
  output [7:0]   indexedLoadStorePort_aw_bits_len,
  output [2:0]   indexedLoadStorePort_aw_bits_size,
  output [1:0]   indexedLoadStorePort_aw_bits_burst,
  output         indexedLoadStorePort_aw_bits_lock,
  output [3:0]   indexedLoadStorePort_aw_bits_cache,
  output [2:0]   indexedLoadStorePort_aw_bits_prot,
  output [3:0]   indexedLoadStorePort_aw_bits_qos,
                 indexedLoadStorePort_aw_bits_region,
  input          indexedLoadStorePort_w_ready,
  output         indexedLoadStorePort_w_valid,
  output [31:0]  indexedLoadStorePort_w_bits_data,
  output [3:0]   indexedLoadStorePort_w_bits_strb,
  output         indexedLoadStorePort_w_bits_last,
                 indexedLoadStorePort_b_ready,
  input          indexedLoadStorePort_b_valid,
  input  [1:0]   indexedLoadStorePort_b_bits_id,
                 indexedLoadStorePort_b_bits_resp,
  input          indexedLoadStorePort_ar_ready,
  output         indexedLoadStorePort_ar_valid,
  output [1:0]   indexedLoadStorePort_ar_bits_id,
  output [31:0]  indexedLoadStorePort_ar_bits_addr,
  output [7:0]   indexedLoadStorePort_ar_bits_len,
  output [2:0]   indexedLoadStorePort_ar_bits_size,
  output [1:0]   indexedLoadStorePort_ar_bits_burst,
  output         indexedLoadStorePort_ar_bits_lock,
  output [3:0]   indexedLoadStorePort_ar_bits_cache,
  output [2:0]   indexedLoadStorePort_ar_bits_prot,
  output [3:0]   indexedLoadStorePort_ar_bits_qos,
                 indexedLoadStorePort_ar_bits_region,
  output         indexedLoadStorePort_r_ready,
  input          indexedLoadStorePort_r_valid,
  input  [1:0]   indexedLoadStorePort_r_bits_id,
  input  [31:0]  indexedLoadStorePort_r_bits_data,
  input  [1:0]   indexedLoadStorePort_r_bits_resp,
  input          indexedLoadStorePort_r_bits_last,
                 highBandwidthLoadStorePort_aw_ready,
  output         highBandwidthLoadStorePort_aw_valid,
  output [1:0]   highBandwidthLoadStorePort_aw_bits_id,
  output [31:0]  highBandwidthLoadStorePort_aw_bits_addr,
  output [7:0]   highBandwidthLoadStorePort_aw_bits_len,
  output [2:0]   highBandwidthLoadStorePort_aw_bits_size,
  output [1:0]   highBandwidthLoadStorePort_aw_bits_burst,
  output         highBandwidthLoadStorePort_aw_bits_lock,
  output [3:0]   highBandwidthLoadStorePort_aw_bits_cache,
  output [2:0]   highBandwidthLoadStorePort_aw_bits_prot,
  output [3:0]   highBandwidthLoadStorePort_aw_bits_qos,
                 highBandwidthLoadStorePort_aw_bits_region,
  input          highBandwidthLoadStorePort_w_ready,
  output         highBandwidthLoadStorePort_w_valid,
  output [511:0] highBandwidthLoadStorePort_w_bits_data,
  output [63:0]  highBandwidthLoadStorePort_w_bits_strb,
  output         highBandwidthLoadStorePort_w_bits_last,
                 highBandwidthLoadStorePort_b_ready,
  input          highBandwidthLoadStorePort_b_valid,
  input  [1:0]   highBandwidthLoadStorePort_b_bits_id,
                 highBandwidthLoadStorePort_b_bits_resp,
  input          highBandwidthLoadStorePort_ar_ready,
  output         highBandwidthLoadStorePort_ar_valid,
  output [1:0]   highBandwidthLoadStorePort_ar_bits_id,
  output [31:0]  highBandwidthLoadStorePort_ar_bits_addr,
  output [7:0]   highBandwidthLoadStorePort_ar_bits_len,
  output [2:0]   highBandwidthLoadStorePort_ar_bits_size,
  output [1:0]   highBandwidthLoadStorePort_ar_bits_burst,
  output         highBandwidthLoadStorePort_ar_bits_lock,
  output [3:0]   highBandwidthLoadStorePort_ar_bits_cache,
  output [2:0]   highBandwidthLoadStorePort_ar_bits_prot,
  output [3:0]   highBandwidthLoadStorePort_ar_bits_qos,
                 highBandwidthLoadStorePort_ar_bits_region,
  output         highBandwidthLoadStorePort_r_ready,
  input          highBandwidthLoadStorePort_r_valid,
  input  [1:0]   highBandwidthLoadStorePort_r_bits_id,
  input  [511:0] highBandwidthLoadStorePort_r_bits_data,
  input  [1:0]   highBandwidthLoadStorePort_r_bits_resp,
  input          highBandwidthLoadStorePort_r_bits_last,
  output         retire_rd_valid,
  output [4:0]   retire_rd_bits_rdAddress,
  output [31:0]  retire_rd_bits_rdData,
  output         retire_rd_bits_isFp,
                 retire_csr_valid,
  output [31:0]  retire_csr_bits_vxsat,
                 retire_csr_bits_fflag,
  output         retire_mem_valid,
                 issue_ready,
  input          issue_valid,
  input  [31:0]  issue_bits_instruction,
                 issue_bits_rs1Data,
                 issue_bits_rs2Data,
                 issue_bits_vtype,
                 issue_bits_vl,
                 issue_bits_vstart,
                 issue_bits_vcsr,
  input          reset,
                 clock
);

  wire         _sinkVec_queue_fifo_63_empty;
  wire         _sinkVec_queue_fifo_63_full;
  wire         _sinkVec_queue_fifo_63_error;
  wire [46:0]  _sinkVec_queue_fifo_63_data_out;
  wire         _sinkVec_queue_fifo_62_empty;
  wire         _sinkVec_queue_fifo_62_full;
  wire         _sinkVec_queue_fifo_62_error;
  wire [46:0]  _sinkVec_queue_fifo_62_data_out;
  wire         _sinkVec_queue_fifo_61_empty;
  wire         _sinkVec_queue_fifo_61_full;
  wire         _sinkVec_queue_fifo_61_error;
  wire [11:0]  _sinkVec_queue_fifo_61_data_out;
  wire         _sinkVec_queue_fifo_60_empty;
  wire         _sinkVec_queue_fifo_60_full;
  wire         _sinkVec_queue_fifo_60_error;
  wire [11:0]  _sinkVec_queue_fifo_60_data_out;
  wire         _laneVec_15_readBusPort_0_enqRelease;
  wire         _laneVec_15_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_15_readBusPort_0_deq_bits_data;
  wire         _laneVec_15_readBusPort_1_enqRelease;
  wire         _laneVec_15_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_15_readBusPort_1_deq_bits_data;
  wire         _laneVec_15_writeBusPort_0_enqRelease;
  wire         _laneVec_15_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_15_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_15_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_15_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_15_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_15_writeBusPort_1_enqRelease;
  wire         _laneVec_15_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_15_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_15_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_15_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_15_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_15_laneRequest_ready;
  wire         _laneVec_15_maskUnitRequest_valid;
  wire [31:0]  _laneVec_15_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_15_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_15_maskUnitRequest_bits_index;
  wire         _laneVec_15_maskUnitRequest_bits_ffo;
  wire         _laneVec_15_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_15_maskRequestToLSU;
  wire [31:0]  _laneVec_15_vrfReadDataChannel;
  wire [7:0]   _laneVec_15_instructionFinished;
  wire [7:0]   _laneVec_15_vxsatReport;
  wire         _laneVec_15_v0Update_valid;
  wire [31:0]  _laneVec_15_v0Update_bits_data;
  wire [1:0]   _laneVec_15_v0Update_bits_offset;
  wire [3:0]   _laneVec_15_v0Update_bits_mask;
  wire [5:0]   _laneVec_15_maskSelect;
  wire [1:0]   _laneVec_15_maskSelectSew;
  wire         _sinkVec_queue_fifo_59_empty;
  wire         _sinkVec_queue_fifo_59_full;
  wire         _sinkVec_queue_fifo_59_error;
  wire [46:0]  _sinkVec_queue_fifo_59_data_out;
  wire         _sinkVec_queue_fifo_58_empty;
  wire         _sinkVec_queue_fifo_58_full;
  wire         _sinkVec_queue_fifo_58_error;
  wire [46:0]  _sinkVec_queue_fifo_58_data_out;
  wire         _sinkVec_queue_fifo_57_empty;
  wire         _sinkVec_queue_fifo_57_full;
  wire         _sinkVec_queue_fifo_57_error;
  wire [11:0]  _sinkVec_queue_fifo_57_data_out;
  wire         _sinkVec_queue_fifo_56_empty;
  wire         _sinkVec_queue_fifo_56_full;
  wire         _sinkVec_queue_fifo_56_error;
  wire [11:0]  _sinkVec_queue_fifo_56_data_out;
  wire         _laneVec_14_readBusPort_0_enqRelease;
  wire         _laneVec_14_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_14_readBusPort_0_deq_bits_data;
  wire         _laneVec_14_readBusPort_1_enqRelease;
  wire         _laneVec_14_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_14_readBusPort_1_deq_bits_data;
  wire         _laneVec_14_writeBusPort_0_enqRelease;
  wire         _laneVec_14_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_14_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_14_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_14_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_14_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_14_writeBusPort_1_enqRelease;
  wire         _laneVec_14_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_14_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_14_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_14_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_14_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_14_laneRequest_ready;
  wire         _laneVec_14_maskUnitRequest_valid;
  wire [31:0]  _laneVec_14_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_14_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_14_maskUnitRequest_bits_index;
  wire         _laneVec_14_maskUnitRequest_bits_ffo;
  wire         _laneVec_14_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_14_maskRequestToLSU;
  wire [31:0]  _laneVec_14_vrfReadDataChannel;
  wire [7:0]   _laneVec_14_instructionFinished;
  wire [7:0]   _laneVec_14_vxsatReport;
  wire         _laneVec_14_v0Update_valid;
  wire [31:0]  _laneVec_14_v0Update_bits_data;
  wire [1:0]   _laneVec_14_v0Update_bits_offset;
  wire [3:0]   _laneVec_14_v0Update_bits_mask;
  wire [5:0]   _laneVec_14_maskSelect;
  wire [1:0]   _laneVec_14_maskSelectSew;
  wire         _sinkVec_queue_fifo_55_empty;
  wire         _sinkVec_queue_fifo_55_full;
  wire         _sinkVec_queue_fifo_55_error;
  wire [46:0]  _sinkVec_queue_fifo_55_data_out;
  wire         _sinkVec_queue_fifo_54_empty;
  wire         _sinkVec_queue_fifo_54_full;
  wire         _sinkVec_queue_fifo_54_error;
  wire [46:0]  _sinkVec_queue_fifo_54_data_out;
  wire         _sinkVec_queue_fifo_53_empty;
  wire         _sinkVec_queue_fifo_53_full;
  wire         _sinkVec_queue_fifo_53_error;
  wire [11:0]  _sinkVec_queue_fifo_53_data_out;
  wire         _sinkVec_queue_fifo_52_empty;
  wire         _sinkVec_queue_fifo_52_full;
  wire         _sinkVec_queue_fifo_52_error;
  wire [11:0]  _sinkVec_queue_fifo_52_data_out;
  wire         _laneVec_13_readBusPort_0_enqRelease;
  wire         _laneVec_13_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_13_readBusPort_0_deq_bits_data;
  wire         _laneVec_13_readBusPort_1_enqRelease;
  wire         _laneVec_13_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_13_readBusPort_1_deq_bits_data;
  wire         _laneVec_13_writeBusPort_0_enqRelease;
  wire         _laneVec_13_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_13_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_13_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_13_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_13_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_13_writeBusPort_1_enqRelease;
  wire         _laneVec_13_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_13_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_13_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_13_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_13_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_13_laneRequest_ready;
  wire         _laneVec_13_maskUnitRequest_valid;
  wire [31:0]  _laneVec_13_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_13_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_13_maskUnitRequest_bits_index;
  wire         _laneVec_13_maskUnitRequest_bits_ffo;
  wire         _laneVec_13_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_13_maskRequestToLSU;
  wire [31:0]  _laneVec_13_vrfReadDataChannel;
  wire [7:0]   _laneVec_13_instructionFinished;
  wire [7:0]   _laneVec_13_vxsatReport;
  wire         _laneVec_13_v0Update_valid;
  wire [31:0]  _laneVec_13_v0Update_bits_data;
  wire [1:0]   _laneVec_13_v0Update_bits_offset;
  wire [3:0]   _laneVec_13_v0Update_bits_mask;
  wire [5:0]   _laneVec_13_maskSelect;
  wire [1:0]   _laneVec_13_maskSelectSew;
  wire         _sinkVec_queue_fifo_51_empty;
  wire         _sinkVec_queue_fifo_51_full;
  wire         _sinkVec_queue_fifo_51_error;
  wire [46:0]  _sinkVec_queue_fifo_51_data_out;
  wire         _sinkVec_queue_fifo_50_empty;
  wire         _sinkVec_queue_fifo_50_full;
  wire         _sinkVec_queue_fifo_50_error;
  wire [46:0]  _sinkVec_queue_fifo_50_data_out;
  wire         _sinkVec_queue_fifo_49_empty;
  wire         _sinkVec_queue_fifo_49_full;
  wire         _sinkVec_queue_fifo_49_error;
  wire [11:0]  _sinkVec_queue_fifo_49_data_out;
  wire         _sinkVec_queue_fifo_48_empty;
  wire         _sinkVec_queue_fifo_48_full;
  wire         _sinkVec_queue_fifo_48_error;
  wire [11:0]  _sinkVec_queue_fifo_48_data_out;
  wire         _laneVec_12_readBusPort_0_enqRelease;
  wire         _laneVec_12_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_12_readBusPort_0_deq_bits_data;
  wire         _laneVec_12_readBusPort_1_enqRelease;
  wire         _laneVec_12_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_12_readBusPort_1_deq_bits_data;
  wire         _laneVec_12_writeBusPort_0_enqRelease;
  wire         _laneVec_12_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_12_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_12_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_12_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_12_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_12_writeBusPort_1_enqRelease;
  wire         _laneVec_12_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_12_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_12_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_12_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_12_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_12_laneRequest_ready;
  wire         _laneVec_12_maskUnitRequest_valid;
  wire [31:0]  _laneVec_12_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_12_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_12_maskUnitRequest_bits_index;
  wire         _laneVec_12_maskUnitRequest_bits_ffo;
  wire         _laneVec_12_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_12_maskRequestToLSU;
  wire [31:0]  _laneVec_12_vrfReadDataChannel;
  wire [7:0]   _laneVec_12_instructionFinished;
  wire [7:0]   _laneVec_12_vxsatReport;
  wire         _laneVec_12_v0Update_valid;
  wire [31:0]  _laneVec_12_v0Update_bits_data;
  wire [1:0]   _laneVec_12_v0Update_bits_offset;
  wire [3:0]   _laneVec_12_v0Update_bits_mask;
  wire [5:0]   _laneVec_12_maskSelect;
  wire [1:0]   _laneVec_12_maskSelectSew;
  wire         _sinkVec_queue_fifo_47_empty;
  wire         _sinkVec_queue_fifo_47_full;
  wire         _sinkVec_queue_fifo_47_error;
  wire [46:0]  _sinkVec_queue_fifo_47_data_out;
  wire         _sinkVec_queue_fifo_46_empty;
  wire         _sinkVec_queue_fifo_46_full;
  wire         _sinkVec_queue_fifo_46_error;
  wire [46:0]  _sinkVec_queue_fifo_46_data_out;
  wire         _sinkVec_queue_fifo_45_empty;
  wire         _sinkVec_queue_fifo_45_full;
  wire         _sinkVec_queue_fifo_45_error;
  wire [11:0]  _sinkVec_queue_fifo_45_data_out;
  wire         _sinkVec_queue_fifo_44_empty;
  wire         _sinkVec_queue_fifo_44_full;
  wire         _sinkVec_queue_fifo_44_error;
  wire [11:0]  _sinkVec_queue_fifo_44_data_out;
  wire         _laneVec_11_readBusPort_0_enqRelease;
  wire         _laneVec_11_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_11_readBusPort_0_deq_bits_data;
  wire         _laneVec_11_readBusPort_1_enqRelease;
  wire         _laneVec_11_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_11_readBusPort_1_deq_bits_data;
  wire         _laneVec_11_writeBusPort_0_enqRelease;
  wire         _laneVec_11_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_11_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_11_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_11_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_11_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_11_writeBusPort_1_enqRelease;
  wire         _laneVec_11_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_11_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_11_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_11_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_11_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_11_laneRequest_ready;
  wire         _laneVec_11_maskUnitRequest_valid;
  wire [31:0]  _laneVec_11_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_11_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_11_maskUnitRequest_bits_index;
  wire         _laneVec_11_maskUnitRequest_bits_ffo;
  wire         _laneVec_11_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_11_maskRequestToLSU;
  wire [31:0]  _laneVec_11_vrfReadDataChannel;
  wire [7:0]   _laneVec_11_instructionFinished;
  wire [7:0]   _laneVec_11_vxsatReport;
  wire         _laneVec_11_v0Update_valid;
  wire [31:0]  _laneVec_11_v0Update_bits_data;
  wire [1:0]   _laneVec_11_v0Update_bits_offset;
  wire [3:0]   _laneVec_11_v0Update_bits_mask;
  wire [5:0]   _laneVec_11_maskSelect;
  wire [1:0]   _laneVec_11_maskSelectSew;
  wire         _sinkVec_queue_fifo_43_empty;
  wire         _sinkVec_queue_fifo_43_full;
  wire         _sinkVec_queue_fifo_43_error;
  wire [46:0]  _sinkVec_queue_fifo_43_data_out;
  wire         _sinkVec_queue_fifo_42_empty;
  wire         _sinkVec_queue_fifo_42_full;
  wire         _sinkVec_queue_fifo_42_error;
  wire [46:0]  _sinkVec_queue_fifo_42_data_out;
  wire         _sinkVec_queue_fifo_41_empty;
  wire         _sinkVec_queue_fifo_41_full;
  wire         _sinkVec_queue_fifo_41_error;
  wire [11:0]  _sinkVec_queue_fifo_41_data_out;
  wire         _sinkVec_queue_fifo_40_empty;
  wire         _sinkVec_queue_fifo_40_full;
  wire         _sinkVec_queue_fifo_40_error;
  wire [11:0]  _sinkVec_queue_fifo_40_data_out;
  wire         _laneVec_10_readBusPort_0_enqRelease;
  wire         _laneVec_10_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_10_readBusPort_0_deq_bits_data;
  wire         _laneVec_10_readBusPort_1_enqRelease;
  wire         _laneVec_10_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_10_readBusPort_1_deq_bits_data;
  wire         _laneVec_10_writeBusPort_0_enqRelease;
  wire         _laneVec_10_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_10_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_10_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_10_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_10_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_10_writeBusPort_1_enqRelease;
  wire         _laneVec_10_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_10_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_10_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_10_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_10_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_10_laneRequest_ready;
  wire         _laneVec_10_maskUnitRequest_valid;
  wire [31:0]  _laneVec_10_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_10_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_10_maskUnitRequest_bits_index;
  wire         _laneVec_10_maskUnitRequest_bits_ffo;
  wire         _laneVec_10_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_10_maskRequestToLSU;
  wire [31:0]  _laneVec_10_vrfReadDataChannel;
  wire [7:0]   _laneVec_10_instructionFinished;
  wire [7:0]   _laneVec_10_vxsatReport;
  wire         _laneVec_10_v0Update_valid;
  wire [31:0]  _laneVec_10_v0Update_bits_data;
  wire [1:0]   _laneVec_10_v0Update_bits_offset;
  wire [3:0]   _laneVec_10_v0Update_bits_mask;
  wire [5:0]   _laneVec_10_maskSelect;
  wire [1:0]   _laneVec_10_maskSelectSew;
  wire         _sinkVec_queue_fifo_39_empty;
  wire         _sinkVec_queue_fifo_39_full;
  wire         _sinkVec_queue_fifo_39_error;
  wire [46:0]  _sinkVec_queue_fifo_39_data_out;
  wire         _sinkVec_queue_fifo_38_empty;
  wire         _sinkVec_queue_fifo_38_full;
  wire         _sinkVec_queue_fifo_38_error;
  wire [46:0]  _sinkVec_queue_fifo_38_data_out;
  wire         _sinkVec_queue_fifo_37_empty;
  wire         _sinkVec_queue_fifo_37_full;
  wire         _sinkVec_queue_fifo_37_error;
  wire [11:0]  _sinkVec_queue_fifo_37_data_out;
  wire         _sinkVec_queue_fifo_36_empty;
  wire         _sinkVec_queue_fifo_36_full;
  wire         _sinkVec_queue_fifo_36_error;
  wire [11:0]  _sinkVec_queue_fifo_36_data_out;
  wire         _laneVec_9_readBusPort_0_enqRelease;
  wire         _laneVec_9_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_9_readBusPort_0_deq_bits_data;
  wire         _laneVec_9_readBusPort_1_enqRelease;
  wire         _laneVec_9_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_9_readBusPort_1_deq_bits_data;
  wire         _laneVec_9_writeBusPort_0_enqRelease;
  wire         _laneVec_9_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_9_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_9_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_9_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_9_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_9_writeBusPort_1_enqRelease;
  wire         _laneVec_9_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_9_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_9_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_9_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_9_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_9_laneRequest_ready;
  wire         _laneVec_9_maskUnitRequest_valid;
  wire [31:0]  _laneVec_9_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_9_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_9_maskUnitRequest_bits_index;
  wire         _laneVec_9_maskUnitRequest_bits_ffo;
  wire         _laneVec_9_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_9_maskRequestToLSU;
  wire [31:0]  _laneVec_9_vrfReadDataChannel;
  wire [7:0]   _laneVec_9_instructionFinished;
  wire [7:0]   _laneVec_9_vxsatReport;
  wire         _laneVec_9_v0Update_valid;
  wire [31:0]  _laneVec_9_v0Update_bits_data;
  wire [1:0]   _laneVec_9_v0Update_bits_offset;
  wire [3:0]   _laneVec_9_v0Update_bits_mask;
  wire [5:0]   _laneVec_9_maskSelect;
  wire [1:0]   _laneVec_9_maskSelectSew;
  wire         _sinkVec_queue_fifo_35_empty;
  wire         _sinkVec_queue_fifo_35_full;
  wire         _sinkVec_queue_fifo_35_error;
  wire [46:0]  _sinkVec_queue_fifo_35_data_out;
  wire         _sinkVec_queue_fifo_34_empty;
  wire         _sinkVec_queue_fifo_34_full;
  wire         _sinkVec_queue_fifo_34_error;
  wire [46:0]  _sinkVec_queue_fifo_34_data_out;
  wire         _sinkVec_queue_fifo_33_empty;
  wire         _sinkVec_queue_fifo_33_full;
  wire         _sinkVec_queue_fifo_33_error;
  wire [11:0]  _sinkVec_queue_fifo_33_data_out;
  wire         _sinkVec_queue_fifo_32_empty;
  wire         _sinkVec_queue_fifo_32_full;
  wire         _sinkVec_queue_fifo_32_error;
  wire [11:0]  _sinkVec_queue_fifo_32_data_out;
  wire         _laneVec_8_readBusPort_0_enqRelease;
  wire         _laneVec_8_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_8_readBusPort_0_deq_bits_data;
  wire         _laneVec_8_readBusPort_1_enqRelease;
  wire         _laneVec_8_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_8_readBusPort_1_deq_bits_data;
  wire         _laneVec_8_writeBusPort_0_enqRelease;
  wire         _laneVec_8_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_8_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_8_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_8_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_8_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_8_writeBusPort_1_enqRelease;
  wire         _laneVec_8_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_8_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_8_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_8_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_8_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_8_laneRequest_ready;
  wire         _laneVec_8_maskUnitRequest_valid;
  wire [31:0]  _laneVec_8_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_8_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_8_maskUnitRequest_bits_index;
  wire         _laneVec_8_maskUnitRequest_bits_ffo;
  wire         _laneVec_8_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_8_maskRequestToLSU;
  wire [31:0]  _laneVec_8_vrfReadDataChannel;
  wire [7:0]   _laneVec_8_instructionFinished;
  wire [7:0]   _laneVec_8_vxsatReport;
  wire         _laneVec_8_v0Update_valid;
  wire [31:0]  _laneVec_8_v0Update_bits_data;
  wire [1:0]   _laneVec_8_v0Update_bits_offset;
  wire [3:0]   _laneVec_8_v0Update_bits_mask;
  wire [5:0]   _laneVec_8_maskSelect;
  wire [1:0]   _laneVec_8_maskSelectSew;
  wire         _sinkVec_queue_fifo_31_empty;
  wire         _sinkVec_queue_fifo_31_full;
  wire         _sinkVec_queue_fifo_31_error;
  wire [46:0]  _sinkVec_queue_fifo_31_data_out;
  wire         _sinkVec_queue_fifo_30_empty;
  wire         _sinkVec_queue_fifo_30_full;
  wire         _sinkVec_queue_fifo_30_error;
  wire [46:0]  _sinkVec_queue_fifo_30_data_out;
  wire         _sinkVec_queue_fifo_29_empty;
  wire         _sinkVec_queue_fifo_29_full;
  wire         _sinkVec_queue_fifo_29_error;
  wire [11:0]  _sinkVec_queue_fifo_29_data_out;
  wire         _sinkVec_queue_fifo_28_empty;
  wire         _sinkVec_queue_fifo_28_full;
  wire         _sinkVec_queue_fifo_28_error;
  wire [11:0]  _sinkVec_queue_fifo_28_data_out;
  wire         _laneVec_7_readBusPort_0_enqRelease;
  wire         _laneVec_7_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_7_readBusPort_0_deq_bits_data;
  wire         _laneVec_7_readBusPort_1_enqRelease;
  wire         _laneVec_7_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_7_readBusPort_1_deq_bits_data;
  wire         _laneVec_7_writeBusPort_0_enqRelease;
  wire         _laneVec_7_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_7_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_7_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_7_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_7_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_7_writeBusPort_1_enqRelease;
  wire         _laneVec_7_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_7_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_7_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_7_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_7_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_7_laneRequest_ready;
  wire         _laneVec_7_maskUnitRequest_valid;
  wire [31:0]  _laneVec_7_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_7_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_7_maskUnitRequest_bits_index;
  wire         _laneVec_7_maskUnitRequest_bits_ffo;
  wire         _laneVec_7_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_7_maskRequestToLSU;
  wire [31:0]  _laneVec_7_vrfReadDataChannel;
  wire [7:0]   _laneVec_7_instructionFinished;
  wire [7:0]   _laneVec_7_vxsatReport;
  wire         _laneVec_7_v0Update_valid;
  wire [31:0]  _laneVec_7_v0Update_bits_data;
  wire [1:0]   _laneVec_7_v0Update_bits_offset;
  wire [3:0]   _laneVec_7_v0Update_bits_mask;
  wire [5:0]   _laneVec_7_maskSelect;
  wire [1:0]   _laneVec_7_maskSelectSew;
  wire         _sinkVec_queue_fifo_27_empty;
  wire         _sinkVec_queue_fifo_27_full;
  wire         _sinkVec_queue_fifo_27_error;
  wire [46:0]  _sinkVec_queue_fifo_27_data_out;
  wire         _sinkVec_queue_fifo_26_empty;
  wire         _sinkVec_queue_fifo_26_full;
  wire         _sinkVec_queue_fifo_26_error;
  wire [46:0]  _sinkVec_queue_fifo_26_data_out;
  wire         _sinkVec_queue_fifo_25_empty;
  wire         _sinkVec_queue_fifo_25_full;
  wire         _sinkVec_queue_fifo_25_error;
  wire [11:0]  _sinkVec_queue_fifo_25_data_out;
  wire         _sinkVec_queue_fifo_24_empty;
  wire         _sinkVec_queue_fifo_24_full;
  wire         _sinkVec_queue_fifo_24_error;
  wire [11:0]  _sinkVec_queue_fifo_24_data_out;
  wire         _laneVec_6_readBusPort_0_enqRelease;
  wire         _laneVec_6_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_6_readBusPort_0_deq_bits_data;
  wire         _laneVec_6_readBusPort_1_enqRelease;
  wire         _laneVec_6_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_6_readBusPort_1_deq_bits_data;
  wire         _laneVec_6_writeBusPort_0_enqRelease;
  wire         _laneVec_6_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_6_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_6_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_6_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_6_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_6_writeBusPort_1_enqRelease;
  wire         _laneVec_6_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_6_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_6_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_6_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_6_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_6_laneRequest_ready;
  wire         _laneVec_6_maskUnitRequest_valid;
  wire [31:0]  _laneVec_6_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_6_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_6_maskUnitRequest_bits_index;
  wire         _laneVec_6_maskUnitRequest_bits_ffo;
  wire         _laneVec_6_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_6_maskRequestToLSU;
  wire [31:0]  _laneVec_6_vrfReadDataChannel;
  wire [7:0]   _laneVec_6_instructionFinished;
  wire [7:0]   _laneVec_6_vxsatReport;
  wire         _laneVec_6_v0Update_valid;
  wire [31:0]  _laneVec_6_v0Update_bits_data;
  wire [1:0]   _laneVec_6_v0Update_bits_offset;
  wire [3:0]   _laneVec_6_v0Update_bits_mask;
  wire [5:0]   _laneVec_6_maskSelect;
  wire [1:0]   _laneVec_6_maskSelectSew;
  wire         _sinkVec_queue_fifo_23_empty;
  wire         _sinkVec_queue_fifo_23_full;
  wire         _sinkVec_queue_fifo_23_error;
  wire [46:0]  _sinkVec_queue_fifo_23_data_out;
  wire         _sinkVec_queue_fifo_22_empty;
  wire         _sinkVec_queue_fifo_22_full;
  wire         _sinkVec_queue_fifo_22_error;
  wire [46:0]  _sinkVec_queue_fifo_22_data_out;
  wire         _sinkVec_queue_fifo_21_empty;
  wire         _sinkVec_queue_fifo_21_full;
  wire         _sinkVec_queue_fifo_21_error;
  wire [11:0]  _sinkVec_queue_fifo_21_data_out;
  wire         _sinkVec_queue_fifo_20_empty;
  wire         _sinkVec_queue_fifo_20_full;
  wire         _sinkVec_queue_fifo_20_error;
  wire [11:0]  _sinkVec_queue_fifo_20_data_out;
  wire         _laneVec_5_readBusPort_0_enqRelease;
  wire         _laneVec_5_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_5_readBusPort_0_deq_bits_data;
  wire         _laneVec_5_readBusPort_1_enqRelease;
  wire         _laneVec_5_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_5_readBusPort_1_deq_bits_data;
  wire         _laneVec_5_writeBusPort_0_enqRelease;
  wire         _laneVec_5_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_5_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_5_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_5_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_5_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_5_writeBusPort_1_enqRelease;
  wire         _laneVec_5_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_5_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_5_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_5_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_5_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_5_laneRequest_ready;
  wire         _laneVec_5_maskUnitRequest_valid;
  wire [31:0]  _laneVec_5_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_5_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_5_maskUnitRequest_bits_index;
  wire         _laneVec_5_maskUnitRequest_bits_ffo;
  wire         _laneVec_5_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_5_maskRequestToLSU;
  wire [31:0]  _laneVec_5_vrfReadDataChannel;
  wire [7:0]   _laneVec_5_instructionFinished;
  wire [7:0]   _laneVec_5_vxsatReport;
  wire         _laneVec_5_v0Update_valid;
  wire [31:0]  _laneVec_5_v0Update_bits_data;
  wire [1:0]   _laneVec_5_v0Update_bits_offset;
  wire [3:0]   _laneVec_5_v0Update_bits_mask;
  wire [5:0]   _laneVec_5_maskSelect;
  wire [1:0]   _laneVec_5_maskSelectSew;
  wire         _sinkVec_queue_fifo_19_empty;
  wire         _sinkVec_queue_fifo_19_full;
  wire         _sinkVec_queue_fifo_19_error;
  wire [46:0]  _sinkVec_queue_fifo_19_data_out;
  wire         _sinkVec_queue_fifo_18_empty;
  wire         _sinkVec_queue_fifo_18_full;
  wire         _sinkVec_queue_fifo_18_error;
  wire [46:0]  _sinkVec_queue_fifo_18_data_out;
  wire         _sinkVec_queue_fifo_17_empty;
  wire         _sinkVec_queue_fifo_17_full;
  wire         _sinkVec_queue_fifo_17_error;
  wire [11:0]  _sinkVec_queue_fifo_17_data_out;
  wire         _sinkVec_queue_fifo_16_empty;
  wire         _sinkVec_queue_fifo_16_full;
  wire         _sinkVec_queue_fifo_16_error;
  wire [11:0]  _sinkVec_queue_fifo_16_data_out;
  wire         _laneVec_4_readBusPort_0_enqRelease;
  wire         _laneVec_4_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_4_readBusPort_0_deq_bits_data;
  wire         _laneVec_4_readBusPort_1_enqRelease;
  wire         _laneVec_4_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_4_readBusPort_1_deq_bits_data;
  wire         _laneVec_4_writeBusPort_0_enqRelease;
  wire         _laneVec_4_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_4_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_4_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_4_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_4_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_4_writeBusPort_1_enqRelease;
  wire         _laneVec_4_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_4_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_4_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_4_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_4_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_4_laneRequest_ready;
  wire         _laneVec_4_maskUnitRequest_valid;
  wire [31:0]  _laneVec_4_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_4_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_4_maskUnitRequest_bits_index;
  wire         _laneVec_4_maskUnitRequest_bits_ffo;
  wire         _laneVec_4_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_4_maskRequestToLSU;
  wire [31:0]  _laneVec_4_vrfReadDataChannel;
  wire [7:0]   _laneVec_4_instructionFinished;
  wire [7:0]   _laneVec_4_vxsatReport;
  wire         _laneVec_4_v0Update_valid;
  wire [31:0]  _laneVec_4_v0Update_bits_data;
  wire [1:0]   _laneVec_4_v0Update_bits_offset;
  wire [3:0]   _laneVec_4_v0Update_bits_mask;
  wire [5:0]   _laneVec_4_maskSelect;
  wire [1:0]   _laneVec_4_maskSelectSew;
  wire         _sinkVec_queue_fifo_15_empty;
  wire         _sinkVec_queue_fifo_15_full;
  wire         _sinkVec_queue_fifo_15_error;
  wire [46:0]  _sinkVec_queue_fifo_15_data_out;
  wire         _sinkVec_queue_fifo_14_empty;
  wire         _sinkVec_queue_fifo_14_full;
  wire         _sinkVec_queue_fifo_14_error;
  wire [46:0]  _sinkVec_queue_fifo_14_data_out;
  wire         _sinkVec_queue_fifo_13_empty;
  wire         _sinkVec_queue_fifo_13_full;
  wire         _sinkVec_queue_fifo_13_error;
  wire [11:0]  _sinkVec_queue_fifo_13_data_out;
  wire         _sinkVec_queue_fifo_12_empty;
  wire         _sinkVec_queue_fifo_12_full;
  wire         _sinkVec_queue_fifo_12_error;
  wire [11:0]  _sinkVec_queue_fifo_12_data_out;
  wire         _laneVec_3_readBusPort_0_enqRelease;
  wire         _laneVec_3_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_3_readBusPort_0_deq_bits_data;
  wire         _laneVec_3_readBusPort_1_enqRelease;
  wire         _laneVec_3_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_3_readBusPort_1_deq_bits_data;
  wire         _laneVec_3_writeBusPort_0_enqRelease;
  wire         _laneVec_3_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_3_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_3_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_3_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_3_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_3_writeBusPort_1_enqRelease;
  wire         _laneVec_3_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_3_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_3_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_3_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_3_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_3_laneRequest_ready;
  wire         _laneVec_3_maskUnitRequest_valid;
  wire [31:0]  _laneVec_3_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_3_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_3_maskUnitRequest_bits_index;
  wire         _laneVec_3_maskUnitRequest_bits_ffo;
  wire         _laneVec_3_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_3_maskRequestToLSU;
  wire [31:0]  _laneVec_3_vrfReadDataChannel;
  wire [7:0]   _laneVec_3_instructionFinished;
  wire [7:0]   _laneVec_3_vxsatReport;
  wire         _laneVec_3_v0Update_valid;
  wire [31:0]  _laneVec_3_v0Update_bits_data;
  wire [1:0]   _laneVec_3_v0Update_bits_offset;
  wire [3:0]   _laneVec_3_v0Update_bits_mask;
  wire [5:0]   _laneVec_3_maskSelect;
  wire [1:0]   _laneVec_3_maskSelectSew;
  wire         _sinkVec_queue_fifo_11_empty;
  wire         _sinkVec_queue_fifo_11_full;
  wire         _sinkVec_queue_fifo_11_error;
  wire [46:0]  _sinkVec_queue_fifo_11_data_out;
  wire         _sinkVec_queue_fifo_10_empty;
  wire         _sinkVec_queue_fifo_10_full;
  wire         _sinkVec_queue_fifo_10_error;
  wire [46:0]  _sinkVec_queue_fifo_10_data_out;
  wire         _sinkVec_queue_fifo_9_empty;
  wire         _sinkVec_queue_fifo_9_full;
  wire         _sinkVec_queue_fifo_9_error;
  wire [11:0]  _sinkVec_queue_fifo_9_data_out;
  wire         _sinkVec_queue_fifo_8_empty;
  wire         _sinkVec_queue_fifo_8_full;
  wire         _sinkVec_queue_fifo_8_error;
  wire [11:0]  _sinkVec_queue_fifo_8_data_out;
  wire         _laneVec_2_readBusPort_0_enqRelease;
  wire         _laneVec_2_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_2_readBusPort_0_deq_bits_data;
  wire         _laneVec_2_readBusPort_1_enqRelease;
  wire         _laneVec_2_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_2_readBusPort_1_deq_bits_data;
  wire         _laneVec_2_writeBusPort_0_enqRelease;
  wire         _laneVec_2_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_2_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_2_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_2_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_2_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_2_writeBusPort_1_enqRelease;
  wire         _laneVec_2_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_2_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_2_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_2_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_2_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_2_laneRequest_ready;
  wire         _laneVec_2_maskUnitRequest_valid;
  wire [31:0]  _laneVec_2_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_2_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_2_maskUnitRequest_bits_index;
  wire         _laneVec_2_maskUnitRequest_bits_ffo;
  wire         _laneVec_2_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_2_maskRequestToLSU;
  wire [31:0]  _laneVec_2_vrfReadDataChannel;
  wire [7:0]   _laneVec_2_instructionFinished;
  wire [7:0]   _laneVec_2_vxsatReport;
  wire         _laneVec_2_v0Update_valid;
  wire [31:0]  _laneVec_2_v0Update_bits_data;
  wire [1:0]   _laneVec_2_v0Update_bits_offset;
  wire [3:0]   _laneVec_2_v0Update_bits_mask;
  wire [5:0]   _laneVec_2_maskSelect;
  wire [1:0]   _laneVec_2_maskSelectSew;
  wire         _sinkVec_queue_fifo_7_empty;
  wire         _sinkVec_queue_fifo_7_full;
  wire         _sinkVec_queue_fifo_7_error;
  wire [46:0]  _sinkVec_queue_fifo_7_data_out;
  wire         _sinkVec_queue_fifo_6_empty;
  wire         _sinkVec_queue_fifo_6_full;
  wire         _sinkVec_queue_fifo_6_error;
  wire [46:0]  _sinkVec_queue_fifo_6_data_out;
  wire         _sinkVec_queue_fifo_5_empty;
  wire         _sinkVec_queue_fifo_5_full;
  wire         _sinkVec_queue_fifo_5_error;
  wire [11:0]  _sinkVec_queue_fifo_5_data_out;
  wire         _sinkVec_queue_fifo_4_empty;
  wire         _sinkVec_queue_fifo_4_full;
  wire         _sinkVec_queue_fifo_4_error;
  wire [11:0]  _sinkVec_queue_fifo_4_data_out;
  wire         _laneVec_1_readBusPort_0_enqRelease;
  wire         _laneVec_1_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_1_readBusPort_0_deq_bits_data;
  wire         _laneVec_1_readBusPort_1_enqRelease;
  wire         _laneVec_1_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_1_readBusPort_1_deq_bits_data;
  wire         _laneVec_1_writeBusPort_0_enqRelease;
  wire         _laneVec_1_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_1_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_1_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_1_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_1_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_1_writeBusPort_1_enqRelease;
  wire         _laneVec_1_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_1_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_1_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_1_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_1_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_1_laneRequest_ready;
  wire         _laneVec_1_maskUnitRequest_valid;
  wire [31:0]  _laneVec_1_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_1_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_1_maskUnitRequest_bits_index;
  wire         _laneVec_1_maskUnitRequest_bits_ffo;
  wire         _laneVec_1_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_1_maskRequestToLSU;
  wire [31:0]  _laneVec_1_vrfReadDataChannel;
  wire [7:0]   _laneVec_1_instructionFinished;
  wire [7:0]   _laneVec_1_vxsatReport;
  wire         _laneVec_1_v0Update_valid;
  wire [31:0]  _laneVec_1_v0Update_bits_data;
  wire [1:0]   _laneVec_1_v0Update_bits_offset;
  wire [3:0]   _laneVec_1_v0Update_bits_mask;
  wire [5:0]   _laneVec_1_maskSelect;
  wire [1:0]   _laneVec_1_maskSelectSew;
  wire         _sinkVec_queue_fifo_3_empty;
  wire         _sinkVec_queue_fifo_3_full;
  wire         _sinkVec_queue_fifo_3_error;
  wire [46:0]  _sinkVec_queue_fifo_3_data_out;
  wire         _sinkVec_queue_fifo_2_empty;
  wire         _sinkVec_queue_fifo_2_full;
  wire         _sinkVec_queue_fifo_2_error;
  wire [46:0]  _sinkVec_queue_fifo_2_data_out;
  wire         _sinkVec_queue_fifo_1_empty;
  wire         _sinkVec_queue_fifo_1_full;
  wire         _sinkVec_queue_fifo_1_error;
  wire [11:0]  _sinkVec_queue_fifo_1_data_out;
  wire         _sinkVec_queue_fifo_empty;
  wire         _sinkVec_queue_fifo_full;
  wire         _sinkVec_queue_fifo_error;
  wire [11:0]  _sinkVec_queue_fifo_data_out;
  wire         _laneVec_0_readBusPort_0_enqRelease;
  wire         _laneVec_0_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_0_readBusPort_0_deq_bits_data;
  wire         _laneVec_0_readBusPort_1_enqRelease;
  wire         _laneVec_0_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_0_readBusPort_1_deq_bits_data;
  wire         _laneVec_0_writeBusPort_0_enqRelease;
  wire         _laneVec_0_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_0_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_0_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_0_writeBusPort_0_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_0_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_0_writeBusPort_1_enqRelease;
  wire         _laneVec_0_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_0_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_0_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_0_writeBusPort_1_deq_bits_instructionIndex;
  wire [5:0]   _laneVec_0_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_0_laneRequest_ready;
  wire         _laneVec_0_maskUnitRequest_valid;
  wire [31:0]  _laneVec_0_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_0_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_0_maskUnitRequest_bits_index;
  wire         _laneVec_0_maskUnitRequest_bits_ffo;
  wire         _laneVec_0_maskUnitRequest_bits_fpReduceValid;
  wire         _laneVec_0_maskRequestToLSU;
  wire [31:0]  _laneVec_0_vrfReadDataChannel;
  wire [7:0]   _laneVec_0_instructionFinished;
  wire [7:0]   _laneVec_0_vxsatReport;
  wire         _laneVec_0_v0Update_valid;
  wire [31:0]  _laneVec_0_v0Update_bits_data;
  wire [1:0]   _laneVec_0_v0Update_bits_offset;
  wire [3:0]   _laneVec_0_v0Update_bits_mask;
  wire [5:0]   _laneVec_0_maskSelect;
  wire [1:0]   _laneVec_0_maskSelectSew;
  wire         _queue_fifo_15_empty;
  wire         _queue_fifo_15_full;
  wire         _queue_fifo_15_error;
  wire [149:0] _queue_fifo_15_data_out;
  wire         _queue_fifo_14_empty;
  wire         _queue_fifo_14_full;
  wire         _queue_fifo_14_error;
  wire [149:0] _queue_fifo_14_data_out;
  wire         _queue_fifo_13_empty;
  wire         _queue_fifo_13_full;
  wire         _queue_fifo_13_error;
  wire [149:0] _queue_fifo_13_data_out;
  wire         _queue_fifo_12_empty;
  wire         _queue_fifo_12_full;
  wire         _queue_fifo_12_error;
  wire [149:0] _queue_fifo_12_data_out;
  wire         _queue_fifo_11_empty;
  wire         _queue_fifo_11_full;
  wire         _queue_fifo_11_error;
  wire [149:0] _queue_fifo_11_data_out;
  wire         _queue_fifo_10_empty;
  wire         _queue_fifo_10_full;
  wire         _queue_fifo_10_error;
  wire [149:0] _queue_fifo_10_data_out;
  wire         _queue_fifo_9_empty;
  wire         _queue_fifo_9_full;
  wire         _queue_fifo_9_error;
  wire [149:0] _queue_fifo_9_data_out;
  wire         _queue_fifo_8_empty;
  wire         _queue_fifo_8_full;
  wire         _queue_fifo_8_error;
  wire [149:0] _queue_fifo_8_data_out;
  wire         _queue_fifo_7_empty;
  wire         _queue_fifo_7_full;
  wire         _queue_fifo_7_error;
  wire [149:0] _queue_fifo_7_data_out;
  wire         _queue_fifo_6_empty;
  wire         _queue_fifo_6_full;
  wire         _queue_fifo_6_error;
  wire [149:0] _queue_fifo_6_data_out;
  wire         _queue_fifo_5_empty;
  wire         _queue_fifo_5_full;
  wire         _queue_fifo_5_error;
  wire [149:0] _queue_fifo_5_data_out;
  wire         _queue_fifo_4_empty;
  wire         _queue_fifo_4_full;
  wire         _queue_fifo_4_error;
  wire [149:0] _queue_fifo_4_data_out;
  wire         _queue_fifo_3_empty;
  wire         _queue_fifo_3_full;
  wire         _queue_fifo_3_error;
  wire [149:0] _queue_fifo_3_data_out;
  wire         _queue_fifo_2_empty;
  wire         _queue_fifo_2_full;
  wire         _queue_fifo_2_error;
  wire [149:0] _queue_fifo_2_data_out;
  wire         _queue_fifo_1_empty;
  wire         _queue_fifo_1_full;
  wire         _queue_fifo_1_error;
  wire [149:0] _queue_fifo_1_data_out;
  wire         _queue_fifo_empty;
  wire         _queue_fifo_full;
  wire         _queue_fifo_error;
  wire [149:0] _queue_fifo_data_out;
  wire         _tokenManager_issueAllow;
  wire [7:0]   _tokenManager_v0WriteValid;
  wire         _maskUnit_exeResp_0_valid;
  wire [3:0]   _maskUnit_exeResp_0_bits_mask;
  wire [2:0]   _maskUnit_exeResp_0_bits_instructionIndex;
  wire         _maskUnit_exeResp_1_valid;
  wire [3:0]   _maskUnit_exeResp_1_bits_mask;
  wire [2:0]   _maskUnit_exeResp_1_bits_instructionIndex;
  wire         _maskUnit_exeResp_2_valid;
  wire [3:0]   _maskUnit_exeResp_2_bits_mask;
  wire [2:0]   _maskUnit_exeResp_2_bits_instructionIndex;
  wire         _maskUnit_exeResp_3_valid;
  wire [3:0]   _maskUnit_exeResp_3_bits_mask;
  wire [2:0]   _maskUnit_exeResp_3_bits_instructionIndex;
  wire         _maskUnit_exeResp_4_valid;
  wire [3:0]   _maskUnit_exeResp_4_bits_mask;
  wire [2:0]   _maskUnit_exeResp_4_bits_instructionIndex;
  wire         _maskUnit_exeResp_5_valid;
  wire [3:0]   _maskUnit_exeResp_5_bits_mask;
  wire [2:0]   _maskUnit_exeResp_5_bits_instructionIndex;
  wire         _maskUnit_exeResp_6_valid;
  wire [3:0]   _maskUnit_exeResp_6_bits_mask;
  wire [2:0]   _maskUnit_exeResp_6_bits_instructionIndex;
  wire         _maskUnit_exeResp_7_valid;
  wire [3:0]   _maskUnit_exeResp_7_bits_mask;
  wire [2:0]   _maskUnit_exeResp_7_bits_instructionIndex;
  wire         _maskUnit_exeResp_8_valid;
  wire [3:0]   _maskUnit_exeResp_8_bits_mask;
  wire [2:0]   _maskUnit_exeResp_8_bits_instructionIndex;
  wire         _maskUnit_exeResp_9_valid;
  wire [3:0]   _maskUnit_exeResp_9_bits_mask;
  wire [2:0]   _maskUnit_exeResp_9_bits_instructionIndex;
  wire         _maskUnit_exeResp_10_valid;
  wire [3:0]   _maskUnit_exeResp_10_bits_mask;
  wire [2:0]   _maskUnit_exeResp_10_bits_instructionIndex;
  wire         _maskUnit_exeResp_11_valid;
  wire [3:0]   _maskUnit_exeResp_11_bits_mask;
  wire [2:0]   _maskUnit_exeResp_11_bits_instructionIndex;
  wire         _maskUnit_exeResp_12_valid;
  wire [3:0]   _maskUnit_exeResp_12_bits_mask;
  wire [2:0]   _maskUnit_exeResp_12_bits_instructionIndex;
  wire         _maskUnit_exeResp_13_valid;
  wire [3:0]   _maskUnit_exeResp_13_bits_mask;
  wire [2:0]   _maskUnit_exeResp_13_bits_instructionIndex;
  wire         _maskUnit_exeResp_14_valid;
  wire [3:0]   _maskUnit_exeResp_14_bits_mask;
  wire [2:0]   _maskUnit_exeResp_14_bits_instructionIndex;
  wire         _maskUnit_exeResp_15_valid;
  wire [3:0]   _maskUnit_exeResp_15_bits_mask;
  wire [2:0]   _maskUnit_exeResp_15_bits_instructionIndex;
  wire         _maskUnit_tokenIO_0_maskRequestRelease;
  wire         _maskUnit_tokenIO_1_maskRequestRelease;
  wire         _maskUnit_tokenIO_2_maskRequestRelease;
  wire         _maskUnit_tokenIO_3_maskRequestRelease;
  wire         _maskUnit_tokenIO_4_maskRequestRelease;
  wire         _maskUnit_tokenIO_5_maskRequestRelease;
  wire         _maskUnit_tokenIO_6_maskRequestRelease;
  wire         _maskUnit_tokenIO_7_maskRequestRelease;
  wire         _maskUnit_tokenIO_8_maskRequestRelease;
  wire         _maskUnit_tokenIO_9_maskRequestRelease;
  wire         _maskUnit_tokenIO_10_maskRequestRelease;
  wire         _maskUnit_tokenIO_11_maskRequestRelease;
  wire         _maskUnit_tokenIO_12_maskRequestRelease;
  wire         _maskUnit_tokenIO_13_maskRequestRelease;
  wire         _maskUnit_tokenIO_14_maskRequestRelease;
  wire         _maskUnit_tokenIO_15_maskRequestRelease;
  wire [7:0]   _maskUnit_lastReport;
  wire [31:0]  _maskUnit_laneMaskInput_0;
  wire [31:0]  _maskUnit_laneMaskInput_1;
  wire [31:0]  _maskUnit_laneMaskInput_2;
  wire [31:0]  _maskUnit_laneMaskInput_3;
  wire [31:0]  _maskUnit_laneMaskInput_4;
  wire [31:0]  _maskUnit_laneMaskInput_5;
  wire [31:0]  _maskUnit_laneMaskInput_6;
  wire [31:0]  _maskUnit_laneMaskInput_7;
  wire [31:0]  _maskUnit_laneMaskInput_8;
  wire [31:0]  _maskUnit_laneMaskInput_9;
  wire [31:0]  _maskUnit_laneMaskInput_10;
  wire [31:0]  _maskUnit_laneMaskInput_11;
  wire [31:0]  _maskUnit_laneMaskInput_12;
  wire [31:0]  _maskUnit_laneMaskInput_13;
  wire [31:0]  _maskUnit_laneMaskInput_14;
  wire [31:0]  _maskUnit_laneMaskInput_15;
  wire         _maskUnit_gatherData_valid;
  wire [31:0]  _maskUnit_gatherData_bits;
  wire         _decode_decodeResult_orderReduce;
  wire         _decode_decodeResult_floatMul;
  wire [1:0]   _decode_decodeResult_fpExecutionType;
  wire         _decode_decodeResult_float;
  wire         _decode_decodeResult_specialSlot;
  wire [4:0]   _decode_decodeResult_topUop;
  wire         _decode_decodeResult_popCount;
  wire         _decode_decodeResult_ffo;
  wire         _decode_decodeResult_average;
  wire         _decode_decodeResult_reverse;
  wire         _decode_decodeResult_dontNeedExecuteInLane;
  wire         _decode_decodeResult_scheduler;
  wire         _decode_decodeResult_sReadVD;
  wire         _decode_decodeResult_vtype;
  wire         _decode_decodeResult_sWrite;
  wire         _decode_decodeResult_crossRead;
  wire         _decode_decodeResult_crossWrite;
  wire         _decode_decodeResult_maskUnit;
  wire         _decode_decodeResult_special;
  wire         _decode_decodeResult_saturate;
  wire         _decode_decodeResult_vwmacc;
  wire         _decode_decodeResult_readOnly;
  wire         _decode_decodeResult_maskSource;
  wire         _decode_decodeResult_maskDestination;
  wire         _decode_decodeResult_maskLogic;
  wire [3:0]   _decode_decodeResult_uop;
  wire         _decode_decodeResult_iota;
  wire         _decode_decodeResult_mv;
  wire         _decode_decodeResult_extend;
  wire         _decode_decodeResult_unOrderWrite;
  wire         _decode_decodeResult_compress;
  wire         _decode_decodeResult_gather16;
  wire         _decode_decodeResult_gather;
  wire         _decode_decodeResult_slid;
  wire         _decode_decodeResult_targetRd;
  wire         _decode_decodeResult_widenReduce;
  wire         _decode_decodeResult_red;
  wire         _decode_decodeResult_nr;
  wire         _decode_decodeResult_itype;
  wire         _decode_decodeResult_unsigned1;
  wire         _decode_decodeResult_unsigned0;
  wire         _decode_decodeResult_other;
  wire         _decode_decodeResult_multiCycle;
  wire         _decode_decodeResult_divider;
  wire         _decode_decodeResult_multiplier;
  wire         _decode_decodeResult_shift;
  wire         _decode_decodeResult_adder;
  wire         _decode_decodeResult_logic;
  wire         _lsu_request_ready;
  wire         _lsu_vrfWritePort_0_valid;
  wire [4:0]   _lsu_vrfWritePort_0_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_0_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_0_bits_instructionIndex;
  wire         _lsu_vrfWritePort_1_valid;
  wire [4:0]   _lsu_vrfWritePort_1_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_1_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_1_bits_instructionIndex;
  wire         _lsu_vrfWritePort_2_valid;
  wire [4:0]   _lsu_vrfWritePort_2_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_2_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_2_bits_instructionIndex;
  wire         _lsu_vrfWritePort_3_valid;
  wire [4:0]   _lsu_vrfWritePort_3_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_3_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_3_bits_instructionIndex;
  wire         _lsu_vrfWritePort_4_valid;
  wire [4:0]   _lsu_vrfWritePort_4_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_4_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_4_bits_instructionIndex;
  wire         _lsu_vrfWritePort_5_valid;
  wire [4:0]   _lsu_vrfWritePort_5_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_5_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_5_bits_instructionIndex;
  wire         _lsu_vrfWritePort_6_valid;
  wire [4:0]   _lsu_vrfWritePort_6_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_6_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_6_bits_instructionIndex;
  wire         _lsu_vrfWritePort_7_valid;
  wire [4:0]   _lsu_vrfWritePort_7_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_7_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_7_bits_instructionIndex;
  wire         _lsu_vrfWritePort_8_valid;
  wire [4:0]   _lsu_vrfWritePort_8_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_8_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_8_bits_instructionIndex;
  wire         _lsu_vrfWritePort_9_valid;
  wire [4:0]   _lsu_vrfWritePort_9_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_9_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_9_bits_instructionIndex;
  wire         _lsu_vrfWritePort_10_valid;
  wire [4:0]   _lsu_vrfWritePort_10_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_10_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_10_bits_instructionIndex;
  wire         _lsu_vrfWritePort_11_valid;
  wire [4:0]   _lsu_vrfWritePort_11_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_11_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_11_bits_instructionIndex;
  wire         _lsu_vrfWritePort_12_valid;
  wire [4:0]   _lsu_vrfWritePort_12_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_12_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_12_bits_instructionIndex;
  wire         _lsu_vrfWritePort_13_valid;
  wire [4:0]   _lsu_vrfWritePort_13_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_13_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_13_bits_instructionIndex;
  wire         _lsu_vrfWritePort_14_valid;
  wire [4:0]   _lsu_vrfWritePort_14_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_14_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_14_bits_instructionIndex;
  wire         _lsu_vrfWritePort_15_valid;
  wire [4:0]   _lsu_vrfWritePort_15_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_15_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_15_bits_instructionIndex;
  wire [7:0]   _lsu_dataInWriteQueue_0;
  wire [7:0]   _lsu_dataInWriteQueue_1;
  wire [7:0]   _lsu_dataInWriteQueue_2;
  wire [7:0]   _lsu_dataInWriteQueue_3;
  wire [7:0]   _lsu_dataInWriteQueue_4;
  wire [7:0]   _lsu_dataInWriteQueue_5;
  wire [7:0]   _lsu_dataInWriteQueue_6;
  wire [7:0]   _lsu_dataInWriteQueue_7;
  wire [7:0]   _lsu_dataInWriteQueue_8;
  wire [7:0]   _lsu_dataInWriteQueue_9;
  wire [7:0]   _lsu_dataInWriteQueue_10;
  wire [7:0]   _lsu_dataInWriteQueue_11;
  wire [7:0]   _lsu_dataInWriteQueue_12;
  wire [7:0]   _lsu_dataInWriteQueue_13;
  wire [7:0]   _lsu_dataInWriteQueue_14;
  wire [7:0]   _lsu_dataInWriteQueue_15;
  wire [7:0]   _lsu_lastReport;
  wire [15:0]  _lsu_tokenIO_offsetGroupRelease;
  wire         sinkVec_queue_63_almostFull;
  wire         sinkVec_queue_63_almostEmpty;
  wire         sinkVec_queue_62_almostFull;
  wire         sinkVec_queue_62_almostEmpty;
  wire         sinkVec_queue_61_almostFull;
  wire         sinkVec_queue_61_almostEmpty;
  wire         sinkVec_queue_60_almostFull;
  wire         sinkVec_queue_60_almostEmpty;
  wire         sinkVec_queue_59_almostFull;
  wire         sinkVec_queue_59_almostEmpty;
  wire         sinkVec_queue_58_almostFull;
  wire         sinkVec_queue_58_almostEmpty;
  wire         sinkVec_queue_57_almostFull;
  wire         sinkVec_queue_57_almostEmpty;
  wire         sinkVec_queue_56_almostFull;
  wire         sinkVec_queue_56_almostEmpty;
  wire         sinkVec_queue_55_almostFull;
  wire         sinkVec_queue_55_almostEmpty;
  wire         sinkVec_queue_54_almostFull;
  wire         sinkVec_queue_54_almostEmpty;
  wire         sinkVec_queue_53_almostFull;
  wire         sinkVec_queue_53_almostEmpty;
  wire         sinkVec_queue_52_almostFull;
  wire         sinkVec_queue_52_almostEmpty;
  wire         sinkVec_queue_51_almostFull;
  wire         sinkVec_queue_51_almostEmpty;
  wire         sinkVec_queue_50_almostFull;
  wire         sinkVec_queue_50_almostEmpty;
  wire         sinkVec_queue_49_almostFull;
  wire         sinkVec_queue_49_almostEmpty;
  wire         sinkVec_queue_48_almostFull;
  wire         sinkVec_queue_48_almostEmpty;
  wire         sinkVec_queue_47_almostFull;
  wire         sinkVec_queue_47_almostEmpty;
  wire         sinkVec_queue_46_almostFull;
  wire         sinkVec_queue_46_almostEmpty;
  wire         sinkVec_queue_45_almostFull;
  wire         sinkVec_queue_45_almostEmpty;
  wire         sinkVec_queue_44_almostFull;
  wire         sinkVec_queue_44_almostEmpty;
  wire         sinkVec_queue_43_almostFull;
  wire         sinkVec_queue_43_almostEmpty;
  wire         sinkVec_queue_42_almostFull;
  wire         sinkVec_queue_42_almostEmpty;
  wire         sinkVec_queue_41_almostFull;
  wire         sinkVec_queue_41_almostEmpty;
  wire         sinkVec_queue_40_almostFull;
  wire         sinkVec_queue_40_almostEmpty;
  wire         sinkVec_queue_39_almostFull;
  wire         sinkVec_queue_39_almostEmpty;
  wire         sinkVec_queue_38_almostFull;
  wire         sinkVec_queue_38_almostEmpty;
  wire         sinkVec_queue_37_almostFull;
  wire         sinkVec_queue_37_almostEmpty;
  wire         sinkVec_queue_36_almostFull;
  wire         sinkVec_queue_36_almostEmpty;
  wire         sinkVec_queue_35_almostFull;
  wire         sinkVec_queue_35_almostEmpty;
  wire         sinkVec_queue_34_almostFull;
  wire         sinkVec_queue_34_almostEmpty;
  wire         sinkVec_queue_33_almostFull;
  wire         sinkVec_queue_33_almostEmpty;
  wire         sinkVec_queue_32_almostFull;
  wire         sinkVec_queue_32_almostEmpty;
  wire         sinkVec_queue_31_almostFull;
  wire         sinkVec_queue_31_almostEmpty;
  wire         sinkVec_queue_30_almostFull;
  wire         sinkVec_queue_30_almostEmpty;
  wire         sinkVec_queue_29_almostFull;
  wire         sinkVec_queue_29_almostEmpty;
  wire         sinkVec_queue_28_almostFull;
  wire         sinkVec_queue_28_almostEmpty;
  wire         sinkVec_queue_27_almostFull;
  wire         sinkVec_queue_27_almostEmpty;
  wire         sinkVec_queue_26_almostFull;
  wire         sinkVec_queue_26_almostEmpty;
  wire         sinkVec_queue_25_almostFull;
  wire         sinkVec_queue_25_almostEmpty;
  wire         sinkVec_queue_24_almostFull;
  wire         sinkVec_queue_24_almostEmpty;
  wire         sinkVec_queue_23_almostFull;
  wire         sinkVec_queue_23_almostEmpty;
  wire         sinkVec_queue_22_almostFull;
  wire         sinkVec_queue_22_almostEmpty;
  wire         sinkVec_queue_21_almostFull;
  wire         sinkVec_queue_21_almostEmpty;
  wire         sinkVec_queue_20_almostFull;
  wire         sinkVec_queue_20_almostEmpty;
  wire         sinkVec_queue_19_almostFull;
  wire         sinkVec_queue_19_almostEmpty;
  wire         sinkVec_queue_18_almostFull;
  wire         sinkVec_queue_18_almostEmpty;
  wire         sinkVec_queue_17_almostFull;
  wire         sinkVec_queue_17_almostEmpty;
  wire         sinkVec_queue_16_almostFull;
  wire         sinkVec_queue_16_almostEmpty;
  wire         sinkVec_queue_15_almostFull;
  wire         sinkVec_queue_15_almostEmpty;
  wire         sinkVec_queue_14_almostFull;
  wire         sinkVec_queue_14_almostEmpty;
  wire         sinkVec_queue_13_almostFull;
  wire         sinkVec_queue_13_almostEmpty;
  wire         sinkVec_queue_12_almostFull;
  wire         sinkVec_queue_12_almostEmpty;
  wire         sinkVec_queue_11_almostFull;
  wire         sinkVec_queue_11_almostEmpty;
  wire         sinkVec_queue_10_almostFull;
  wire         sinkVec_queue_10_almostEmpty;
  wire         sinkVec_queue_9_almostFull;
  wire         sinkVec_queue_9_almostEmpty;
  wire         sinkVec_queue_8_almostFull;
  wire         sinkVec_queue_8_almostEmpty;
  wire         sinkVec_queue_7_almostFull;
  wire         sinkVec_queue_7_almostEmpty;
  wire         sinkVec_queue_6_almostFull;
  wire         sinkVec_queue_6_almostEmpty;
  wire         sinkVec_queue_5_almostFull;
  wire         sinkVec_queue_5_almostEmpty;
  wire         sinkVec_queue_4_almostFull;
  wire         sinkVec_queue_4_almostEmpty;
  wire         sinkVec_queue_3_almostFull;
  wire         sinkVec_queue_3_almostEmpty;
  wire         sinkVec_queue_2_almostFull;
  wire         sinkVec_queue_2_almostEmpty;
  wire         sinkVec_queue_1_almostFull;
  wire         sinkVec_queue_1_almostEmpty;
  wire         sinkVec_queue_almostFull;
  wire         sinkVec_queue_almostEmpty;
  wire         queue_15_almostFull;
  wire         queue_15_almostEmpty;
  wire         queue_14_almostFull;
  wire         queue_14_almostEmpty;
  wire         queue_13_almostFull;
  wire         queue_13_almostEmpty;
  wire         queue_12_almostFull;
  wire         queue_12_almostEmpty;
  wire         queue_11_almostFull;
  wire         queue_11_almostEmpty;
  wire         queue_10_almostFull;
  wire         queue_10_almostEmpty;
  wire         queue_9_almostFull;
  wire         queue_9_almostEmpty;
  wire         queue_8_almostFull;
  wire         queue_8_almostEmpty;
  wire         queue_7_almostFull;
  wire         queue_7_almostEmpty;
  wire         queue_6_almostFull;
  wire         queue_6_almostEmpty;
  wire         queue_5_almostFull;
  wire         queue_5_almostEmpty;
  wire         queue_4_almostFull;
  wire         queue_4_almostEmpty;
  wire         queue_3_almostFull;
  wire         queue_3_almostEmpty;
  wire         queue_2_almostFull;
  wire         queue_2_almostEmpty;
  wire         queue_1_almostFull;
  wire         queue_1_almostEmpty;
  wire         queue_almostFull;
  wire         queue_almostEmpty;
  wire [31:0]  retire_rd_bits_rdData_0;
  wire         highBandwidthLoadStorePort_r_ready_0;
  wire [31:0]  highBandwidthLoadStorePort_ar_bits_addr_0;
  wire         highBandwidthLoadStorePort_ar_valid_0;
  wire [63:0]  highBandwidthLoadStorePort_w_bits_strb_0;
  wire [511:0] highBandwidthLoadStorePort_w_bits_data_0;
  wire         highBandwidthLoadStorePort_w_valid_0;
  wire [31:0]  highBandwidthLoadStorePort_aw_bits_addr_0;
  wire [1:0]   highBandwidthLoadStorePort_aw_bits_id_0;
  wire         highBandwidthLoadStorePort_aw_valid_0;
  wire         indexedLoadStorePort_r_ready_0;
  wire [31:0]  indexedLoadStorePort_ar_bits_addr_0;
  wire         indexedLoadStorePort_ar_valid_0;
  wire [3:0]   indexedLoadStorePort_w_bits_strb_0;
  wire [31:0]  indexedLoadStorePort_w_bits_data_0;
  wire         indexedLoadStorePort_w_valid_0;
  wire [2:0]   indexedLoadStorePort_aw_bits_size_0;
  wire [31:0]  indexedLoadStorePort_aw_bits_addr_0;
  wire [1:0]   indexedLoadStorePort_aw_bits_id_0;
  wire         indexedLoadStorePort_aw_valid_0;
  wire [2:0]   x22_15_1_bits_instructionIndex;
  wire         x22_15_1_bits_last;
  wire [31:0]  x22_15_1_bits_data;
  wire [3:0]   x22_15_1_bits_mask;
  wire [1:0]   x22_15_1_bits_offset;
  wire [4:0]   x22_15_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_63_bits_instructionIndex;
  wire         sinkVec_sinkWire_63_bits_last;
  wire [31:0]  sinkVec_sinkWire_63_bits_data;
  wire [3:0]   sinkVec_sinkWire_63_bits_mask;
  wire [1:0]   sinkVec_sinkWire_63_bits_offset;
  wire [4:0]   sinkVec_sinkWire_63_bits_vd;
  wire         sinkVec_sinkWire_63_valid;
  wire         sinkVec_sinkWire_63_ready;
  wire [2:0]   x22_15_0_bits_instructionIndex;
  wire [31:0]  x22_15_0_bits_data;
  wire [3:0]   x22_15_0_bits_mask;
  wire [1:0]   x22_15_0_bits_offset;
  wire [4:0]   x22_15_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_62_bits_instructionIndex;
  wire         sinkVec_sinkWire_62_bits_last;
  wire [31:0]  sinkVec_sinkWire_62_bits_data;
  wire [3:0]   sinkVec_sinkWire_62_bits_mask;
  wire [1:0]   sinkVec_sinkWire_62_bits_offset;
  wire [4:0]   sinkVec_sinkWire_62_bits_vd;
  wire         sinkVec_sinkWire_62_valid;
  wire         sinkVec_sinkWire_62_ready;
  wire [2:0]   x13_15_1_bits_instructionIndex;
  wire [1:0]   x13_15_1_bits_offset;
  wire [4:0]   x13_15_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_61_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_61_bits_offset;
  wire [1:0]   sinkVec_sinkWire_61_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_61_bits_vs;
  wire         sinkVec_sinkWire_61_valid;
  wire         sinkVec_sinkWire_61_ready;
  wire [2:0]   x13_15_0_bits_instructionIndex;
  wire [1:0]   x13_15_0_bits_offset;
  wire [4:0]   x13_15_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_60_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_60_bits_offset;
  wire [1:0]   sinkVec_sinkWire_60_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_60_bits_vs;
  wire         sinkVec_sinkWire_60_valid;
  wire         sinkVec_sinkWire_60_ready;
  wire [2:0]   x22_14_1_bits_instructionIndex;
  wire         x22_14_1_bits_last;
  wire [31:0]  x22_14_1_bits_data;
  wire [3:0]   x22_14_1_bits_mask;
  wire [1:0]   x22_14_1_bits_offset;
  wire [4:0]   x22_14_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_59_bits_instructionIndex;
  wire         sinkVec_sinkWire_59_bits_last;
  wire [31:0]  sinkVec_sinkWire_59_bits_data;
  wire [3:0]   sinkVec_sinkWire_59_bits_mask;
  wire [1:0]   sinkVec_sinkWire_59_bits_offset;
  wire [4:0]   sinkVec_sinkWire_59_bits_vd;
  wire         sinkVec_sinkWire_59_valid;
  wire         sinkVec_sinkWire_59_ready;
  wire [2:0]   x22_14_0_bits_instructionIndex;
  wire [31:0]  x22_14_0_bits_data;
  wire [3:0]   x22_14_0_bits_mask;
  wire [1:0]   x22_14_0_bits_offset;
  wire [4:0]   x22_14_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_58_bits_instructionIndex;
  wire         sinkVec_sinkWire_58_bits_last;
  wire [31:0]  sinkVec_sinkWire_58_bits_data;
  wire [3:0]   sinkVec_sinkWire_58_bits_mask;
  wire [1:0]   sinkVec_sinkWire_58_bits_offset;
  wire [4:0]   sinkVec_sinkWire_58_bits_vd;
  wire         sinkVec_sinkWire_58_valid;
  wire         sinkVec_sinkWire_58_ready;
  wire [2:0]   x13_14_1_bits_instructionIndex;
  wire [1:0]   x13_14_1_bits_offset;
  wire [4:0]   x13_14_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_57_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_57_bits_offset;
  wire [1:0]   sinkVec_sinkWire_57_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_57_bits_vs;
  wire         sinkVec_sinkWire_57_valid;
  wire         sinkVec_sinkWire_57_ready;
  wire [2:0]   x13_14_0_bits_instructionIndex;
  wire [1:0]   x13_14_0_bits_offset;
  wire [4:0]   x13_14_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_56_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_56_bits_offset;
  wire [1:0]   sinkVec_sinkWire_56_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_56_bits_vs;
  wire         sinkVec_sinkWire_56_valid;
  wire         sinkVec_sinkWire_56_ready;
  wire [2:0]   x22_13_1_bits_instructionIndex;
  wire         x22_13_1_bits_last;
  wire [31:0]  x22_13_1_bits_data;
  wire [3:0]   x22_13_1_bits_mask;
  wire [1:0]   x22_13_1_bits_offset;
  wire [4:0]   x22_13_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_55_bits_instructionIndex;
  wire         sinkVec_sinkWire_55_bits_last;
  wire [31:0]  sinkVec_sinkWire_55_bits_data;
  wire [3:0]   sinkVec_sinkWire_55_bits_mask;
  wire [1:0]   sinkVec_sinkWire_55_bits_offset;
  wire [4:0]   sinkVec_sinkWire_55_bits_vd;
  wire         sinkVec_sinkWire_55_valid;
  wire         sinkVec_sinkWire_55_ready;
  wire [2:0]   x22_13_0_bits_instructionIndex;
  wire [31:0]  x22_13_0_bits_data;
  wire [3:0]   x22_13_0_bits_mask;
  wire [1:0]   x22_13_0_bits_offset;
  wire [4:0]   x22_13_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_54_bits_instructionIndex;
  wire         sinkVec_sinkWire_54_bits_last;
  wire [31:0]  sinkVec_sinkWire_54_bits_data;
  wire [3:0]   sinkVec_sinkWire_54_bits_mask;
  wire [1:0]   sinkVec_sinkWire_54_bits_offset;
  wire [4:0]   sinkVec_sinkWire_54_bits_vd;
  wire         sinkVec_sinkWire_54_valid;
  wire         sinkVec_sinkWire_54_ready;
  wire [2:0]   x13_13_1_bits_instructionIndex;
  wire [1:0]   x13_13_1_bits_offset;
  wire [4:0]   x13_13_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_53_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_53_bits_offset;
  wire [1:0]   sinkVec_sinkWire_53_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_53_bits_vs;
  wire         sinkVec_sinkWire_53_valid;
  wire         sinkVec_sinkWire_53_ready;
  wire [2:0]   x13_13_0_bits_instructionIndex;
  wire [1:0]   x13_13_0_bits_offset;
  wire [4:0]   x13_13_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_52_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_52_bits_offset;
  wire [1:0]   sinkVec_sinkWire_52_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_52_bits_vs;
  wire         sinkVec_sinkWire_52_valid;
  wire         sinkVec_sinkWire_52_ready;
  wire [2:0]   x22_12_1_bits_instructionIndex;
  wire         x22_12_1_bits_last;
  wire [31:0]  x22_12_1_bits_data;
  wire [3:0]   x22_12_1_bits_mask;
  wire [1:0]   x22_12_1_bits_offset;
  wire [4:0]   x22_12_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_51_bits_instructionIndex;
  wire         sinkVec_sinkWire_51_bits_last;
  wire [31:0]  sinkVec_sinkWire_51_bits_data;
  wire [3:0]   sinkVec_sinkWire_51_bits_mask;
  wire [1:0]   sinkVec_sinkWire_51_bits_offset;
  wire [4:0]   sinkVec_sinkWire_51_bits_vd;
  wire         sinkVec_sinkWire_51_valid;
  wire         sinkVec_sinkWire_51_ready;
  wire [2:0]   x22_12_0_bits_instructionIndex;
  wire [31:0]  x22_12_0_bits_data;
  wire [3:0]   x22_12_0_bits_mask;
  wire [1:0]   x22_12_0_bits_offset;
  wire [4:0]   x22_12_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_50_bits_instructionIndex;
  wire         sinkVec_sinkWire_50_bits_last;
  wire [31:0]  sinkVec_sinkWire_50_bits_data;
  wire [3:0]   sinkVec_sinkWire_50_bits_mask;
  wire [1:0]   sinkVec_sinkWire_50_bits_offset;
  wire [4:0]   sinkVec_sinkWire_50_bits_vd;
  wire         sinkVec_sinkWire_50_valid;
  wire         sinkVec_sinkWire_50_ready;
  wire [2:0]   x13_12_1_bits_instructionIndex;
  wire [1:0]   x13_12_1_bits_offset;
  wire [4:0]   x13_12_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_49_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_49_bits_offset;
  wire [1:0]   sinkVec_sinkWire_49_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_49_bits_vs;
  wire         sinkVec_sinkWire_49_valid;
  wire         sinkVec_sinkWire_49_ready;
  wire [2:0]   x13_12_0_bits_instructionIndex;
  wire [1:0]   x13_12_0_bits_offset;
  wire [4:0]   x13_12_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_48_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_48_bits_offset;
  wire [1:0]   sinkVec_sinkWire_48_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_48_bits_vs;
  wire         sinkVec_sinkWire_48_valid;
  wire         sinkVec_sinkWire_48_ready;
  wire [2:0]   x22_11_1_bits_instructionIndex;
  wire         x22_11_1_bits_last;
  wire [31:0]  x22_11_1_bits_data;
  wire [3:0]   x22_11_1_bits_mask;
  wire [1:0]   x22_11_1_bits_offset;
  wire [4:0]   x22_11_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_47_bits_instructionIndex;
  wire         sinkVec_sinkWire_47_bits_last;
  wire [31:0]  sinkVec_sinkWire_47_bits_data;
  wire [3:0]   sinkVec_sinkWire_47_bits_mask;
  wire [1:0]   sinkVec_sinkWire_47_bits_offset;
  wire [4:0]   sinkVec_sinkWire_47_bits_vd;
  wire         sinkVec_sinkWire_47_valid;
  wire         sinkVec_sinkWire_47_ready;
  wire [2:0]   x22_11_0_bits_instructionIndex;
  wire [31:0]  x22_11_0_bits_data;
  wire [3:0]   x22_11_0_bits_mask;
  wire [1:0]   x22_11_0_bits_offset;
  wire [4:0]   x22_11_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_46_bits_instructionIndex;
  wire         sinkVec_sinkWire_46_bits_last;
  wire [31:0]  sinkVec_sinkWire_46_bits_data;
  wire [3:0]   sinkVec_sinkWire_46_bits_mask;
  wire [1:0]   sinkVec_sinkWire_46_bits_offset;
  wire [4:0]   sinkVec_sinkWire_46_bits_vd;
  wire         sinkVec_sinkWire_46_valid;
  wire         sinkVec_sinkWire_46_ready;
  wire [2:0]   x13_11_1_bits_instructionIndex;
  wire [1:0]   x13_11_1_bits_offset;
  wire [4:0]   x13_11_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_45_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_45_bits_offset;
  wire [1:0]   sinkVec_sinkWire_45_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_45_bits_vs;
  wire         sinkVec_sinkWire_45_valid;
  wire         sinkVec_sinkWire_45_ready;
  wire [2:0]   x13_11_0_bits_instructionIndex;
  wire [1:0]   x13_11_0_bits_offset;
  wire [4:0]   x13_11_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_44_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_44_bits_offset;
  wire [1:0]   sinkVec_sinkWire_44_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_44_bits_vs;
  wire         sinkVec_sinkWire_44_valid;
  wire         sinkVec_sinkWire_44_ready;
  wire [2:0]   x22_10_1_bits_instructionIndex;
  wire         x22_10_1_bits_last;
  wire [31:0]  x22_10_1_bits_data;
  wire [3:0]   x22_10_1_bits_mask;
  wire [1:0]   x22_10_1_bits_offset;
  wire [4:0]   x22_10_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_43_bits_instructionIndex;
  wire         sinkVec_sinkWire_43_bits_last;
  wire [31:0]  sinkVec_sinkWire_43_bits_data;
  wire [3:0]   sinkVec_sinkWire_43_bits_mask;
  wire [1:0]   sinkVec_sinkWire_43_bits_offset;
  wire [4:0]   sinkVec_sinkWire_43_bits_vd;
  wire         sinkVec_sinkWire_43_valid;
  wire         sinkVec_sinkWire_43_ready;
  wire [2:0]   x22_10_0_bits_instructionIndex;
  wire [31:0]  x22_10_0_bits_data;
  wire [3:0]   x22_10_0_bits_mask;
  wire [1:0]   x22_10_0_bits_offset;
  wire [4:0]   x22_10_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_42_bits_instructionIndex;
  wire         sinkVec_sinkWire_42_bits_last;
  wire [31:0]  sinkVec_sinkWire_42_bits_data;
  wire [3:0]   sinkVec_sinkWire_42_bits_mask;
  wire [1:0]   sinkVec_sinkWire_42_bits_offset;
  wire [4:0]   sinkVec_sinkWire_42_bits_vd;
  wire         sinkVec_sinkWire_42_valid;
  wire         sinkVec_sinkWire_42_ready;
  wire [2:0]   x13_10_1_bits_instructionIndex;
  wire [1:0]   x13_10_1_bits_offset;
  wire [4:0]   x13_10_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_41_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_41_bits_offset;
  wire [1:0]   sinkVec_sinkWire_41_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_41_bits_vs;
  wire         sinkVec_sinkWire_41_valid;
  wire         sinkVec_sinkWire_41_ready;
  wire [2:0]   x13_10_0_bits_instructionIndex;
  wire [1:0]   x13_10_0_bits_offset;
  wire [4:0]   x13_10_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_40_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_40_bits_offset;
  wire [1:0]   sinkVec_sinkWire_40_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_40_bits_vs;
  wire         sinkVec_sinkWire_40_valid;
  wire         sinkVec_sinkWire_40_ready;
  wire [2:0]   x22_9_1_bits_instructionIndex;
  wire         x22_9_1_bits_last;
  wire [31:0]  x22_9_1_bits_data;
  wire [3:0]   x22_9_1_bits_mask;
  wire [1:0]   x22_9_1_bits_offset;
  wire [4:0]   x22_9_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_39_bits_instructionIndex;
  wire         sinkVec_sinkWire_39_bits_last;
  wire [31:0]  sinkVec_sinkWire_39_bits_data;
  wire [3:0]   sinkVec_sinkWire_39_bits_mask;
  wire [1:0]   sinkVec_sinkWire_39_bits_offset;
  wire [4:0]   sinkVec_sinkWire_39_bits_vd;
  wire         sinkVec_sinkWire_39_valid;
  wire         sinkVec_sinkWire_39_ready;
  wire [2:0]   x22_9_0_bits_instructionIndex;
  wire [31:0]  x22_9_0_bits_data;
  wire [3:0]   x22_9_0_bits_mask;
  wire [1:0]   x22_9_0_bits_offset;
  wire [4:0]   x22_9_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_38_bits_instructionIndex;
  wire         sinkVec_sinkWire_38_bits_last;
  wire [31:0]  sinkVec_sinkWire_38_bits_data;
  wire [3:0]   sinkVec_sinkWire_38_bits_mask;
  wire [1:0]   sinkVec_sinkWire_38_bits_offset;
  wire [4:0]   sinkVec_sinkWire_38_bits_vd;
  wire         sinkVec_sinkWire_38_valid;
  wire         sinkVec_sinkWire_38_ready;
  wire [2:0]   x13_9_1_bits_instructionIndex;
  wire [1:0]   x13_9_1_bits_offset;
  wire [4:0]   x13_9_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_37_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_37_bits_offset;
  wire [1:0]   sinkVec_sinkWire_37_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_37_bits_vs;
  wire         sinkVec_sinkWire_37_valid;
  wire         sinkVec_sinkWire_37_ready;
  wire [2:0]   x13_9_0_bits_instructionIndex;
  wire [1:0]   x13_9_0_bits_offset;
  wire [4:0]   x13_9_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_36_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_36_bits_offset;
  wire [1:0]   sinkVec_sinkWire_36_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_36_bits_vs;
  wire         sinkVec_sinkWire_36_valid;
  wire         sinkVec_sinkWire_36_ready;
  wire [2:0]   x22_8_1_bits_instructionIndex;
  wire         x22_8_1_bits_last;
  wire [31:0]  x22_8_1_bits_data;
  wire [3:0]   x22_8_1_bits_mask;
  wire [1:0]   x22_8_1_bits_offset;
  wire [4:0]   x22_8_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_35_bits_instructionIndex;
  wire         sinkVec_sinkWire_35_bits_last;
  wire [31:0]  sinkVec_sinkWire_35_bits_data;
  wire [3:0]   sinkVec_sinkWire_35_bits_mask;
  wire [1:0]   sinkVec_sinkWire_35_bits_offset;
  wire [4:0]   sinkVec_sinkWire_35_bits_vd;
  wire         sinkVec_sinkWire_35_valid;
  wire         sinkVec_sinkWire_35_ready;
  wire [2:0]   x22_8_0_bits_instructionIndex;
  wire [31:0]  x22_8_0_bits_data;
  wire [3:0]   x22_8_0_bits_mask;
  wire [1:0]   x22_8_0_bits_offset;
  wire [4:0]   x22_8_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_34_bits_instructionIndex;
  wire         sinkVec_sinkWire_34_bits_last;
  wire [31:0]  sinkVec_sinkWire_34_bits_data;
  wire [3:0]   sinkVec_sinkWire_34_bits_mask;
  wire [1:0]   sinkVec_sinkWire_34_bits_offset;
  wire [4:0]   sinkVec_sinkWire_34_bits_vd;
  wire         sinkVec_sinkWire_34_valid;
  wire         sinkVec_sinkWire_34_ready;
  wire [2:0]   x13_8_1_bits_instructionIndex;
  wire [1:0]   x13_8_1_bits_offset;
  wire [4:0]   x13_8_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_33_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_33_bits_offset;
  wire [1:0]   sinkVec_sinkWire_33_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_33_bits_vs;
  wire         sinkVec_sinkWire_33_valid;
  wire         sinkVec_sinkWire_33_ready;
  wire [2:0]   x13_8_0_bits_instructionIndex;
  wire [1:0]   x13_8_0_bits_offset;
  wire [4:0]   x13_8_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_32_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_32_bits_offset;
  wire [1:0]   sinkVec_sinkWire_32_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_32_bits_vs;
  wire         sinkVec_sinkWire_32_valid;
  wire         sinkVec_sinkWire_32_ready;
  wire [2:0]   x22_7_1_bits_instructionIndex;
  wire         x22_7_1_bits_last;
  wire [31:0]  x22_7_1_bits_data;
  wire [3:0]   x22_7_1_bits_mask;
  wire [1:0]   x22_7_1_bits_offset;
  wire [4:0]   x22_7_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_31_bits_instructionIndex;
  wire         sinkVec_sinkWire_31_bits_last;
  wire [31:0]  sinkVec_sinkWire_31_bits_data;
  wire [3:0]   sinkVec_sinkWire_31_bits_mask;
  wire [1:0]   sinkVec_sinkWire_31_bits_offset;
  wire [4:0]   sinkVec_sinkWire_31_bits_vd;
  wire         sinkVec_sinkWire_31_valid;
  wire         sinkVec_sinkWire_31_ready;
  wire [2:0]   x22_7_0_bits_instructionIndex;
  wire [31:0]  x22_7_0_bits_data;
  wire [3:0]   x22_7_0_bits_mask;
  wire [1:0]   x22_7_0_bits_offset;
  wire [4:0]   x22_7_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_30_bits_instructionIndex;
  wire         sinkVec_sinkWire_30_bits_last;
  wire [31:0]  sinkVec_sinkWire_30_bits_data;
  wire [3:0]   sinkVec_sinkWire_30_bits_mask;
  wire [1:0]   sinkVec_sinkWire_30_bits_offset;
  wire [4:0]   sinkVec_sinkWire_30_bits_vd;
  wire         sinkVec_sinkWire_30_valid;
  wire         sinkVec_sinkWire_30_ready;
  wire [2:0]   x13_7_1_bits_instructionIndex;
  wire [1:0]   x13_7_1_bits_offset;
  wire [4:0]   x13_7_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_29_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_29_bits_offset;
  wire [1:0]   sinkVec_sinkWire_29_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_29_bits_vs;
  wire         sinkVec_sinkWire_29_valid;
  wire         sinkVec_sinkWire_29_ready;
  wire [2:0]   x13_7_0_bits_instructionIndex;
  wire [1:0]   x13_7_0_bits_offset;
  wire [4:0]   x13_7_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_28_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_28_bits_offset;
  wire [1:0]   sinkVec_sinkWire_28_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_28_bits_vs;
  wire         sinkVec_sinkWire_28_valid;
  wire         sinkVec_sinkWire_28_ready;
  wire [2:0]   x22_6_1_bits_instructionIndex;
  wire         x22_6_1_bits_last;
  wire [31:0]  x22_6_1_bits_data;
  wire [3:0]   x22_6_1_bits_mask;
  wire [1:0]   x22_6_1_bits_offset;
  wire [4:0]   x22_6_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_27_bits_instructionIndex;
  wire         sinkVec_sinkWire_27_bits_last;
  wire [31:0]  sinkVec_sinkWire_27_bits_data;
  wire [3:0]   sinkVec_sinkWire_27_bits_mask;
  wire [1:0]   sinkVec_sinkWire_27_bits_offset;
  wire [4:0]   sinkVec_sinkWire_27_bits_vd;
  wire         sinkVec_sinkWire_27_valid;
  wire         sinkVec_sinkWire_27_ready;
  wire [2:0]   x22_6_0_bits_instructionIndex;
  wire [31:0]  x22_6_0_bits_data;
  wire [3:0]   x22_6_0_bits_mask;
  wire [1:0]   x22_6_0_bits_offset;
  wire [4:0]   x22_6_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_26_bits_instructionIndex;
  wire         sinkVec_sinkWire_26_bits_last;
  wire [31:0]  sinkVec_sinkWire_26_bits_data;
  wire [3:0]   sinkVec_sinkWire_26_bits_mask;
  wire [1:0]   sinkVec_sinkWire_26_bits_offset;
  wire [4:0]   sinkVec_sinkWire_26_bits_vd;
  wire         sinkVec_sinkWire_26_valid;
  wire         sinkVec_sinkWire_26_ready;
  wire [2:0]   x13_6_1_bits_instructionIndex;
  wire [1:0]   x13_6_1_bits_offset;
  wire [4:0]   x13_6_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_25_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_25_bits_offset;
  wire [1:0]   sinkVec_sinkWire_25_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_25_bits_vs;
  wire         sinkVec_sinkWire_25_valid;
  wire         sinkVec_sinkWire_25_ready;
  wire [2:0]   x13_6_0_bits_instructionIndex;
  wire [1:0]   x13_6_0_bits_offset;
  wire [4:0]   x13_6_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_24_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_24_bits_offset;
  wire [1:0]   sinkVec_sinkWire_24_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_24_bits_vs;
  wire         sinkVec_sinkWire_24_valid;
  wire         sinkVec_sinkWire_24_ready;
  wire [2:0]   x22_5_1_bits_instructionIndex;
  wire         x22_5_1_bits_last;
  wire [31:0]  x22_5_1_bits_data;
  wire [3:0]   x22_5_1_bits_mask;
  wire [1:0]   x22_5_1_bits_offset;
  wire [4:0]   x22_5_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_23_bits_instructionIndex;
  wire         sinkVec_sinkWire_23_bits_last;
  wire [31:0]  sinkVec_sinkWire_23_bits_data;
  wire [3:0]   sinkVec_sinkWire_23_bits_mask;
  wire [1:0]   sinkVec_sinkWire_23_bits_offset;
  wire [4:0]   sinkVec_sinkWire_23_bits_vd;
  wire         sinkVec_sinkWire_23_valid;
  wire         sinkVec_sinkWire_23_ready;
  wire [2:0]   x22_5_0_bits_instructionIndex;
  wire [31:0]  x22_5_0_bits_data;
  wire [3:0]   x22_5_0_bits_mask;
  wire [1:0]   x22_5_0_bits_offset;
  wire [4:0]   x22_5_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_22_bits_instructionIndex;
  wire         sinkVec_sinkWire_22_bits_last;
  wire [31:0]  sinkVec_sinkWire_22_bits_data;
  wire [3:0]   sinkVec_sinkWire_22_bits_mask;
  wire [1:0]   sinkVec_sinkWire_22_bits_offset;
  wire [4:0]   sinkVec_sinkWire_22_bits_vd;
  wire         sinkVec_sinkWire_22_valid;
  wire         sinkVec_sinkWire_22_ready;
  wire [2:0]   x13_5_1_bits_instructionIndex;
  wire [1:0]   x13_5_1_bits_offset;
  wire [4:0]   x13_5_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_21_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_21_bits_offset;
  wire [1:0]   sinkVec_sinkWire_21_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_21_bits_vs;
  wire         sinkVec_sinkWire_21_valid;
  wire         sinkVec_sinkWire_21_ready;
  wire [2:0]   x13_5_0_bits_instructionIndex;
  wire [1:0]   x13_5_0_bits_offset;
  wire [4:0]   x13_5_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_20_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_20_bits_offset;
  wire [1:0]   sinkVec_sinkWire_20_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_20_bits_vs;
  wire         sinkVec_sinkWire_20_valid;
  wire         sinkVec_sinkWire_20_ready;
  wire [2:0]   x22_4_1_bits_instructionIndex;
  wire         x22_4_1_bits_last;
  wire [31:0]  x22_4_1_bits_data;
  wire [3:0]   x22_4_1_bits_mask;
  wire [1:0]   x22_4_1_bits_offset;
  wire [4:0]   x22_4_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_19_bits_instructionIndex;
  wire         sinkVec_sinkWire_19_bits_last;
  wire [31:0]  sinkVec_sinkWire_19_bits_data;
  wire [3:0]   sinkVec_sinkWire_19_bits_mask;
  wire [1:0]   sinkVec_sinkWire_19_bits_offset;
  wire [4:0]   sinkVec_sinkWire_19_bits_vd;
  wire         sinkVec_sinkWire_19_valid;
  wire         sinkVec_sinkWire_19_ready;
  wire [2:0]   x22_4_0_bits_instructionIndex;
  wire [31:0]  x22_4_0_bits_data;
  wire [3:0]   x22_4_0_bits_mask;
  wire [1:0]   x22_4_0_bits_offset;
  wire [4:0]   x22_4_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_18_bits_instructionIndex;
  wire         sinkVec_sinkWire_18_bits_last;
  wire [31:0]  sinkVec_sinkWire_18_bits_data;
  wire [3:0]   sinkVec_sinkWire_18_bits_mask;
  wire [1:0]   sinkVec_sinkWire_18_bits_offset;
  wire [4:0]   sinkVec_sinkWire_18_bits_vd;
  wire         sinkVec_sinkWire_18_valid;
  wire         sinkVec_sinkWire_18_ready;
  wire [2:0]   x13_4_1_bits_instructionIndex;
  wire [1:0]   x13_4_1_bits_offset;
  wire [4:0]   x13_4_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_17_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_17_bits_offset;
  wire [1:0]   sinkVec_sinkWire_17_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_17_bits_vs;
  wire         sinkVec_sinkWire_17_valid;
  wire         sinkVec_sinkWire_17_ready;
  wire [2:0]   x13_4_0_bits_instructionIndex;
  wire [1:0]   x13_4_0_bits_offset;
  wire [4:0]   x13_4_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_16_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_16_bits_offset;
  wire [1:0]   sinkVec_sinkWire_16_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_16_bits_vs;
  wire         sinkVec_sinkWire_16_valid;
  wire         sinkVec_sinkWire_16_ready;
  wire [2:0]   x22_3_1_bits_instructionIndex;
  wire         x22_3_1_bits_last;
  wire [31:0]  x22_3_1_bits_data;
  wire [3:0]   x22_3_1_bits_mask;
  wire [1:0]   x22_3_1_bits_offset;
  wire [4:0]   x22_3_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_15_bits_instructionIndex;
  wire         sinkVec_sinkWire_15_bits_last;
  wire [31:0]  sinkVec_sinkWire_15_bits_data;
  wire [3:0]   sinkVec_sinkWire_15_bits_mask;
  wire [1:0]   sinkVec_sinkWire_15_bits_offset;
  wire [4:0]   sinkVec_sinkWire_15_bits_vd;
  wire         sinkVec_sinkWire_15_valid;
  wire         sinkVec_sinkWire_15_ready;
  wire [2:0]   x22_3_0_bits_instructionIndex;
  wire [31:0]  x22_3_0_bits_data;
  wire [3:0]   x22_3_0_bits_mask;
  wire [1:0]   x22_3_0_bits_offset;
  wire [4:0]   x22_3_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_14_bits_instructionIndex;
  wire         sinkVec_sinkWire_14_bits_last;
  wire [31:0]  sinkVec_sinkWire_14_bits_data;
  wire [3:0]   sinkVec_sinkWire_14_bits_mask;
  wire [1:0]   sinkVec_sinkWire_14_bits_offset;
  wire [4:0]   sinkVec_sinkWire_14_bits_vd;
  wire         sinkVec_sinkWire_14_valid;
  wire         sinkVec_sinkWire_14_ready;
  wire [2:0]   x13_3_1_bits_instructionIndex;
  wire [1:0]   x13_3_1_bits_offset;
  wire [4:0]   x13_3_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_13_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_13_bits_offset;
  wire [1:0]   sinkVec_sinkWire_13_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_13_bits_vs;
  wire         sinkVec_sinkWire_13_valid;
  wire         sinkVec_sinkWire_13_ready;
  wire [2:0]   x13_3_0_bits_instructionIndex;
  wire [1:0]   x13_3_0_bits_offset;
  wire [4:0]   x13_3_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_12_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_12_bits_offset;
  wire [1:0]   sinkVec_sinkWire_12_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_12_bits_vs;
  wire         sinkVec_sinkWire_12_valid;
  wire         sinkVec_sinkWire_12_ready;
  wire [2:0]   x22_2_1_bits_instructionIndex;
  wire         x22_2_1_bits_last;
  wire [31:0]  x22_2_1_bits_data;
  wire [3:0]   x22_2_1_bits_mask;
  wire [1:0]   x22_2_1_bits_offset;
  wire [4:0]   x22_2_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_11_bits_instructionIndex;
  wire         sinkVec_sinkWire_11_bits_last;
  wire [31:0]  sinkVec_sinkWire_11_bits_data;
  wire [3:0]   sinkVec_sinkWire_11_bits_mask;
  wire [1:0]   sinkVec_sinkWire_11_bits_offset;
  wire [4:0]   sinkVec_sinkWire_11_bits_vd;
  wire         sinkVec_sinkWire_11_valid;
  wire         sinkVec_sinkWire_11_ready;
  wire [2:0]   x22_2_0_bits_instructionIndex;
  wire [31:0]  x22_2_0_bits_data;
  wire [3:0]   x22_2_0_bits_mask;
  wire [1:0]   x22_2_0_bits_offset;
  wire [4:0]   x22_2_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_10_bits_instructionIndex;
  wire         sinkVec_sinkWire_10_bits_last;
  wire [31:0]  sinkVec_sinkWire_10_bits_data;
  wire [3:0]   sinkVec_sinkWire_10_bits_mask;
  wire [1:0]   sinkVec_sinkWire_10_bits_offset;
  wire [4:0]   sinkVec_sinkWire_10_bits_vd;
  wire         sinkVec_sinkWire_10_valid;
  wire         sinkVec_sinkWire_10_ready;
  wire [2:0]   x13_2_1_bits_instructionIndex;
  wire [1:0]   x13_2_1_bits_offset;
  wire [4:0]   x13_2_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_9_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_9_bits_offset;
  wire [1:0]   sinkVec_sinkWire_9_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_9_bits_vs;
  wire         sinkVec_sinkWire_9_valid;
  wire         sinkVec_sinkWire_9_ready;
  wire [2:0]   x13_2_0_bits_instructionIndex;
  wire [1:0]   x13_2_0_bits_offset;
  wire [4:0]   x13_2_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_8_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_8_bits_offset;
  wire [1:0]   sinkVec_sinkWire_8_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_8_bits_vs;
  wire         sinkVec_sinkWire_8_valid;
  wire         sinkVec_sinkWire_8_ready;
  wire [2:0]   x22_1_1_bits_instructionIndex;
  wire         x22_1_1_bits_last;
  wire [31:0]  x22_1_1_bits_data;
  wire [3:0]   x22_1_1_bits_mask;
  wire [1:0]   x22_1_1_bits_offset;
  wire [4:0]   x22_1_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_7_bits_instructionIndex;
  wire         sinkVec_sinkWire_7_bits_last;
  wire [31:0]  sinkVec_sinkWire_7_bits_data;
  wire [3:0]   sinkVec_sinkWire_7_bits_mask;
  wire [1:0]   sinkVec_sinkWire_7_bits_offset;
  wire [4:0]   sinkVec_sinkWire_7_bits_vd;
  wire         sinkVec_sinkWire_7_valid;
  wire         sinkVec_sinkWire_7_ready;
  wire [2:0]   x22_1_0_bits_instructionIndex;
  wire [31:0]  x22_1_0_bits_data;
  wire [3:0]   x22_1_0_bits_mask;
  wire [1:0]   x22_1_0_bits_offset;
  wire [4:0]   x22_1_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_6_bits_instructionIndex;
  wire         sinkVec_sinkWire_6_bits_last;
  wire [31:0]  sinkVec_sinkWire_6_bits_data;
  wire [3:0]   sinkVec_sinkWire_6_bits_mask;
  wire [1:0]   sinkVec_sinkWire_6_bits_offset;
  wire [4:0]   sinkVec_sinkWire_6_bits_vd;
  wire         sinkVec_sinkWire_6_valid;
  wire         sinkVec_sinkWire_6_ready;
  wire [2:0]   x13_1_1_bits_instructionIndex;
  wire [1:0]   x13_1_1_bits_offset;
  wire [4:0]   x13_1_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_5_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_5_bits_offset;
  wire [1:0]   sinkVec_sinkWire_5_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_5_bits_vs;
  wire         sinkVec_sinkWire_5_valid;
  wire         sinkVec_sinkWire_5_ready;
  wire [2:0]   x13_1_0_bits_instructionIndex;
  wire [1:0]   x13_1_0_bits_offset;
  wire [4:0]   x13_1_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_4_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_4_bits_offset;
  wire [1:0]   sinkVec_sinkWire_4_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_4_bits_vs;
  wire         sinkVec_sinkWire_4_valid;
  wire         sinkVec_sinkWire_4_ready;
  wire [2:0]   x22_1_bits_instructionIndex;
  wire         x22_1_bits_last;
  wire [31:0]  x22_1_bits_data;
  wire [3:0]   x22_1_bits_mask;
  wire [1:0]   x22_1_bits_offset;
  wire [4:0]   x22_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_3_bits_instructionIndex;
  wire         sinkVec_sinkWire_3_bits_last;
  wire [31:0]  sinkVec_sinkWire_3_bits_data;
  wire [3:0]   sinkVec_sinkWire_3_bits_mask;
  wire [1:0]   sinkVec_sinkWire_3_bits_offset;
  wire [4:0]   sinkVec_sinkWire_3_bits_vd;
  wire         sinkVec_sinkWire_3_valid;
  wire         sinkVec_sinkWire_3_ready;
  wire [2:0]   x22_0_bits_instructionIndex;
  wire [31:0]  x22_0_bits_data;
  wire [3:0]   x22_0_bits_mask;
  wire [1:0]   x22_0_bits_offset;
  wire [4:0]   x22_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_2_bits_instructionIndex;
  wire         sinkVec_sinkWire_2_bits_last;
  wire [31:0]  sinkVec_sinkWire_2_bits_data;
  wire [3:0]   sinkVec_sinkWire_2_bits_mask;
  wire [1:0]   sinkVec_sinkWire_2_bits_offset;
  wire [4:0]   sinkVec_sinkWire_2_bits_vd;
  wire         sinkVec_sinkWire_2_valid;
  wire         sinkVec_sinkWire_2_ready;
  wire [2:0]   x13_1_bits_instructionIndex;
  wire [1:0]   x13_1_bits_offset;
  wire [4:0]   x13_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_1_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_1_bits_offset;
  wire [1:0]   sinkVec_sinkWire_1_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_1_bits_vs;
  wire         sinkVec_sinkWire_1_valid;
  wire         sinkVec_sinkWire_1_ready;
  wire [2:0]   x13_0_bits_instructionIndex;
  wire [1:0]   x13_0_bits_offset;
  wire [4:0]   x13_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_bits_instructionIndex;
  wire [1:0]   sinkVec_sinkWire_bits_offset;
  wire [1:0]   sinkVec_sinkWire_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_bits_vs;
  wire         sinkVec_sinkWire_valid;
  wire         sinkVec_sinkWire_ready;
  wire [1:0]   laneRequestSourceWire_15_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_15_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_15_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_15_bits_segment;
  wire [1:0]   laneRequestSourceWire_15_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_15_bits_vd;
  wire [4:0]   laneRequestSourceWire_15_bits_vs1;
  wire         laneRequestSourceWire_15_bits_issueInst;
  wire         laneRequestSinkWire_15_ready;
  wire [1:0]   laneRequestSourceWire_14_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_14_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_14_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_14_bits_segment;
  wire [1:0]   laneRequestSourceWire_14_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_14_bits_vd;
  wire [4:0]   laneRequestSourceWire_14_bits_vs1;
  wire         laneRequestSourceWire_14_bits_issueInst;
  wire         laneRequestSinkWire_14_ready;
  wire [1:0]   laneRequestSourceWire_13_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_13_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_13_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_13_bits_segment;
  wire [1:0]   laneRequestSourceWire_13_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_13_bits_vd;
  wire [4:0]   laneRequestSourceWire_13_bits_vs1;
  wire         laneRequestSourceWire_13_bits_issueInst;
  wire         laneRequestSinkWire_13_ready;
  wire [1:0]   laneRequestSourceWire_12_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_12_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_12_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_12_bits_segment;
  wire [1:0]   laneRequestSourceWire_12_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_12_bits_vd;
  wire [4:0]   laneRequestSourceWire_12_bits_vs1;
  wire         laneRequestSourceWire_12_bits_issueInst;
  wire         laneRequestSinkWire_12_ready;
  wire [1:0]   laneRequestSourceWire_11_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_11_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_11_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_11_bits_segment;
  wire [1:0]   laneRequestSourceWire_11_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_11_bits_vd;
  wire [4:0]   laneRequestSourceWire_11_bits_vs1;
  wire         laneRequestSourceWire_11_bits_issueInst;
  wire         laneRequestSinkWire_11_ready;
  wire [1:0]   laneRequestSourceWire_10_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_10_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_10_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_10_bits_segment;
  wire [1:0]   laneRequestSourceWire_10_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_10_bits_vd;
  wire [4:0]   laneRequestSourceWire_10_bits_vs1;
  wire         laneRequestSourceWire_10_bits_issueInst;
  wire         laneRequestSinkWire_10_ready;
  wire [1:0]   laneRequestSourceWire_9_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_9_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_9_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_9_bits_segment;
  wire [1:0]   laneRequestSourceWire_9_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_9_bits_vd;
  wire [4:0]   laneRequestSourceWire_9_bits_vs1;
  wire         laneRequestSourceWire_9_bits_issueInst;
  wire         laneRequestSinkWire_9_ready;
  wire [1:0]   laneRequestSourceWire_8_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_8_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_8_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_8_bits_segment;
  wire [1:0]   laneRequestSourceWire_8_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_8_bits_vd;
  wire [4:0]   laneRequestSourceWire_8_bits_vs1;
  wire         laneRequestSourceWire_8_bits_issueInst;
  wire         laneRequestSinkWire_8_ready;
  wire [1:0]   laneRequestSourceWire_7_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_7_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_7_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_7_bits_segment;
  wire [1:0]   laneRequestSourceWire_7_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_7_bits_vd;
  wire [4:0]   laneRequestSourceWire_7_bits_vs1;
  wire         laneRequestSourceWire_7_bits_issueInst;
  wire         laneRequestSinkWire_7_ready;
  wire [1:0]   laneRequestSourceWire_6_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_6_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_6_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_6_bits_segment;
  wire [1:0]   laneRequestSourceWire_6_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_6_bits_vd;
  wire [4:0]   laneRequestSourceWire_6_bits_vs1;
  wire         laneRequestSourceWire_6_bits_issueInst;
  wire         laneRequestSinkWire_6_ready;
  wire [1:0]   laneRequestSourceWire_5_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_5_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_5_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_5_bits_segment;
  wire [1:0]   laneRequestSourceWire_5_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_5_bits_vd;
  wire [4:0]   laneRequestSourceWire_5_bits_vs1;
  wire         laneRequestSourceWire_5_bits_issueInst;
  wire         laneRequestSinkWire_5_ready;
  wire [1:0]   laneRequestSourceWire_4_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_4_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_4_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_4_bits_segment;
  wire [1:0]   laneRequestSourceWire_4_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_4_bits_vd;
  wire [4:0]   laneRequestSourceWire_4_bits_vs1;
  wire         laneRequestSourceWire_4_bits_issueInst;
  wire         laneRequestSinkWire_4_ready;
  wire [1:0]   laneRequestSourceWire_3_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_3_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_3_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_3_bits_segment;
  wire [1:0]   laneRequestSourceWire_3_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_3_bits_vd;
  wire [4:0]   laneRequestSourceWire_3_bits_vs1;
  wire         laneRequestSourceWire_3_bits_issueInst;
  wire         laneRequestSinkWire_3_ready;
  wire [1:0]   laneRequestSourceWire_2_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_2_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_2_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_2_bits_segment;
  wire [1:0]   laneRequestSourceWire_2_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_2_bits_vd;
  wire [4:0]   laneRequestSourceWire_2_bits_vs1;
  wire         laneRequestSourceWire_2_bits_issueInst;
  wire         laneRequestSinkWire_2_ready;
  wire [1:0]   laneRequestSourceWire_1_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_1_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_1_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_1_bits_segment;
  wire [1:0]   laneRequestSourceWire_1_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_1_bits_vd;
  wire [4:0]   laneRequestSourceWire_1_bits_vs1;
  wire         laneRequestSourceWire_1_bits_issueInst;
  wire         laneRequestSinkWire_1_ready;
  wire [1:0]   laneRequestSourceWire_0_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_0_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_0_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_0_bits_segment;
  wire [1:0]   laneRequestSourceWire_0_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_0_bits_vd;
  wire [4:0]   laneRequestSourceWire_0_bits_vs1;
  wire         laneRequestSourceWire_0_bits_issueInst;
  wire         laneRequestSinkWire_0_ready;
  wire [1:0]   requestRegCSR_vxrm;
  wire [11:0]  requestRegCSR_vStart;
  wire         requestRegCSR_vma;
  wire         requestRegCSR_vta;
  wire [2:0]   requestRegCSR_vlmul;
  wire         indexedLoadStorePort_aw_ready_0 = indexedLoadStorePort_aw_ready;
  wire         indexedLoadStorePort_w_ready_0 = indexedLoadStorePort_w_ready;
  wire         indexedLoadStorePort_b_valid_0 = indexedLoadStorePort_b_valid;
  wire [1:0]   indexedLoadStorePort_b_bits_id_0 = indexedLoadStorePort_b_bits_id;
  wire [1:0]   indexedLoadStorePort_b_bits_resp_0 = indexedLoadStorePort_b_bits_resp;
  wire         indexedLoadStorePort_ar_ready_0 = indexedLoadStorePort_ar_ready;
  wire         indexedLoadStorePort_r_valid_0 = indexedLoadStorePort_r_valid;
  wire [1:0]   indexedLoadStorePort_r_bits_id_0 = indexedLoadStorePort_r_bits_id;
  wire [31:0]  indexedLoadStorePort_r_bits_data_0 = indexedLoadStorePort_r_bits_data;
  wire [1:0]   indexedLoadStorePort_r_bits_resp_0 = indexedLoadStorePort_r_bits_resp;
  wire         indexedLoadStorePort_r_bits_last_0 = indexedLoadStorePort_r_bits_last;
  wire         highBandwidthLoadStorePort_aw_ready_0 = highBandwidthLoadStorePort_aw_ready;
  wire         highBandwidthLoadStorePort_w_ready_0 = highBandwidthLoadStorePort_w_ready;
  wire         highBandwidthLoadStorePort_b_valid_0 = highBandwidthLoadStorePort_b_valid;
  wire [1:0]   highBandwidthLoadStorePort_b_bits_id_0 = highBandwidthLoadStorePort_b_bits_id;
  wire [1:0]   highBandwidthLoadStorePort_b_bits_resp_0 = highBandwidthLoadStorePort_b_bits_resp;
  wire         highBandwidthLoadStorePort_ar_ready_0 = highBandwidthLoadStorePort_ar_ready;
  wire         highBandwidthLoadStorePort_r_valid_0 = highBandwidthLoadStorePort_r_valid;
  wire [1:0]   highBandwidthLoadStorePort_r_bits_id_0 = highBandwidthLoadStorePort_r_bits_id;
  wire [511:0] highBandwidthLoadStorePort_r_bits_data_0 = highBandwidthLoadStorePort_r_bits_data;
  wire [1:0]   highBandwidthLoadStorePort_r_bits_resp_0 = highBandwidthLoadStorePort_r_bits_resp;
  wire         highBandwidthLoadStorePort_r_bits_last_0 = highBandwidthLoadStorePort_r_bits_last;
  wire         issue_valid_0 = issue_valid;
  wire [31:0]  issue_bits_instruction_0 = issue_bits_instruction;
  wire [31:0]  issue_bits_rs1Data_0 = issue_bits_rs1Data;
  wire [31:0]  issue_bits_rs2Data_0 = issue_bits_rs2Data;
  wire [31:0]  issue_bits_vtype_0 = issue_bits_vtype;
  wire [31:0]  issue_bits_vl_0 = issue_bits_vl;
  wire [31:0]  issue_bits_vstart_0 = issue_bits_vstart;
  wire [31:0]  issue_bits_vcsr_0 = issue_bits_vcsr;
  wire [2:0]   highBandwidthLoadStorePort_aw_bits_size_0 = 3'h6;
  wire [2:0]   highBandwidthLoadStorePort_ar_bits_size_0 = 3'h6;
  wire [1:0]   indexedLoadStorePort_ar_bits_id_0 = 2'h0;
  wire [1:0]   highBandwidthLoadStorePort_ar_bits_id_0 = 2'h0;
  wire [7:0]   indexedLoadStorePort_aw_bits_len_0 = 8'h0;
  wire [7:0]   indexedLoadStorePort_ar_bits_len_0 = 8'h0;
  wire [7:0]   highBandwidthLoadStorePort_aw_bits_len_0 = 8'h0;
  wire [7:0]   highBandwidthLoadStorePort_ar_bits_len_0 = 8'h0;
  wire [2:0]   indexedLoadStorePort_ar_bits_size_0 = 3'h2;
  wire [1:0]   indexedLoadStorePort_aw_bits_burst_0 = 2'h1;
  wire [1:0]   indexedLoadStorePort_ar_bits_burst_0 = 2'h1;
  wire [1:0]   highBandwidthLoadStorePort_aw_bits_burst_0 = 2'h1;
  wire [1:0]   highBandwidthLoadStorePort_ar_bits_burst_0 = 2'h1;
  wire [2:0]   indexedLoadStorePort_aw_bits_prot_0 = 3'h0;
  wire [2:0]   indexedLoadStorePort_ar_bits_prot_0 = 3'h0;
  wire [2:0]   highBandwidthLoadStorePort_aw_bits_prot_0 = 3'h0;
  wire [2:0]   highBandwidthLoadStorePort_ar_bits_prot_0 = 3'h0;
  wire [31:0]  retire_csr_bits_fflag_0 = 32'h0;
  wire [3:0]   indexedLoadStorePort_aw_bits_cache_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_aw_bits_qos_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_aw_bits_region_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_cache_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_qos_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_region_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_cache_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_qos_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_region_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_cache_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_qos_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_region_0 = 4'h0;
  wire [1:0]   x13_0_bits_readSource = 2'h2;
  wire [1:0]   x13_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_1_bits_readSource = 2'h2;
  wire [1:0]   x13_1_0_bits_readSource = 2'h2;
  wire [1:0]   x13_1_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_4_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_5_bits_readSource = 2'h2;
  wire [1:0]   x13_2_0_bits_readSource = 2'h2;
  wire [1:0]   x13_2_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_8_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_9_bits_readSource = 2'h2;
  wire [1:0]   x13_3_0_bits_readSource = 2'h2;
  wire [1:0]   x13_3_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_12_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_13_bits_readSource = 2'h2;
  wire [1:0]   x13_4_0_bits_readSource = 2'h2;
  wire [1:0]   x13_4_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_16_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_17_bits_readSource = 2'h2;
  wire [1:0]   x13_5_0_bits_readSource = 2'h2;
  wire [1:0]   x13_5_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_20_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_21_bits_readSource = 2'h2;
  wire [1:0]   x13_6_0_bits_readSource = 2'h2;
  wire [1:0]   x13_6_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_24_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_25_bits_readSource = 2'h2;
  wire [1:0]   x13_7_0_bits_readSource = 2'h2;
  wire [1:0]   x13_7_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_28_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_29_bits_readSource = 2'h2;
  wire [1:0]   x13_8_0_bits_readSource = 2'h2;
  wire [1:0]   x13_8_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_32_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_33_bits_readSource = 2'h2;
  wire [1:0]   x13_9_0_bits_readSource = 2'h2;
  wire [1:0]   x13_9_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_36_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_37_bits_readSource = 2'h2;
  wire [1:0]   x13_10_0_bits_readSource = 2'h2;
  wire [1:0]   x13_10_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_40_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_41_bits_readSource = 2'h2;
  wire [1:0]   x13_11_0_bits_readSource = 2'h2;
  wire [1:0]   x13_11_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_44_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_45_bits_readSource = 2'h2;
  wire [1:0]   x13_12_0_bits_readSource = 2'h2;
  wire [1:0]   x13_12_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_48_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_49_bits_readSource = 2'h2;
  wire [1:0]   x13_13_0_bits_readSource = 2'h2;
  wire [1:0]   x13_13_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_52_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_53_bits_readSource = 2'h2;
  wire [1:0]   x13_14_0_bits_readSource = 2'h2;
  wire [1:0]   x13_14_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_56_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_57_bits_readSource = 2'h2;
  wire [1:0]   x13_15_0_bits_readSource = 2'h2;
  wire [1:0]   x13_15_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_60_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_61_bits_readSource = 2'h2;
  wire [1:0]   lo_lo_lo = 2'h3;
  wire [1:0]   lo_lo_hi = 2'h3;
  wire [1:0]   lo_hi_lo = 2'h3;
  wire [1:0]   lo_hi_hi = 2'h3;
  wire [1:0]   hi_lo_lo = 2'h3;
  wire [1:0]   hi_lo_hi = 2'h3;
  wire [1:0]   hi_hi_lo = 2'h3;
  wire [1:0]   hi_hi_hi = 2'h3;
  wire [1:0]   lo_lo_lo_1 = 2'h3;
  wire [1:0]   lo_lo_hi_1 = 2'h3;
  wire [1:0]   lo_hi_lo_1 = 2'h3;
  wire [1:0]   lo_hi_hi_1 = 2'h3;
  wire [1:0]   hi_lo_lo_1 = 2'h3;
  wire [1:0]   hi_lo_hi_1 = 2'h3;
  wire [1:0]   hi_hi_lo_1 = 2'h3;
  wire [1:0]   hi_hi_hi_1 = 2'h3;
  wire [3:0]   lo_lo = 4'hF;
  wire [3:0]   lo_hi = 4'hF;
  wire [3:0]   hi_lo = 4'hF;
  wire [3:0]   hi_hi = 4'hF;
  wire [3:0]   lo_lo_1 = 4'hF;
  wire [3:0]   lo_hi_1 = 4'hF;
  wire [3:0]   hi_lo_1 = 4'hF;
  wire [3:0]   hi_hi_1 = 4'hF;
  wire [7:0]   lo = 8'hFF;
  wire [7:0]   hi = 8'hFF;
  wire [7:0]   lo_1 = 8'hFF;
  wire [7:0]   hi_1 = 8'hFF;
  wire         indexedLoadStorePort_w_bits_last_0 = 1'h1;
  wire         indexedLoadStorePort_b_ready_0 = 1'h1;
  wire         highBandwidthLoadStorePort_w_bits_last_0 = 1'h1;
  wire         highBandwidthLoadStorePort_b_ready_0 = 1'h1;
  wire [2:0]   vSewOHForMask = 3'h1;
  wire         indexedLoadStorePort_aw_bits_lock_0 = 1'h0;
  wire         indexedLoadStorePort_ar_bits_lock_0 = 1'h0;
  wire         highBandwidthLoadStorePort_aw_bits_lock_0 = 1'h0;
  wire         highBandwidthLoadStorePort_ar_bits_lock_0 = 1'h0;
  wire         retire_csr_valid_0 = 1'h0;
  wire         x22_0_bits_last = 1'h0;
  wire         sinkVec_queue_2_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_2_bits_last = 1'h0;
  wire         sinkVec_validSink_2_bits_last = 1'h0;
  wire         x22_1_0_bits_last = 1'h0;
  wire         sinkVec_queue_6_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_6_bits_last = 1'h0;
  wire         sinkVec_validSink_6_bits_last = 1'h0;
  wire         x22_2_0_bits_last = 1'h0;
  wire         sinkVec_queue_10_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_10_bits_last = 1'h0;
  wire         sinkVec_validSink_10_bits_last = 1'h0;
  wire         x22_3_0_bits_last = 1'h0;
  wire         sinkVec_queue_14_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_14_bits_last = 1'h0;
  wire         sinkVec_validSink_14_bits_last = 1'h0;
  wire         x22_4_0_bits_last = 1'h0;
  wire         sinkVec_queue_18_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_18_bits_last = 1'h0;
  wire         sinkVec_validSink_18_bits_last = 1'h0;
  wire         x22_5_0_bits_last = 1'h0;
  wire         sinkVec_queue_22_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_22_bits_last = 1'h0;
  wire         sinkVec_validSink_22_bits_last = 1'h0;
  wire         x22_6_0_bits_last = 1'h0;
  wire         sinkVec_queue_26_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_26_bits_last = 1'h0;
  wire         sinkVec_validSink_26_bits_last = 1'h0;
  wire         x22_7_0_bits_last = 1'h0;
  wire         sinkVec_queue_30_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_30_bits_last = 1'h0;
  wire         sinkVec_validSink_30_bits_last = 1'h0;
  wire         x22_8_0_bits_last = 1'h0;
  wire         sinkVec_queue_34_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_34_bits_last = 1'h0;
  wire         sinkVec_validSink_34_bits_last = 1'h0;
  wire         x22_9_0_bits_last = 1'h0;
  wire         sinkVec_queue_38_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_38_bits_last = 1'h0;
  wire         sinkVec_validSink_38_bits_last = 1'h0;
  wire         x22_10_0_bits_last = 1'h0;
  wire         sinkVec_queue_42_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_42_bits_last = 1'h0;
  wire         sinkVec_validSink_42_bits_last = 1'h0;
  wire         x22_11_0_bits_last = 1'h0;
  wire         sinkVec_queue_46_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_46_bits_last = 1'h0;
  wire         sinkVec_validSink_46_bits_last = 1'h0;
  wire         x22_12_0_bits_last = 1'h0;
  wire         sinkVec_queue_50_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_50_bits_last = 1'h0;
  wire         sinkVec_validSink_50_bits_last = 1'h0;
  wire         x22_13_0_bits_last = 1'h0;
  wire         sinkVec_queue_54_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_54_bits_last = 1'h0;
  wire         sinkVec_validSink_54_bits_last = 1'h0;
  wire         x22_14_0_bits_last = 1'h0;
  wire         sinkVec_queue_58_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_58_bits_last = 1'h0;
  wire         sinkVec_validSink_58_bits_last = 1'h0;
  wire         x22_15_0_bits_last = 1'h0;
  wire         sinkVec_queue_62_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_62_bits_last = 1'h0;
  wire         sinkVec_validSink_62_bits_last = 1'h0;
  reg  [2:0]   instructionCounter;
  wire [2:0]   nextInstructionCounter = instructionCounter + 3'h1;
  wire         issue_ready_0;
  wire         _probeWire_issue_valid_T = issue_ready_0 & issue_valid_0;
  reg  [2:0]   responseCounter;
  wire [2:0]   nextResponseCounter = responseCounter + 3'h1;
  reg          requestReg_valid;
  wire         requestRegDequeue_valid = requestReg_valid;
  reg  [31:0]  requestReg_bits_issue_instruction;
  wire [31:0]  requestRegDequeue_bits_instruction = requestReg_bits_issue_instruction;
  reg  [31:0]  requestReg_bits_issue_rs1Data;
  wire [31:0]  requestRegDequeue_bits_rs1Data = requestReg_bits_issue_rs1Data;
  reg  [31:0]  requestReg_bits_issue_rs2Data;
  wire [31:0]  requestRegDequeue_bits_rs2Data = requestReg_bits_issue_rs2Data;
  reg  [31:0]  requestReg_bits_issue_vtype;
  wire [31:0]  requestRegDequeue_bits_vtype = requestReg_bits_issue_vtype;
  reg  [31:0]  requestReg_bits_issue_vl;
  wire [31:0]  requestRegDequeue_bits_vl = requestReg_bits_issue_vl;
  reg  [31:0]  requestReg_bits_issue_vstart;
  wire [31:0]  requestRegDequeue_bits_vstart = requestReg_bits_issue_vstart;
  reg  [31:0]  requestReg_bits_issue_vcsr;
  wire [31:0]  requestRegDequeue_bits_vcsr = requestReg_bits_issue_vcsr;
  reg          requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_0_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_1_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_2_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_3_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_4_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_5_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_6_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_7_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_8_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_9_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_10_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_11_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_12_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_13_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_14_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  wire         laneRequestSourceWire_15_bits_decodeResult_orderReduce = requestReg_bits_decodeResult_orderReduce;
  reg          requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_0_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_1_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_2_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_3_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_4_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_5_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_6_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_7_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_8_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_9_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_10_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_11_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_12_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_13_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_14_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  wire         laneRequestSourceWire_15_bits_decodeResult_floatMul = requestReg_bits_decodeResult_floatMul;
  reg  [1:0]   requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_0_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_1_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_2_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_3_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_4_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_5_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_6_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_7_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_8_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_9_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_10_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_11_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_12_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_13_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_14_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  wire [1:0]   laneRequestSourceWire_15_bits_decodeResult_fpExecutionType = requestReg_bits_decodeResult_fpExecutionType;
  reg          requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_0_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_1_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_2_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_3_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_4_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_5_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_6_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_7_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_8_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_9_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_10_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_11_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_12_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_13_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_14_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  wire         laneRequestSourceWire_15_bits_decodeResult_float = requestReg_bits_decodeResult_float;
  reg          requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_0_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_1_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_2_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_3_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_4_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_5_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_6_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_7_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_8_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_9_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_10_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_11_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_12_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_13_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_14_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_15_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  reg  [4:0]   requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_0_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_1_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_2_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_3_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_4_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_5_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_6_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_7_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_8_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_9_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_10_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_11_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_12_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_13_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_14_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_15_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  reg          requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_0_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_1_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_2_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_3_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_4_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_5_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_6_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_7_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_8_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_9_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_10_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_11_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_12_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_13_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_14_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_15_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  reg          requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_0_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_1_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_2_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_3_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_4_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_5_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_6_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_7_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_8_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_9_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_10_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_11_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_12_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_13_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_14_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_15_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  reg          requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_0_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_1_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_2_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_3_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_4_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_5_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_6_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_7_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_8_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_9_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_10_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_11_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_12_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_13_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_14_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_15_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  reg          requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_0_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_1_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_2_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_3_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_4_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_5_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_6_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_7_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_8_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_9_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_10_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_11_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_12_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_13_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_14_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_15_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  reg          requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_0_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_1_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_2_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_3_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_4_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_5_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_6_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_7_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_8_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_9_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_10_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_11_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_12_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_13_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_14_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_15_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  reg          requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_0_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_1_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_2_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_3_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_4_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_5_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_6_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_7_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_8_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_9_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_10_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_11_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_12_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_13_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_14_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_15_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  reg          requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_0_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_1_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_2_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_3_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_4_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_5_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_6_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_7_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_8_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_9_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_10_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_11_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_12_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_13_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_14_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_15_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  reg          requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_0_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_1_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_2_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_3_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_4_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_5_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_6_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_7_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_8_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_9_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_10_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_11_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_12_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_13_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_14_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_15_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  reg          requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_8_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_9_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_10_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_11_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_12_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_13_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_14_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_15_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  reg          requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_0_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_1_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_2_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_3_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_4_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_5_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_6_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_7_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_8_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_9_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_10_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_11_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_12_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_13_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_14_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_15_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  reg          requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_8_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_9_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_10_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_11_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_12_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_13_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_14_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_15_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  reg          requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_8_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_9_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_10_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_11_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_12_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_13_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_14_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_15_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  reg          requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_0_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_1_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_2_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_3_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_4_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_5_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_6_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_7_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_8_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_9_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_10_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_11_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_12_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_13_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_14_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_15_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  reg          requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_0_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_1_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_2_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_3_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_4_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_5_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_6_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_7_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_8_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_9_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_10_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_11_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_12_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_13_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_14_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_15_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  reg          requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_0_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_1_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_2_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_3_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_4_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_5_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_6_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_7_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_8_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_9_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_10_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_11_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_12_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_13_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_14_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_15_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  reg          requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_0_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_1_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_2_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_3_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_4_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_5_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_6_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_7_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_8_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_9_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_10_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_11_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_12_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_13_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_14_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_15_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  reg          requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_8_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_9_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_10_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_11_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_12_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_13_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_14_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_15_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  reg          requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_8_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_9_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_10_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_11_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_12_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_13_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_14_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_15_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  reg          requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_8_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_9_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_10_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_11_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_12_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_13_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_14_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_15_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  reg  [3:0]   requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_0_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_1_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_2_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_3_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_4_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_5_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_6_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_7_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_8_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_9_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_10_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_11_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_12_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_13_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_14_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_15_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  reg          requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_0_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_1_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_2_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_3_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_4_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_5_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_6_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_7_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_8_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_9_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_10_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_11_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_12_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_13_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_14_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_15_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  reg          requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_0_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_1_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_2_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_3_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_4_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_5_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_6_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_7_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_8_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_9_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_10_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_11_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_12_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_13_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_14_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_15_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  reg          requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_0_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_1_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_2_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_3_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_4_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_5_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_6_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_7_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_8_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_9_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_10_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_11_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_12_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_13_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_14_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_15_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  reg          requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_8_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_9_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_10_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_11_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_12_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_13_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_14_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_15_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  reg          requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_0_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_1_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_2_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_3_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_4_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_5_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_6_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_7_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_8_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_9_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_10_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_11_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_12_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_13_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_14_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_15_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  reg          requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_0_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_1_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_2_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_3_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_4_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_5_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_6_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_7_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_8_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_9_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_10_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_11_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_12_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_13_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_14_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_15_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  reg          requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_0_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_1_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_2_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_3_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_4_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_5_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_6_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_7_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_8_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_9_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_10_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_11_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_12_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_13_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_14_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_15_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  reg          requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_0_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_1_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_2_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_3_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_4_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_5_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_6_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_7_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_8_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_9_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_10_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_11_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_12_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_13_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_14_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_15_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  reg          requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_0_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_1_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_2_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_3_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_4_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_5_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_6_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_7_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_8_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_9_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_10_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_11_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_12_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_13_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_14_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_15_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  reg          requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_0_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_1_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_2_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_3_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_4_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_5_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_6_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_7_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_8_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_9_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_10_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_11_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_12_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_13_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_14_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_15_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  reg          requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_0_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_1_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_2_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_3_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_4_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_5_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_6_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_7_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_8_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_9_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_10_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_11_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_12_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_13_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_14_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_15_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  reg          requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_0_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_1_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_2_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_3_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_4_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_5_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_6_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_7_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_8_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_9_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_10_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_11_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_12_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_13_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_14_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_15_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  reg          requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_0_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_1_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_2_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_3_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_4_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_5_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_6_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_7_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_8_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_9_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_10_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_11_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_12_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_13_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_14_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_15_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  reg          requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_0_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_1_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_2_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_3_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_4_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_5_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_6_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_7_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_8_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_9_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_10_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_11_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_12_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_13_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_14_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_15_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  reg          requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_0_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_1_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_2_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_3_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_4_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_5_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_6_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_7_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_8_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_9_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_10_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_11_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_12_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_13_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_14_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_15_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  reg          requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_0_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_1_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_2_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_3_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_4_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_5_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_6_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_7_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_8_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_9_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_10_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_11_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_12_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_13_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_14_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_15_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  reg          requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_0_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_1_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_2_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_3_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_4_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_5_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_6_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_7_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_8_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_9_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_10_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_11_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_12_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_13_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_14_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_15_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  reg          requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_0_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_1_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_2_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_3_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_4_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_5_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_6_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_7_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_8_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_9_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_10_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_11_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_12_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_13_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_14_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_15_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  reg          requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_0_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_1_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_2_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_3_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_4_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_5_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_6_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_7_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_8_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_9_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_10_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_11_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_12_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_13_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_14_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_15_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  reg          requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_0_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_1_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_2_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_3_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_4_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_5_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_6_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_7_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_8_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_9_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_10_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_11_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_12_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_13_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_14_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_15_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  reg          requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_0_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_1_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_2_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_3_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_4_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_5_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_6_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_7_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_8_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_9_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_10_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_11_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_12_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_13_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_14_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_15_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  reg          requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_0_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_1_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_2_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_3_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_4_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_5_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_6_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_7_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_8_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_9_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_10_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_11_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_12_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_13_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_14_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_15_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  reg  [2:0]   requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_0_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_1_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_2_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_3_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_4_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_5_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_6_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_7_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_8_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_9_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_10_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_11_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_12_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_13_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_14_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_15_bits_instructionIndex = requestReg_bits_instructionIndex;
  reg          requestReg_bits_vdIsV0;
  reg  [11:0]  requestReg_bits_writeByte;
  wire [11:0]  laneRequestSourceWire_0_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_1_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_2_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_3_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_4_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_5_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_6_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_7_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_8_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_9_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_10_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_11_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_12_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_13_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_14_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_15_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [2:0]   laneRequestSourceWire_0_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_1_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_2_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_3_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_4_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_5_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_6_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_7_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_8_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_9_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_10_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_11_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_12_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_13_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_14_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_15_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [1:0]   laneRequestSourceWire_0_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_1_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_2_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_3_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_4_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_5_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_6_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_7_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_8_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_9_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_10_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_11_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_12_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_13_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_14_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_15_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire         laneRequestSourceWire_0_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_1_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_2_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_3_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_4_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_5_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_6_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_7_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_8_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_9_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_10_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_11_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_12_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_13_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_14_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_15_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_0_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_1_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_2_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_3_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_4_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_5_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_6_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_7_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_8_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_9_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_10_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_11_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_12_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_13_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_14_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_15_bits_csrInterface_vma = requestRegCSR_vma;
  assign requestRegCSR_vlmul = requestReg_bits_issue_vtype[2:0];
  wire [1:0]   requestRegCSR_vSew = requestReg_bits_issue_vtype[4:3];
  assign requestRegCSR_vta = requestReg_bits_issue_vtype[6];
  assign requestRegCSR_vma = requestReg_bits_issue_vtype[7];
  wire [11:0]  requestRegCSR_vl = requestReg_bits_issue_vl[11:0];
  assign requestRegCSR_vStart = requestReg_bits_issue_vstart[11:0];
  assign requestRegCSR_vxrm = requestReg_bits_issue_vcsr[2:1];
  wire         requestRegDequeue_ready;
  wire         maskUnit_gatherData_ready = requestRegDequeue_ready & requestRegDequeue_valid;
  wire         laneRequestSourceWire_0_valid;
  assign laneRequestSourceWire_0_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_1_valid;
  assign laneRequestSourceWire_1_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_2_valid;
  assign laneRequestSourceWire_2_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_3_valid;
  assign laneRequestSourceWire_3_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_4_valid;
  assign laneRequestSourceWire_4_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_5_valid;
  assign laneRequestSourceWire_5_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_6_valid;
  assign laneRequestSourceWire_6_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_7_valid;
  assign laneRequestSourceWire_7_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_8_valid;
  assign laneRequestSourceWire_8_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_9_valid;
  assign laneRequestSourceWire_9_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_10_valid;
  assign laneRequestSourceWire_10_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_11_valid;
  assign laneRequestSourceWire_11_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_12_valid;
  assign laneRequestSourceWire_12_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_13_valid;
  assign laneRequestSourceWire_13_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_14_valid;
  assign laneRequestSourceWire_14_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_15_valid;
  assign laneRequestSourceWire_15_valid = maskUnit_gatherData_ready;
  assign issue_ready_0 = ~requestReg_valid | requestRegDequeue_ready;
  wire         isLoadStoreType = ~(requestRegDequeue_bits_instruction[6]) & requestRegDequeue_valid;
  wire         laneRequestSourceWire_0_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_1_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_2_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_3_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_4_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_5_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_6_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_7_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_8_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_9_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_10_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_11_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_12_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_13_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_14_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_15_bits_loadStore = isLoadStoreType;
  wire         isStoreType = ~(requestRegDequeue_bits_instruction[6]) & requestRegDequeue_bits_instruction[5];
  wire         laneRequestSourceWire_0_bits_store = isStoreType;
  wire         laneRequestSourceWire_1_bits_store = isStoreType;
  wire         laneRequestSourceWire_2_bits_store = isStoreType;
  wire         laneRequestSourceWire_3_bits_store = isStoreType;
  wire         laneRequestSourceWire_4_bits_store = isStoreType;
  wire         laneRequestSourceWire_5_bits_store = isStoreType;
  wire         laneRequestSourceWire_6_bits_store = isStoreType;
  wire         laneRequestSourceWire_7_bits_store = isStoreType;
  wire         laneRequestSourceWire_8_bits_store = isStoreType;
  wire         laneRequestSourceWire_9_bits_store = isStoreType;
  wire         laneRequestSourceWire_10_bits_store = isStoreType;
  wire         laneRequestSourceWire_11_bits_store = isStoreType;
  wire         laneRequestSourceWire_12_bits_store = isStoreType;
  wire         laneRequestSourceWire_13_bits_store = isStoreType;
  wire         laneRequestSourceWire_14_bits_store = isStoreType;
  wire         laneRequestSourceWire_15_bits_store = isStoreType;
  wire         maskType = ~(requestRegDequeue_bits_instruction[25]);
  wire         laneRequestSourceWire_0_bits_mask = maskType;
  wire         laneRequestSourceWire_1_bits_mask = maskType;
  wire         laneRequestSourceWire_2_bits_mask = maskType;
  wire         laneRequestSourceWire_3_bits_mask = maskType;
  wire         laneRequestSourceWire_4_bits_mask = maskType;
  wire         laneRequestSourceWire_5_bits_mask = maskType;
  wire         laneRequestSourceWire_6_bits_mask = maskType;
  wire         laneRequestSourceWire_7_bits_mask = maskType;
  wire         laneRequestSourceWire_8_bits_mask = maskType;
  wire         laneRequestSourceWire_9_bits_mask = maskType;
  wire         laneRequestSourceWire_10_bits_mask = maskType;
  wire         laneRequestSourceWire_11_bits_mask = maskType;
  wire         laneRequestSourceWire_12_bits_mask = maskType;
  wire         laneRequestSourceWire_13_bits_mask = maskType;
  wire         laneRequestSourceWire_14_bits_mask = maskType;
  wire         laneRequestSourceWire_15_bits_mask = maskType;
  wire [4:0]   laneRequestSourceWire_0_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_1_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_2_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_3_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_4_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_5_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_6_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_7_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_8_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_9_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_10_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_11_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_12_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_13_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_14_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_15_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire         lsWholeReg = isLoadStoreType & requestRegDequeue_bits_instruction[27:26] == 2'h0 & requestRegDequeue_bits_instruction[24:20] == 5'h8;
  wire         laneRequestSourceWire_0_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_1_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_2_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_3_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_4_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_5_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_6_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_7_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_8_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_9_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_10_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_11_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_12_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_13_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_14_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_15_bits_lsWholeReg = lsWholeReg;
  wire         maskUnitInstruction = requestReg_bits_decodeResult_slid | requestReg_bits_decodeResult_mv;
  wire         skipLastFromLane = isStoreType | maskUnitInstruction | requestReg_bits_decodeResult_readOnly;
  wire         instructionValid = requestReg_bits_issue_vl > requestReg_bits_issue_vstart;
  wire         noOffsetReadLoadStore = isLoadStoreType & ~(requestRegDequeue_bits_instruction[26]);
  wire [7:0]   vSew1H = 8'h1 << requestReg_bits_issue_vtype[5:3];
  wire [31:0]  source1Extend =
    (vSew1H[0] ? {{24{requestRegDequeue_bits_rs1Data[7] & ~requestReg_bits_decodeResult_unsigned0}}, requestRegDequeue_bits_rs1Data[7:0]} : 32'h0)
    | (vSew1H[1] ? {{16{requestRegDequeue_bits_rs1Data[15] & ~requestReg_bits_decodeResult_unsigned0}}, requestRegDequeue_bits_rs1Data[15:0]} : 32'h0) | (vSew1H[2] ? requestRegDequeue_bits_rs1Data : 32'h0);
  wire         src1IsSInt;
  assign src1IsSInt = ~requestReg_bits_decodeResult_unsigned0;
  wire [4:0]   imm = requestReg_bits_issue_instruction[19:15];
  wire [31:0]  immSignExtend = {{16{imm[4] & (vSew1H[2] | src1IsSInt)}}, {8{imm[4] & (vSew1H[1] | vSew1H[2] | src1IsSInt)}}, {3{imm[4]}}, imm};
  wire         slotCommit_3;
  wire [3:0]   vxsatReportVec_0;
  wire [3:0]   vxsatReportVec_1;
  wire [3:0]   vxsatReportVec_2;
  wire [3:0]   vxsatReportVec_3;
  wire [3:0]   vxsatReportVec_4;
  wire [3:0]   vxsatReportVec_5;
  wire [3:0]   vxsatReportVec_6;
  wire [3:0]   vxsatReportVec_7;
  wire [3:0]   vxsatReportVec_8;
  wire [3:0]   vxsatReportVec_9;
  wire [3:0]   vxsatReportVec_10;
  wire [3:0]   vxsatReportVec_11;
  wire [3:0]   vxsatReportVec_12;
  wire [3:0]   vxsatReportVec_13;
  wire [3:0]   vxsatReportVec_14;
  wire [3:0]   vxsatReportVec_15;
  wire [3:0]   vxsatReport =
    vxsatReportVec_0 | vxsatReportVec_1 | vxsatReportVec_2 | vxsatReportVec_3 | vxsatReportVec_4 | vxsatReportVec_5 | vxsatReportVec_6 | vxsatReportVec_7 | vxsatReportVec_8 | vxsatReportVec_9 | vxsatReportVec_10 | vxsatReportVec_11
    | vxsatReportVec_12 | vxsatReportVec_13 | vxsatReportVec_14 | vxsatReportVec_15;
  wire         specialInstruction = requestReg_bits_decodeResult_special | requestReg_bits_vdIsV0;
  wire         laneRequestSourceWire_0_bits_special = specialInstruction;
  wire         laneRequestSourceWire_1_bits_special = specialInstruction;
  wire         laneRequestSourceWire_2_bits_special = specialInstruction;
  wire         laneRequestSourceWire_3_bits_special = specialInstruction;
  wire         laneRequestSourceWire_4_bits_special = specialInstruction;
  wire         laneRequestSourceWire_5_bits_special = specialInstruction;
  wire         laneRequestSourceWire_6_bits_special = specialInstruction;
  wire         laneRequestSourceWire_7_bits_special = specialInstruction;
  wire         laneRequestSourceWire_8_bits_special = specialInstruction;
  wire         laneRequestSourceWire_9_bits_special = specialInstruction;
  wire         laneRequestSourceWire_10_bits_special = specialInstruction;
  wire         laneRequestSourceWire_11_bits_special = specialInstruction;
  wire         laneRequestSourceWire_12_bits_special = specialInstruction;
  wire         laneRequestSourceWire_13_bits_special = specialInstruction;
  wire         laneRequestSourceWire_14_bits_special = specialInstruction;
  wire         laneRequestSourceWire_15_bits_special = specialInstruction;
  wire [7:0]   dataInWritePipeVec_0;
  wire [7:0]   dataInWritePipeVec_1;
  wire [7:0]   dataInWritePipeVec_2;
  wire [7:0]   dataInWritePipeVec_3;
  wire [7:0]   dataInWritePipeVec_4;
  wire [7:0]   dataInWritePipeVec_5;
  wire [7:0]   dataInWritePipeVec_6;
  wire [7:0]   dataInWritePipeVec_7;
  wire [7:0]   dataInWritePipeVec_8;
  wire [7:0]   dataInWritePipeVec_9;
  wire [7:0]   dataInWritePipeVec_10;
  wire [7:0]   dataInWritePipeVec_11;
  wire [7:0]   dataInWritePipeVec_12;
  wire [7:0]   dataInWritePipeVec_13;
  wire [7:0]   dataInWritePipeVec_14;
  wire [7:0]   dataInWritePipeVec_15;
  wire [7:0]   dataInWritePipe =
    dataInWritePipeVec_0 | dataInWritePipeVec_1 | dataInWritePipeVec_2 | dataInWritePipeVec_3 | dataInWritePipeVec_4 | dataInWritePipeVec_5 | dataInWritePipeVec_6 | dataInWritePipeVec_7 | dataInWritePipeVec_8 | dataInWritePipeVec_9
    | dataInWritePipeVec_10 | dataInWritePipeVec_11 | dataInWritePipeVec_12 | dataInWritePipeVec_13 | dataInWritePipeVec_14 | dataInWritePipeVec_15;
  wire         gatherNeedRead = requestRegDequeue_valid & requestReg_bits_decodeResult_gather & ~requestReg_bits_decodeResult_vtype;
  reg  [2:0]   slots_0_record_instructionIndex;
  reg          slots_0_record_isLoadStore;
  reg          slots_0_record_maskType;
  reg          slots_0_state_wLast;
  reg          slots_0_state_idle;
  reg          slots_0_state_wMaskUnitLast;
  reg          slots_0_state_wVRFWrite;
  reg          slots_0_state_sCommit;
  reg          slots_0_endTag_0;
  reg          slots_0_endTag_1;
  reg          slots_0_endTag_2;
  reg          slots_0_endTag_3;
  reg          slots_0_endTag_4;
  reg          slots_0_endTag_5;
  reg          slots_0_endTag_6;
  reg          slots_0_endTag_7;
  reg          slots_0_endTag_8;
  reg          slots_0_endTag_9;
  reg          slots_0_endTag_10;
  reg          slots_0_endTag_11;
  reg          slots_0_endTag_12;
  reg          slots_0_endTag_13;
  reg          slots_0_endTag_14;
  reg          slots_0_endTag_15;
  reg          slots_0_endTag_16;
  reg          slots_0_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_lo = {slots_0_endTag_1, slots_0_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_hi = {slots_0_endTag_3, slots_0_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_lo = {slots_laneAndLSUFinish_lo_lo_hi, slots_laneAndLSUFinish_lo_lo_lo};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_lo = {slots_0_endTag_5, slots_0_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_hi = {slots_0_endTag_7, slots_0_endTag_6};
  wire [3:0]   slots_laneAndLSUFinish_lo_hi = {slots_laneAndLSUFinish_lo_hi_hi, slots_laneAndLSUFinish_lo_hi_lo};
  wire [7:0]   slots_laneAndLSUFinish_lo = {slots_laneAndLSUFinish_lo_hi, slots_laneAndLSUFinish_lo_lo};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_lo = {slots_0_endTag_9, slots_0_endTag_8};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_hi = {slots_0_endTag_11, slots_0_endTag_10};
  wire [3:0]   slots_laneAndLSUFinish_hi_lo = {slots_laneAndLSUFinish_hi_lo_hi, slots_laneAndLSUFinish_hi_lo_lo};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_lo = {slots_0_endTag_13, slots_0_endTag_12};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_hi = {slots_0_endTag_16, slots_0_endTag_15};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_hi = {slots_laneAndLSUFinish_hi_hi_hi_hi, slots_0_endTag_14};
  wire [4:0]   slots_laneAndLSUFinish_hi_hi = {slots_laneAndLSUFinish_hi_hi_hi, slots_laneAndLSUFinish_hi_hi_lo};
  wire [8:0]   slots_laneAndLSUFinish_hi = {slots_laneAndLSUFinish_hi_hi, slots_laneAndLSUFinish_hi_lo};
  wire         slots_laneAndLSUFinish = &{slots_laneAndLSUFinish_hi, slots_laneAndLSUFinish_lo};
  wire [7:0]   _GEN = {5'h0, slots_0_record_instructionIndex};
  wire         slots_v0WriteFinish = (8'h1 << _GEN & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished = |(8'h1 << _GEN & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_1 = 8'h1 << _GEN;
  wire         slots_vxsatUpdate = |(_slots_vxsatUpdate_T_1[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck = |(8'h1 << _GEN & dataInWritePipe);
  reg  [2:0]   slots_1_record_instructionIndex;
  reg          slots_1_record_isLoadStore;
  reg          slots_1_record_maskType;
  reg          slots_1_state_wLast;
  reg          slots_1_state_idle;
  reg          slots_1_state_wMaskUnitLast;
  reg          slots_1_state_wVRFWrite;
  reg          slots_1_state_sCommit;
  reg          slots_1_endTag_0;
  reg          slots_1_endTag_1;
  reg          slots_1_endTag_2;
  reg          slots_1_endTag_3;
  reg          slots_1_endTag_4;
  reg          slots_1_endTag_5;
  reg          slots_1_endTag_6;
  reg          slots_1_endTag_7;
  reg          slots_1_endTag_8;
  reg          slots_1_endTag_9;
  reg          slots_1_endTag_10;
  reg          slots_1_endTag_11;
  reg          slots_1_endTag_12;
  reg          slots_1_endTag_13;
  reg          slots_1_endTag_14;
  reg          slots_1_endTag_15;
  reg          slots_1_endTag_16;
  reg          slots_1_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_lo_1 = {slots_1_endTag_1, slots_1_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_hi_1 = {slots_1_endTag_3, slots_1_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_lo_1 = {slots_laneAndLSUFinish_lo_lo_hi_1, slots_laneAndLSUFinish_lo_lo_lo_1};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_lo_1 = {slots_1_endTag_5, slots_1_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_hi_1 = {slots_1_endTag_7, slots_1_endTag_6};
  wire [3:0]   slots_laneAndLSUFinish_lo_hi_1 = {slots_laneAndLSUFinish_lo_hi_hi_1, slots_laneAndLSUFinish_lo_hi_lo_1};
  wire [7:0]   slots_laneAndLSUFinish_lo_1 = {slots_laneAndLSUFinish_lo_hi_1, slots_laneAndLSUFinish_lo_lo_1};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_lo_1 = {slots_1_endTag_9, slots_1_endTag_8};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_hi_1 = {slots_1_endTag_11, slots_1_endTag_10};
  wire [3:0]   slots_laneAndLSUFinish_hi_lo_1 = {slots_laneAndLSUFinish_hi_lo_hi_1, slots_laneAndLSUFinish_hi_lo_lo_1};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_lo_1 = {slots_1_endTag_13, slots_1_endTag_12};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_hi_1 = {slots_1_endTag_16, slots_1_endTag_15};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_hi_1 = {slots_laneAndLSUFinish_hi_hi_hi_hi_1, slots_1_endTag_14};
  wire [4:0]   slots_laneAndLSUFinish_hi_hi_1 = {slots_laneAndLSUFinish_hi_hi_hi_1, slots_laneAndLSUFinish_hi_hi_lo_1};
  wire [8:0]   slots_laneAndLSUFinish_hi_1 = {slots_laneAndLSUFinish_hi_hi_1, slots_laneAndLSUFinish_hi_lo_1};
  wire         slots_laneAndLSUFinish_1 = &{slots_laneAndLSUFinish_hi_1, slots_laneAndLSUFinish_lo_1};
  wire [7:0]   _GEN_0 = {5'h0, slots_1_record_instructionIndex};
  wire         slots_v0WriteFinish_1 = (8'h1 << _GEN_0 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_1 = |(8'h1 << _GEN_0 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_4 = 8'h1 << _GEN_0;
  wire         slots_vxsatUpdate_1 = |(_slots_vxsatUpdate_T_4[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_1 = |(8'h1 << _GEN_0 & dataInWritePipe);
  reg  [2:0]   slots_2_record_instructionIndex;
  reg          slots_2_record_isLoadStore;
  reg          slots_2_record_maskType;
  reg          slots_2_state_wLast;
  reg          slots_2_state_idle;
  reg          slots_2_state_wMaskUnitLast;
  reg          slots_2_state_wVRFWrite;
  reg          slots_2_state_sCommit;
  reg          slots_2_endTag_0;
  reg          slots_2_endTag_1;
  reg          slots_2_endTag_2;
  reg          slots_2_endTag_3;
  reg          slots_2_endTag_4;
  reg          slots_2_endTag_5;
  reg          slots_2_endTag_6;
  reg          slots_2_endTag_7;
  reg          slots_2_endTag_8;
  reg          slots_2_endTag_9;
  reg          slots_2_endTag_10;
  reg          slots_2_endTag_11;
  reg          slots_2_endTag_12;
  reg          slots_2_endTag_13;
  reg          slots_2_endTag_14;
  reg          slots_2_endTag_15;
  reg          slots_2_endTag_16;
  reg          slots_2_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_lo_2 = {slots_2_endTag_1, slots_2_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_hi_2 = {slots_2_endTag_3, slots_2_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_lo_2 = {slots_laneAndLSUFinish_lo_lo_hi_2, slots_laneAndLSUFinish_lo_lo_lo_2};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_lo_2 = {slots_2_endTag_5, slots_2_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_hi_2 = {slots_2_endTag_7, slots_2_endTag_6};
  wire [3:0]   slots_laneAndLSUFinish_lo_hi_2 = {slots_laneAndLSUFinish_lo_hi_hi_2, slots_laneAndLSUFinish_lo_hi_lo_2};
  wire [7:0]   slots_laneAndLSUFinish_lo_2 = {slots_laneAndLSUFinish_lo_hi_2, slots_laneAndLSUFinish_lo_lo_2};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_lo_2 = {slots_2_endTag_9, slots_2_endTag_8};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_hi_2 = {slots_2_endTag_11, slots_2_endTag_10};
  wire [3:0]   slots_laneAndLSUFinish_hi_lo_2 = {slots_laneAndLSUFinish_hi_lo_hi_2, slots_laneAndLSUFinish_hi_lo_lo_2};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_lo_2 = {slots_2_endTag_13, slots_2_endTag_12};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_hi_2 = {slots_2_endTag_16, slots_2_endTag_15};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_hi_2 = {slots_laneAndLSUFinish_hi_hi_hi_hi_2, slots_2_endTag_14};
  wire [4:0]   slots_laneAndLSUFinish_hi_hi_2 = {slots_laneAndLSUFinish_hi_hi_hi_2, slots_laneAndLSUFinish_hi_hi_lo_2};
  wire [8:0]   slots_laneAndLSUFinish_hi_2 = {slots_laneAndLSUFinish_hi_hi_2, slots_laneAndLSUFinish_hi_lo_2};
  wire         slots_laneAndLSUFinish_2 = &{slots_laneAndLSUFinish_hi_2, slots_laneAndLSUFinish_lo_2};
  wire [7:0]   _GEN_1 = {5'h0, slots_2_record_instructionIndex};
  wire         slots_v0WriteFinish_2 = (8'h1 << _GEN_1 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_2 = |(8'h1 << _GEN_1 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_7 = 8'h1 << _GEN_1;
  wire         slots_vxsatUpdate_2 = |(_slots_vxsatUpdate_T_7[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_2 = |(8'h1 << _GEN_1 & dataInWritePipe);
  reg  [2:0]   slots_3_record_instructionIndex;
  reg          slots_3_record_isLoadStore;
  reg          slots_3_record_maskType;
  reg          slots_3_state_wLast;
  reg          slots_3_state_idle;
  reg          slots_3_state_wMaskUnitLast;
  reg          slots_3_state_wVRFWrite;
  reg          slots_3_state_sCommit;
  reg          slots_3_endTag_0;
  reg          slots_3_endTag_1;
  reg          slots_3_endTag_2;
  reg          slots_3_endTag_3;
  reg          slots_3_endTag_4;
  reg          slots_3_endTag_5;
  reg          slots_3_endTag_6;
  reg          slots_3_endTag_7;
  reg          slots_3_endTag_8;
  reg          slots_3_endTag_9;
  reg          slots_3_endTag_10;
  reg          slots_3_endTag_11;
  reg          slots_3_endTag_12;
  reg          slots_3_endTag_13;
  reg          slots_3_endTag_14;
  reg          slots_3_endTag_15;
  reg          slots_3_endTag_16;
  reg          slots_3_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_lo_3 = {slots_3_endTag_1, slots_3_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_hi_3 = {slots_3_endTag_3, slots_3_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_lo_3 = {slots_laneAndLSUFinish_lo_lo_hi_3, slots_laneAndLSUFinish_lo_lo_lo_3};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_lo_3 = {slots_3_endTag_5, slots_3_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_hi_3 = {slots_3_endTag_7, slots_3_endTag_6};
  wire [3:0]   slots_laneAndLSUFinish_lo_hi_3 = {slots_laneAndLSUFinish_lo_hi_hi_3, slots_laneAndLSUFinish_lo_hi_lo_3};
  wire [7:0]   slots_laneAndLSUFinish_lo_3 = {slots_laneAndLSUFinish_lo_hi_3, slots_laneAndLSUFinish_lo_lo_3};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_lo_3 = {slots_3_endTag_9, slots_3_endTag_8};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_hi_3 = {slots_3_endTag_11, slots_3_endTag_10};
  wire [3:0]   slots_laneAndLSUFinish_hi_lo_3 = {slots_laneAndLSUFinish_hi_lo_hi_3, slots_laneAndLSUFinish_hi_lo_lo_3};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_lo_3 = {slots_3_endTag_13, slots_3_endTag_12};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_hi_3 = {slots_3_endTag_16, slots_3_endTag_15};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_hi_3 = {slots_laneAndLSUFinish_hi_hi_hi_hi_3, slots_3_endTag_14};
  wire [4:0]   slots_laneAndLSUFinish_hi_hi_3 = {slots_laneAndLSUFinish_hi_hi_hi_3, slots_laneAndLSUFinish_hi_hi_lo_3};
  wire [8:0]   slots_laneAndLSUFinish_hi_3 = {slots_laneAndLSUFinish_hi_hi_3, slots_laneAndLSUFinish_hi_lo_3};
  wire         slots_laneAndLSUFinish_3 = &{slots_laneAndLSUFinish_hi_3, slots_laneAndLSUFinish_lo_3};
  wire [7:0]   _GEN_2 = {5'h0, slots_3_record_instructionIndex};
  wire         slots_v0WriteFinish_3 = (8'h1 << _GEN_2 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_3 = |(8'h1 << _GEN_2 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_10 = 8'h1 << _GEN_2;
  wire         slots_vxsatUpdate_3 = |(_slots_vxsatUpdate_T_10[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_3 = |(8'h1 << _GEN_2 & dataInWritePipe);
  reg          slots_writeRD;
  reg          slots_float;
  wire         retire_rd_bits_isFp_0 = slots_float;
  reg  [4:0]   slots_vd;
  wire [4:0]   retire_rd_bits_rdAddress_0 = slots_vd;
  wire         lastSlotCommit;
  wire         retire_rd_valid_0 = lastSlotCommit & slots_writeRD;
  wire         tokenCheck;
  wire [2:0]   validSource_bits_instructionIndex = laneRequestSourceWire_0_bits_instructionIndex;
  wire         validSource_bits_decodeResult_orderReduce = laneRequestSourceWire_0_bits_decodeResult_orderReduce;
  wire         validSource_bits_decodeResult_floatMul = laneRequestSourceWire_0_bits_decodeResult_floatMul;
  wire [1:0]   validSource_bits_decodeResult_fpExecutionType = laneRequestSourceWire_0_bits_decodeResult_fpExecutionType;
  wire         validSource_bits_decodeResult_float = laneRequestSourceWire_0_bits_decodeResult_float;
  wire         validSource_bits_decodeResult_specialSlot = laneRequestSourceWire_0_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_bits_decodeResult_topUop = laneRequestSourceWire_0_bits_decodeResult_topUop;
  wire         validSource_bits_decodeResult_popCount = laneRequestSourceWire_0_bits_decodeResult_popCount;
  wire         validSource_bits_decodeResult_ffo = laneRequestSourceWire_0_bits_decodeResult_ffo;
  wire         validSource_bits_decodeResult_average = laneRequestSourceWire_0_bits_decodeResult_average;
  wire         validSource_bits_decodeResult_reverse = laneRequestSourceWire_0_bits_decodeResult_reverse;
  wire         validSource_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_0_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_bits_decodeResult_scheduler = laneRequestSourceWire_0_bits_decodeResult_scheduler;
  wire         validSource_bits_decodeResult_sReadVD = laneRequestSourceWire_0_bits_decodeResult_sReadVD;
  wire         validSource_bits_decodeResult_vtype = laneRequestSourceWire_0_bits_decodeResult_vtype;
  wire         validSource_bits_decodeResult_sWrite = laneRequestSourceWire_0_bits_decodeResult_sWrite;
  wire         validSource_bits_decodeResult_crossRead = laneRequestSourceWire_0_bits_decodeResult_crossRead;
  wire         validSource_bits_decodeResult_crossWrite = laneRequestSourceWire_0_bits_decodeResult_crossWrite;
  wire         validSource_bits_decodeResult_maskUnit = laneRequestSourceWire_0_bits_decodeResult_maskUnit;
  wire         validSource_bits_decodeResult_special = laneRequestSourceWire_0_bits_decodeResult_special;
  wire         validSource_bits_decodeResult_saturate = laneRequestSourceWire_0_bits_decodeResult_saturate;
  wire         validSource_bits_decodeResult_vwmacc = laneRequestSourceWire_0_bits_decodeResult_vwmacc;
  wire         validSource_bits_decodeResult_readOnly = laneRequestSourceWire_0_bits_decodeResult_readOnly;
  wire         validSource_bits_decodeResult_maskSource = laneRequestSourceWire_0_bits_decodeResult_maskSource;
  wire         validSource_bits_decodeResult_maskDestination = laneRequestSourceWire_0_bits_decodeResult_maskDestination;
  wire         validSource_bits_decodeResult_maskLogic = laneRequestSourceWire_0_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_bits_decodeResult_uop = laneRequestSourceWire_0_bits_decodeResult_uop;
  wire         validSource_bits_decodeResult_iota = laneRequestSourceWire_0_bits_decodeResult_iota;
  wire         validSource_bits_decodeResult_mv = laneRequestSourceWire_0_bits_decodeResult_mv;
  wire         validSource_bits_decodeResult_extend = laneRequestSourceWire_0_bits_decodeResult_extend;
  wire         validSource_bits_decodeResult_unOrderWrite = laneRequestSourceWire_0_bits_decodeResult_unOrderWrite;
  wire         validSource_bits_decodeResult_compress = laneRequestSourceWire_0_bits_decodeResult_compress;
  wire         validSource_bits_decodeResult_gather16 = laneRequestSourceWire_0_bits_decodeResult_gather16;
  wire         validSource_bits_decodeResult_gather = laneRequestSourceWire_0_bits_decodeResult_gather;
  wire         validSource_bits_decodeResult_slid = laneRequestSourceWire_0_bits_decodeResult_slid;
  wire         validSource_bits_decodeResult_targetRd = laneRequestSourceWire_0_bits_decodeResult_targetRd;
  wire         validSource_bits_decodeResult_widenReduce = laneRequestSourceWire_0_bits_decodeResult_widenReduce;
  wire         validSource_bits_decodeResult_red = laneRequestSourceWire_0_bits_decodeResult_red;
  wire         validSource_bits_decodeResult_nr = laneRequestSourceWire_0_bits_decodeResult_nr;
  wire         validSource_bits_decodeResult_itype = laneRequestSourceWire_0_bits_decodeResult_itype;
  wire         validSource_bits_decodeResult_unsigned1 = laneRequestSourceWire_0_bits_decodeResult_unsigned1;
  wire         validSource_bits_decodeResult_unsigned0 = laneRequestSourceWire_0_bits_decodeResult_unsigned0;
  wire         validSource_bits_decodeResult_other = laneRequestSourceWire_0_bits_decodeResult_other;
  wire         validSource_bits_decodeResult_multiCycle = laneRequestSourceWire_0_bits_decodeResult_multiCycle;
  wire         validSource_bits_decodeResult_divider = laneRequestSourceWire_0_bits_decodeResult_divider;
  wire         validSource_bits_decodeResult_multiplier = laneRequestSourceWire_0_bits_decodeResult_multiplier;
  wire         validSource_bits_decodeResult_shift = laneRequestSourceWire_0_bits_decodeResult_shift;
  wire         validSource_bits_decodeResult_adder = laneRequestSourceWire_0_bits_decodeResult_adder;
  wire         validSource_bits_decodeResult_logic = laneRequestSourceWire_0_bits_decodeResult_logic;
  wire         validSource_bits_loadStore = laneRequestSourceWire_0_bits_loadStore;
  wire         validSource_bits_issueInst = laneRequestSourceWire_0_bits_issueInst;
  wire         validSource_bits_store = laneRequestSourceWire_0_bits_store;
  wire         validSource_bits_special = laneRequestSourceWire_0_bits_special;
  wire         validSource_bits_lsWholeReg = laneRequestSourceWire_0_bits_lsWholeReg;
  wire [4:0]   validSource_bits_vs1 = laneRequestSourceWire_0_bits_vs1;
  wire [4:0]   validSource_bits_vs2 = laneRequestSourceWire_0_bits_vs2;
  wire [4:0]   validSource_bits_vd = laneRequestSourceWire_0_bits_vd;
  wire [1:0]   validSource_bits_loadStoreEEW = laneRequestSourceWire_0_bits_loadStoreEEW;
  wire         validSource_bits_mask = laneRequestSourceWire_0_bits_mask;
  wire [2:0]   validSource_bits_segment = laneRequestSourceWire_0_bits_segment;
  wire [31:0]  source1Select;
  wire [31:0]  validSource_bits_readFromScalar = laneRequestSourceWire_0_bits_readFromScalar;
  wire [11:0]  validSource_bits_csrInterface_vl = laneRequestSourceWire_0_bits_csrInterface_vl;
  wire [11:0]  validSource_bits_csrInterface_vStart = laneRequestSourceWire_0_bits_csrInterface_vStart;
  wire [2:0]   validSource_bits_csrInterface_vlmul = laneRequestSourceWire_0_bits_csrInterface_vlmul;
  wire [1:0]   validSource_bits_csrInterface_vSew = laneRequestSourceWire_0_bits_csrInterface_vSew;
  wire [1:0]   validSource_bits_csrInterface_vxrm = laneRequestSourceWire_0_bits_csrInterface_vxrm;
  wire         validSource_bits_csrInterface_vta = laneRequestSourceWire_0_bits_csrInterface_vta;
  wire         validSource_bits_csrInterface_vma = laneRequestSourceWire_0_bits_csrInterface_vma;
  wire         tokenCheck_1;
  wire [2:0]   validSource_1_bits_instructionIndex = laneRequestSourceWire_1_bits_instructionIndex;
  wire         validSource_1_bits_decodeResult_orderReduce = laneRequestSourceWire_1_bits_decodeResult_orderReduce;
  wire         validSource_1_bits_decodeResult_floatMul = laneRequestSourceWire_1_bits_decodeResult_floatMul;
  wire [1:0]   validSource_1_bits_decodeResult_fpExecutionType = laneRequestSourceWire_1_bits_decodeResult_fpExecutionType;
  wire         validSource_1_bits_decodeResult_float = laneRequestSourceWire_1_bits_decodeResult_float;
  wire         validSource_1_bits_decodeResult_specialSlot = laneRequestSourceWire_1_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_1_bits_decodeResult_topUop = laneRequestSourceWire_1_bits_decodeResult_topUop;
  wire         validSource_1_bits_decodeResult_popCount = laneRequestSourceWire_1_bits_decodeResult_popCount;
  wire         validSource_1_bits_decodeResult_ffo = laneRequestSourceWire_1_bits_decodeResult_ffo;
  wire         validSource_1_bits_decodeResult_average = laneRequestSourceWire_1_bits_decodeResult_average;
  wire         validSource_1_bits_decodeResult_reverse = laneRequestSourceWire_1_bits_decodeResult_reverse;
  wire         validSource_1_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_1_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_1_bits_decodeResult_scheduler = laneRequestSourceWire_1_bits_decodeResult_scheduler;
  wire         validSource_1_bits_decodeResult_sReadVD = laneRequestSourceWire_1_bits_decodeResult_sReadVD;
  wire         validSource_1_bits_decodeResult_vtype = laneRequestSourceWire_1_bits_decodeResult_vtype;
  wire         validSource_1_bits_decodeResult_sWrite = laneRequestSourceWire_1_bits_decodeResult_sWrite;
  wire         validSource_1_bits_decodeResult_crossRead = laneRequestSourceWire_1_bits_decodeResult_crossRead;
  wire         validSource_1_bits_decodeResult_crossWrite = laneRequestSourceWire_1_bits_decodeResult_crossWrite;
  wire         validSource_1_bits_decodeResult_maskUnit = laneRequestSourceWire_1_bits_decodeResult_maskUnit;
  wire         validSource_1_bits_decodeResult_special = laneRequestSourceWire_1_bits_decodeResult_special;
  wire         validSource_1_bits_decodeResult_saturate = laneRequestSourceWire_1_bits_decodeResult_saturate;
  wire         validSource_1_bits_decodeResult_vwmacc = laneRequestSourceWire_1_bits_decodeResult_vwmacc;
  wire         validSource_1_bits_decodeResult_readOnly = laneRequestSourceWire_1_bits_decodeResult_readOnly;
  wire         validSource_1_bits_decodeResult_maskSource = laneRequestSourceWire_1_bits_decodeResult_maskSource;
  wire         validSource_1_bits_decodeResult_maskDestination = laneRequestSourceWire_1_bits_decodeResult_maskDestination;
  wire         validSource_1_bits_decodeResult_maskLogic = laneRequestSourceWire_1_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_1_bits_decodeResult_uop = laneRequestSourceWire_1_bits_decodeResult_uop;
  wire         validSource_1_bits_decodeResult_iota = laneRequestSourceWire_1_bits_decodeResult_iota;
  wire         validSource_1_bits_decodeResult_mv = laneRequestSourceWire_1_bits_decodeResult_mv;
  wire         validSource_1_bits_decodeResult_extend = laneRequestSourceWire_1_bits_decodeResult_extend;
  wire         validSource_1_bits_decodeResult_unOrderWrite = laneRequestSourceWire_1_bits_decodeResult_unOrderWrite;
  wire         validSource_1_bits_decodeResult_compress = laneRequestSourceWire_1_bits_decodeResult_compress;
  wire         validSource_1_bits_decodeResult_gather16 = laneRequestSourceWire_1_bits_decodeResult_gather16;
  wire         validSource_1_bits_decodeResult_gather = laneRequestSourceWire_1_bits_decodeResult_gather;
  wire         validSource_1_bits_decodeResult_slid = laneRequestSourceWire_1_bits_decodeResult_slid;
  wire         validSource_1_bits_decodeResult_targetRd = laneRequestSourceWire_1_bits_decodeResult_targetRd;
  wire         validSource_1_bits_decodeResult_widenReduce = laneRequestSourceWire_1_bits_decodeResult_widenReduce;
  wire         validSource_1_bits_decodeResult_red = laneRequestSourceWire_1_bits_decodeResult_red;
  wire         validSource_1_bits_decodeResult_nr = laneRequestSourceWire_1_bits_decodeResult_nr;
  wire         validSource_1_bits_decodeResult_itype = laneRequestSourceWire_1_bits_decodeResult_itype;
  wire         validSource_1_bits_decodeResult_unsigned1 = laneRequestSourceWire_1_bits_decodeResult_unsigned1;
  wire         validSource_1_bits_decodeResult_unsigned0 = laneRequestSourceWire_1_bits_decodeResult_unsigned0;
  wire         validSource_1_bits_decodeResult_other = laneRequestSourceWire_1_bits_decodeResult_other;
  wire         validSource_1_bits_decodeResult_multiCycle = laneRequestSourceWire_1_bits_decodeResult_multiCycle;
  wire         validSource_1_bits_decodeResult_divider = laneRequestSourceWire_1_bits_decodeResult_divider;
  wire         validSource_1_bits_decodeResult_multiplier = laneRequestSourceWire_1_bits_decodeResult_multiplier;
  wire         validSource_1_bits_decodeResult_shift = laneRequestSourceWire_1_bits_decodeResult_shift;
  wire         validSource_1_bits_decodeResult_adder = laneRequestSourceWire_1_bits_decodeResult_adder;
  wire         validSource_1_bits_decodeResult_logic = laneRequestSourceWire_1_bits_decodeResult_logic;
  wire         validSource_1_bits_loadStore = laneRequestSourceWire_1_bits_loadStore;
  wire         validSource_1_bits_issueInst = laneRequestSourceWire_1_bits_issueInst;
  wire         validSource_1_bits_store = laneRequestSourceWire_1_bits_store;
  wire         validSource_1_bits_special = laneRequestSourceWire_1_bits_special;
  wire         validSource_1_bits_lsWholeReg = laneRequestSourceWire_1_bits_lsWholeReg;
  wire [4:0]   validSource_1_bits_vs1 = laneRequestSourceWire_1_bits_vs1;
  wire [4:0]   validSource_1_bits_vs2 = laneRequestSourceWire_1_bits_vs2;
  wire [4:0]   validSource_1_bits_vd = laneRequestSourceWire_1_bits_vd;
  wire [1:0]   validSource_1_bits_loadStoreEEW = laneRequestSourceWire_1_bits_loadStoreEEW;
  wire         validSource_1_bits_mask = laneRequestSourceWire_1_bits_mask;
  wire [2:0]   validSource_1_bits_segment = laneRequestSourceWire_1_bits_segment;
  wire [31:0]  validSource_1_bits_readFromScalar = laneRequestSourceWire_1_bits_readFromScalar;
  wire [11:0]  validSource_1_bits_csrInterface_vl = laneRequestSourceWire_1_bits_csrInterface_vl;
  wire [11:0]  validSource_1_bits_csrInterface_vStart = laneRequestSourceWire_1_bits_csrInterface_vStart;
  wire [2:0]   validSource_1_bits_csrInterface_vlmul = laneRequestSourceWire_1_bits_csrInterface_vlmul;
  wire [1:0]   validSource_1_bits_csrInterface_vSew = laneRequestSourceWire_1_bits_csrInterface_vSew;
  wire [1:0]   validSource_1_bits_csrInterface_vxrm = laneRequestSourceWire_1_bits_csrInterface_vxrm;
  wire         validSource_1_bits_csrInterface_vta = laneRequestSourceWire_1_bits_csrInterface_vta;
  wire         validSource_1_bits_csrInterface_vma = laneRequestSourceWire_1_bits_csrInterface_vma;
  wire         tokenCheck_2;
  wire [2:0]   validSource_2_bits_instructionIndex = laneRequestSourceWire_2_bits_instructionIndex;
  wire         validSource_2_bits_decodeResult_orderReduce = laneRequestSourceWire_2_bits_decodeResult_orderReduce;
  wire         validSource_2_bits_decodeResult_floatMul = laneRequestSourceWire_2_bits_decodeResult_floatMul;
  wire [1:0]   validSource_2_bits_decodeResult_fpExecutionType = laneRequestSourceWire_2_bits_decodeResult_fpExecutionType;
  wire         validSource_2_bits_decodeResult_float = laneRequestSourceWire_2_bits_decodeResult_float;
  wire         validSource_2_bits_decodeResult_specialSlot = laneRequestSourceWire_2_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_2_bits_decodeResult_topUop = laneRequestSourceWire_2_bits_decodeResult_topUop;
  wire         validSource_2_bits_decodeResult_popCount = laneRequestSourceWire_2_bits_decodeResult_popCount;
  wire         validSource_2_bits_decodeResult_ffo = laneRequestSourceWire_2_bits_decodeResult_ffo;
  wire         validSource_2_bits_decodeResult_average = laneRequestSourceWire_2_bits_decodeResult_average;
  wire         validSource_2_bits_decodeResult_reverse = laneRequestSourceWire_2_bits_decodeResult_reverse;
  wire         validSource_2_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_2_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_2_bits_decodeResult_scheduler = laneRequestSourceWire_2_bits_decodeResult_scheduler;
  wire         validSource_2_bits_decodeResult_sReadVD = laneRequestSourceWire_2_bits_decodeResult_sReadVD;
  wire         validSource_2_bits_decodeResult_vtype = laneRequestSourceWire_2_bits_decodeResult_vtype;
  wire         validSource_2_bits_decodeResult_sWrite = laneRequestSourceWire_2_bits_decodeResult_sWrite;
  wire         validSource_2_bits_decodeResult_crossRead = laneRequestSourceWire_2_bits_decodeResult_crossRead;
  wire         validSource_2_bits_decodeResult_crossWrite = laneRequestSourceWire_2_bits_decodeResult_crossWrite;
  wire         validSource_2_bits_decodeResult_maskUnit = laneRequestSourceWire_2_bits_decodeResult_maskUnit;
  wire         validSource_2_bits_decodeResult_special = laneRequestSourceWire_2_bits_decodeResult_special;
  wire         validSource_2_bits_decodeResult_saturate = laneRequestSourceWire_2_bits_decodeResult_saturate;
  wire         validSource_2_bits_decodeResult_vwmacc = laneRequestSourceWire_2_bits_decodeResult_vwmacc;
  wire         validSource_2_bits_decodeResult_readOnly = laneRequestSourceWire_2_bits_decodeResult_readOnly;
  wire         validSource_2_bits_decodeResult_maskSource = laneRequestSourceWire_2_bits_decodeResult_maskSource;
  wire         validSource_2_bits_decodeResult_maskDestination = laneRequestSourceWire_2_bits_decodeResult_maskDestination;
  wire         validSource_2_bits_decodeResult_maskLogic = laneRequestSourceWire_2_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_2_bits_decodeResult_uop = laneRequestSourceWire_2_bits_decodeResult_uop;
  wire         validSource_2_bits_decodeResult_iota = laneRequestSourceWire_2_bits_decodeResult_iota;
  wire         validSource_2_bits_decodeResult_mv = laneRequestSourceWire_2_bits_decodeResult_mv;
  wire         validSource_2_bits_decodeResult_extend = laneRequestSourceWire_2_bits_decodeResult_extend;
  wire         validSource_2_bits_decodeResult_unOrderWrite = laneRequestSourceWire_2_bits_decodeResult_unOrderWrite;
  wire         validSource_2_bits_decodeResult_compress = laneRequestSourceWire_2_bits_decodeResult_compress;
  wire         validSource_2_bits_decodeResult_gather16 = laneRequestSourceWire_2_bits_decodeResult_gather16;
  wire         validSource_2_bits_decodeResult_gather = laneRequestSourceWire_2_bits_decodeResult_gather;
  wire         validSource_2_bits_decodeResult_slid = laneRequestSourceWire_2_bits_decodeResult_slid;
  wire         validSource_2_bits_decodeResult_targetRd = laneRequestSourceWire_2_bits_decodeResult_targetRd;
  wire         validSource_2_bits_decodeResult_widenReduce = laneRequestSourceWire_2_bits_decodeResult_widenReduce;
  wire         validSource_2_bits_decodeResult_red = laneRequestSourceWire_2_bits_decodeResult_red;
  wire         validSource_2_bits_decodeResult_nr = laneRequestSourceWire_2_bits_decodeResult_nr;
  wire         validSource_2_bits_decodeResult_itype = laneRequestSourceWire_2_bits_decodeResult_itype;
  wire         validSource_2_bits_decodeResult_unsigned1 = laneRequestSourceWire_2_bits_decodeResult_unsigned1;
  wire         validSource_2_bits_decodeResult_unsigned0 = laneRequestSourceWire_2_bits_decodeResult_unsigned0;
  wire         validSource_2_bits_decodeResult_other = laneRequestSourceWire_2_bits_decodeResult_other;
  wire         validSource_2_bits_decodeResult_multiCycle = laneRequestSourceWire_2_bits_decodeResult_multiCycle;
  wire         validSource_2_bits_decodeResult_divider = laneRequestSourceWire_2_bits_decodeResult_divider;
  wire         validSource_2_bits_decodeResult_multiplier = laneRequestSourceWire_2_bits_decodeResult_multiplier;
  wire         validSource_2_bits_decodeResult_shift = laneRequestSourceWire_2_bits_decodeResult_shift;
  wire         validSource_2_bits_decodeResult_adder = laneRequestSourceWire_2_bits_decodeResult_adder;
  wire         validSource_2_bits_decodeResult_logic = laneRequestSourceWire_2_bits_decodeResult_logic;
  wire         validSource_2_bits_loadStore = laneRequestSourceWire_2_bits_loadStore;
  wire         validSource_2_bits_issueInst = laneRequestSourceWire_2_bits_issueInst;
  wire         validSource_2_bits_store = laneRequestSourceWire_2_bits_store;
  wire         validSource_2_bits_special = laneRequestSourceWire_2_bits_special;
  wire         validSource_2_bits_lsWholeReg = laneRequestSourceWire_2_bits_lsWholeReg;
  wire [4:0]   validSource_2_bits_vs1 = laneRequestSourceWire_2_bits_vs1;
  wire [4:0]   validSource_2_bits_vs2 = laneRequestSourceWire_2_bits_vs2;
  wire [4:0]   validSource_2_bits_vd = laneRequestSourceWire_2_bits_vd;
  wire [1:0]   validSource_2_bits_loadStoreEEW = laneRequestSourceWire_2_bits_loadStoreEEW;
  wire         validSource_2_bits_mask = laneRequestSourceWire_2_bits_mask;
  wire [2:0]   validSource_2_bits_segment = laneRequestSourceWire_2_bits_segment;
  wire [31:0]  validSource_2_bits_readFromScalar = laneRequestSourceWire_2_bits_readFromScalar;
  wire [11:0]  validSource_2_bits_csrInterface_vl = laneRequestSourceWire_2_bits_csrInterface_vl;
  wire [11:0]  validSource_2_bits_csrInterface_vStart = laneRequestSourceWire_2_bits_csrInterface_vStart;
  wire [2:0]   validSource_2_bits_csrInterface_vlmul = laneRequestSourceWire_2_bits_csrInterface_vlmul;
  wire [1:0]   validSource_2_bits_csrInterface_vSew = laneRequestSourceWire_2_bits_csrInterface_vSew;
  wire [1:0]   validSource_2_bits_csrInterface_vxrm = laneRequestSourceWire_2_bits_csrInterface_vxrm;
  wire         validSource_2_bits_csrInterface_vta = laneRequestSourceWire_2_bits_csrInterface_vta;
  wire         validSource_2_bits_csrInterface_vma = laneRequestSourceWire_2_bits_csrInterface_vma;
  wire         tokenCheck_3;
  wire [2:0]   validSource_3_bits_instructionIndex = laneRequestSourceWire_3_bits_instructionIndex;
  wire         validSource_3_bits_decodeResult_orderReduce = laneRequestSourceWire_3_bits_decodeResult_orderReduce;
  wire         validSource_3_bits_decodeResult_floatMul = laneRequestSourceWire_3_bits_decodeResult_floatMul;
  wire [1:0]   validSource_3_bits_decodeResult_fpExecutionType = laneRequestSourceWire_3_bits_decodeResult_fpExecutionType;
  wire         validSource_3_bits_decodeResult_float = laneRequestSourceWire_3_bits_decodeResult_float;
  wire         validSource_3_bits_decodeResult_specialSlot = laneRequestSourceWire_3_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_3_bits_decodeResult_topUop = laneRequestSourceWire_3_bits_decodeResult_topUop;
  wire         validSource_3_bits_decodeResult_popCount = laneRequestSourceWire_3_bits_decodeResult_popCount;
  wire         validSource_3_bits_decodeResult_ffo = laneRequestSourceWire_3_bits_decodeResult_ffo;
  wire         validSource_3_bits_decodeResult_average = laneRequestSourceWire_3_bits_decodeResult_average;
  wire         validSource_3_bits_decodeResult_reverse = laneRequestSourceWire_3_bits_decodeResult_reverse;
  wire         validSource_3_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_3_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_3_bits_decodeResult_scheduler = laneRequestSourceWire_3_bits_decodeResult_scheduler;
  wire         validSource_3_bits_decodeResult_sReadVD = laneRequestSourceWire_3_bits_decodeResult_sReadVD;
  wire         validSource_3_bits_decodeResult_vtype = laneRequestSourceWire_3_bits_decodeResult_vtype;
  wire         validSource_3_bits_decodeResult_sWrite = laneRequestSourceWire_3_bits_decodeResult_sWrite;
  wire         validSource_3_bits_decodeResult_crossRead = laneRequestSourceWire_3_bits_decodeResult_crossRead;
  wire         validSource_3_bits_decodeResult_crossWrite = laneRequestSourceWire_3_bits_decodeResult_crossWrite;
  wire         validSource_3_bits_decodeResult_maskUnit = laneRequestSourceWire_3_bits_decodeResult_maskUnit;
  wire         validSource_3_bits_decodeResult_special = laneRequestSourceWire_3_bits_decodeResult_special;
  wire         validSource_3_bits_decodeResult_saturate = laneRequestSourceWire_3_bits_decodeResult_saturate;
  wire         validSource_3_bits_decodeResult_vwmacc = laneRequestSourceWire_3_bits_decodeResult_vwmacc;
  wire         validSource_3_bits_decodeResult_readOnly = laneRequestSourceWire_3_bits_decodeResult_readOnly;
  wire         validSource_3_bits_decodeResult_maskSource = laneRequestSourceWire_3_bits_decodeResult_maskSource;
  wire         validSource_3_bits_decodeResult_maskDestination = laneRequestSourceWire_3_bits_decodeResult_maskDestination;
  wire         validSource_3_bits_decodeResult_maskLogic = laneRequestSourceWire_3_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_3_bits_decodeResult_uop = laneRequestSourceWire_3_bits_decodeResult_uop;
  wire         validSource_3_bits_decodeResult_iota = laneRequestSourceWire_3_bits_decodeResult_iota;
  wire         validSource_3_bits_decodeResult_mv = laneRequestSourceWire_3_bits_decodeResult_mv;
  wire         validSource_3_bits_decodeResult_extend = laneRequestSourceWire_3_bits_decodeResult_extend;
  wire         validSource_3_bits_decodeResult_unOrderWrite = laneRequestSourceWire_3_bits_decodeResult_unOrderWrite;
  wire         validSource_3_bits_decodeResult_compress = laneRequestSourceWire_3_bits_decodeResult_compress;
  wire         validSource_3_bits_decodeResult_gather16 = laneRequestSourceWire_3_bits_decodeResult_gather16;
  wire         validSource_3_bits_decodeResult_gather = laneRequestSourceWire_3_bits_decodeResult_gather;
  wire         validSource_3_bits_decodeResult_slid = laneRequestSourceWire_3_bits_decodeResult_slid;
  wire         validSource_3_bits_decodeResult_targetRd = laneRequestSourceWire_3_bits_decodeResult_targetRd;
  wire         validSource_3_bits_decodeResult_widenReduce = laneRequestSourceWire_3_bits_decodeResult_widenReduce;
  wire         validSource_3_bits_decodeResult_red = laneRequestSourceWire_3_bits_decodeResult_red;
  wire         validSource_3_bits_decodeResult_nr = laneRequestSourceWire_3_bits_decodeResult_nr;
  wire         validSource_3_bits_decodeResult_itype = laneRequestSourceWire_3_bits_decodeResult_itype;
  wire         validSource_3_bits_decodeResult_unsigned1 = laneRequestSourceWire_3_bits_decodeResult_unsigned1;
  wire         validSource_3_bits_decodeResult_unsigned0 = laneRequestSourceWire_3_bits_decodeResult_unsigned0;
  wire         validSource_3_bits_decodeResult_other = laneRequestSourceWire_3_bits_decodeResult_other;
  wire         validSource_3_bits_decodeResult_multiCycle = laneRequestSourceWire_3_bits_decodeResult_multiCycle;
  wire         validSource_3_bits_decodeResult_divider = laneRequestSourceWire_3_bits_decodeResult_divider;
  wire         validSource_3_bits_decodeResult_multiplier = laneRequestSourceWire_3_bits_decodeResult_multiplier;
  wire         validSource_3_bits_decodeResult_shift = laneRequestSourceWire_3_bits_decodeResult_shift;
  wire         validSource_3_bits_decodeResult_adder = laneRequestSourceWire_3_bits_decodeResult_adder;
  wire         validSource_3_bits_decodeResult_logic = laneRequestSourceWire_3_bits_decodeResult_logic;
  wire         validSource_3_bits_loadStore = laneRequestSourceWire_3_bits_loadStore;
  wire         validSource_3_bits_issueInst = laneRequestSourceWire_3_bits_issueInst;
  wire         validSource_3_bits_store = laneRequestSourceWire_3_bits_store;
  wire         validSource_3_bits_special = laneRequestSourceWire_3_bits_special;
  wire         validSource_3_bits_lsWholeReg = laneRequestSourceWire_3_bits_lsWholeReg;
  wire [4:0]   validSource_3_bits_vs1 = laneRequestSourceWire_3_bits_vs1;
  wire [4:0]   validSource_3_bits_vs2 = laneRequestSourceWire_3_bits_vs2;
  wire [4:0]   validSource_3_bits_vd = laneRequestSourceWire_3_bits_vd;
  wire [1:0]   validSource_3_bits_loadStoreEEW = laneRequestSourceWire_3_bits_loadStoreEEW;
  wire         validSource_3_bits_mask = laneRequestSourceWire_3_bits_mask;
  wire [2:0]   validSource_3_bits_segment = laneRequestSourceWire_3_bits_segment;
  wire [31:0]  validSource_3_bits_readFromScalar = laneRequestSourceWire_3_bits_readFromScalar;
  wire [11:0]  validSource_3_bits_csrInterface_vl = laneRequestSourceWire_3_bits_csrInterface_vl;
  wire [11:0]  validSource_3_bits_csrInterface_vStart = laneRequestSourceWire_3_bits_csrInterface_vStart;
  wire [2:0]   validSource_3_bits_csrInterface_vlmul = laneRequestSourceWire_3_bits_csrInterface_vlmul;
  wire [1:0]   validSource_3_bits_csrInterface_vSew = laneRequestSourceWire_3_bits_csrInterface_vSew;
  wire [1:0]   validSource_3_bits_csrInterface_vxrm = laneRequestSourceWire_3_bits_csrInterface_vxrm;
  wire         validSource_3_bits_csrInterface_vta = laneRequestSourceWire_3_bits_csrInterface_vta;
  wire         validSource_3_bits_csrInterface_vma = laneRequestSourceWire_3_bits_csrInterface_vma;
  wire         tokenCheck_4;
  wire [2:0]   validSource_4_bits_instructionIndex = laneRequestSourceWire_4_bits_instructionIndex;
  wire         validSource_4_bits_decodeResult_orderReduce = laneRequestSourceWire_4_bits_decodeResult_orderReduce;
  wire         validSource_4_bits_decodeResult_floatMul = laneRequestSourceWire_4_bits_decodeResult_floatMul;
  wire [1:0]   validSource_4_bits_decodeResult_fpExecutionType = laneRequestSourceWire_4_bits_decodeResult_fpExecutionType;
  wire         validSource_4_bits_decodeResult_float = laneRequestSourceWire_4_bits_decodeResult_float;
  wire         validSource_4_bits_decodeResult_specialSlot = laneRequestSourceWire_4_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_4_bits_decodeResult_topUop = laneRequestSourceWire_4_bits_decodeResult_topUop;
  wire         validSource_4_bits_decodeResult_popCount = laneRequestSourceWire_4_bits_decodeResult_popCount;
  wire         validSource_4_bits_decodeResult_ffo = laneRequestSourceWire_4_bits_decodeResult_ffo;
  wire         validSource_4_bits_decodeResult_average = laneRequestSourceWire_4_bits_decodeResult_average;
  wire         validSource_4_bits_decodeResult_reverse = laneRequestSourceWire_4_bits_decodeResult_reverse;
  wire         validSource_4_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_4_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_4_bits_decodeResult_scheduler = laneRequestSourceWire_4_bits_decodeResult_scheduler;
  wire         validSource_4_bits_decodeResult_sReadVD = laneRequestSourceWire_4_bits_decodeResult_sReadVD;
  wire         validSource_4_bits_decodeResult_vtype = laneRequestSourceWire_4_bits_decodeResult_vtype;
  wire         validSource_4_bits_decodeResult_sWrite = laneRequestSourceWire_4_bits_decodeResult_sWrite;
  wire         validSource_4_bits_decodeResult_crossRead = laneRequestSourceWire_4_bits_decodeResult_crossRead;
  wire         validSource_4_bits_decodeResult_crossWrite = laneRequestSourceWire_4_bits_decodeResult_crossWrite;
  wire         validSource_4_bits_decodeResult_maskUnit = laneRequestSourceWire_4_bits_decodeResult_maskUnit;
  wire         validSource_4_bits_decodeResult_special = laneRequestSourceWire_4_bits_decodeResult_special;
  wire         validSource_4_bits_decodeResult_saturate = laneRequestSourceWire_4_bits_decodeResult_saturate;
  wire         validSource_4_bits_decodeResult_vwmacc = laneRequestSourceWire_4_bits_decodeResult_vwmacc;
  wire         validSource_4_bits_decodeResult_readOnly = laneRequestSourceWire_4_bits_decodeResult_readOnly;
  wire         validSource_4_bits_decodeResult_maskSource = laneRequestSourceWire_4_bits_decodeResult_maskSource;
  wire         validSource_4_bits_decodeResult_maskDestination = laneRequestSourceWire_4_bits_decodeResult_maskDestination;
  wire         validSource_4_bits_decodeResult_maskLogic = laneRequestSourceWire_4_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_4_bits_decodeResult_uop = laneRequestSourceWire_4_bits_decodeResult_uop;
  wire         validSource_4_bits_decodeResult_iota = laneRequestSourceWire_4_bits_decodeResult_iota;
  wire         validSource_4_bits_decodeResult_mv = laneRequestSourceWire_4_bits_decodeResult_mv;
  wire         validSource_4_bits_decodeResult_extend = laneRequestSourceWire_4_bits_decodeResult_extend;
  wire         validSource_4_bits_decodeResult_unOrderWrite = laneRequestSourceWire_4_bits_decodeResult_unOrderWrite;
  wire         validSource_4_bits_decodeResult_compress = laneRequestSourceWire_4_bits_decodeResult_compress;
  wire         validSource_4_bits_decodeResult_gather16 = laneRequestSourceWire_4_bits_decodeResult_gather16;
  wire         validSource_4_bits_decodeResult_gather = laneRequestSourceWire_4_bits_decodeResult_gather;
  wire         validSource_4_bits_decodeResult_slid = laneRequestSourceWire_4_bits_decodeResult_slid;
  wire         validSource_4_bits_decodeResult_targetRd = laneRequestSourceWire_4_bits_decodeResult_targetRd;
  wire         validSource_4_bits_decodeResult_widenReduce = laneRequestSourceWire_4_bits_decodeResult_widenReduce;
  wire         validSource_4_bits_decodeResult_red = laneRequestSourceWire_4_bits_decodeResult_red;
  wire         validSource_4_bits_decodeResult_nr = laneRequestSourceWire_4_bits_decodeResult_nr;
  wire         validSource_4_bits_decodeResult_itype = laneRequestSourceWire_4_bits_decodeResult_itype;
  wire         validSource_4_bits_decodeResult_unsigned1 = laneRequestSourceWire_4_bits_decodeResult_unsigned1;
  wire         validSource_4_bits_decodeResult_unsigned0 = laneRequestSourceWire_4_bits_decodeResult_unsigned0;
  wire         validSource_4_bits_decodeResult_other = laneRequestSourceWire_4_bits_decodeResult_other;
  wire         validSource_4_bits_decodeResult_multiCycle = laneRequestSourceWire_4_bits_decodeResult_multiCycle;
  wire         validSource_4_bits_decodeResult_divider = laneRequestSourceWire_4_bits_decodeResult_divider;
  wire         validSource_4_bits_decodeResult_multiplier = laneRequestSourceWire_4_bits_decodeResult_multiplier;
  wire         validSource_4_bits_decodeResult_shift = laneRequestSourceWire_4_bits_decodeResult_shift;
  wire         validSource_4_bits_decodeResult_adder = laneRequestSourceWire_4_bits_decodeResult_adder;
  wire         validSource_4_bits_decodeResult_logic = laneRequestSourceWire_4_bits_decodeResult_logic;
  wire         validSource_4_bits_loadStore = laneRequestSourceWire_4_bits_loadStore;
  wire         validSource_4_bits_issueInst = laneRequestSourceWire_4_bits_issueInst;
  wire         validSource_4_bits_store = laneRequestSourceWire_4_bits_store;
  wire         validSource_4_bits_special = laneRequestSourceWire_4_bits_special;
  wire         validSource_4_bits_lsWholeReg = laneRequestSourceWire_4_bits_lsWholeReg;
  wire [4:0]   validSource_4_bits_vs1 = laneRequestSourceWire_4_bits_vs1;
  wire [4:0]   validSource_4_bits_vs2 = laneRequestSourceWire_4_bits_vs2;
  wire [4:0]   validSource_4_bits_vd = laneRequestSourceWire_4_bits_vd;
  wire [1:0]   validSource_4_bits_loadStoreEEW = laneRequestSourceWire_4_bits_loadStoreEEW;
  wire         validSource_4_bits_mask = laneRequestSourceWire_4_bits_mask;
  wire [2:0]   validSource_4_bits_segment = laneRequestSourceWire_4_bits_segment;
  wire [31:0]  validSource_4_bits_readFromScalar = laneRequestSourceWire_4_bits_readFromScalar;
  wire [11:0]  validSource_4_bits_csrInterface_vl = laneRequestSourceWire_4_bits_csrInterface_vl;
  wire [11:0]  validSource_4_bits_csrInterface_vStart = laneRequestSourceWire_4_bits_csrInterface_vStart;
  wire [2:0]   validSource_4_bits_csrInterface_vlmul = laneRequestSourceWire_4_bits_csrInterface_vlmul;
  wire [1:0]   validSource_4_bits_csrInterface_vSew = laneRequestSourceWire_4_bits_csrInterface_vSew;
  wire [1:0]   validSource_4_bits_csrInterface_vxrm = laneRequestSourceWire_4_bits_csrInterface_vxrm;
  wire         validSource_4_bits_csrInterface_vta = laneRequestSourceWire_4_bits_csrInterface_vta;
  wire         validSource_4_bits_csrInterface_vma = laneRequestSourceWire_4_bits_csrInterface_vma;
  wire         tokenCheck_5;
  wire [2:0]   validSource_5_bits_instructionIndex = laneRequestSourceWire_5_bits_instructionIndex;
  wire         validSource_5_bits_decodeResult_orderReduce = laneRequestSourceWire_5_bits_decodeResult_orderReduce;
  wire         validSource_5_bits_decodeResult_floatMul = laneRequestSourceWire_5_bits_decodeResult_floatMul;
  wire [1:0]   validSource_5_bits_decodeResult_fpExecutionType = laneRequestSourceWire_5_bits_decodeResult_fpExecutionType;
  wire         validSource_5_bits_decodeResult_float = laneRequestSourceWire_5_bits_decodeResult_float;
  wire         validSource_5_bits_decodeResult_specialSlot = laneRequestSourceWire_5_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_5_bits_decodeResult_topUop = laneRequestSourceWire_5_bits_decodeResult_topUop;
  wire         validSource_5_bits_decodeResult_popCount = laneRequestSourceWire_5_bits_decodeResult_popCount;
  wire         validSource_5_bits_decodeResult_ffo = laneRequestSourceWire_5_bits_decodeResult_ffo;
  wire         validSource_5_bits_decodeResult_average = laneRequestSourceWire_5_bits_decodeResult_average;
  wire         validSource_5_bits_decodeResult_reverse = laneRequestSourceWire_5_bits_decodeResult_reverse;
  wire         validSource_5_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_5_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_5_bits_decodeResult_scheduler = laneRequestSourceWire_5_bits_decodeResult_scheduler;
  wire         validSource_5_bits_decodeResult_sReadVD = laneRequestSourceWire_5_bits_decodeResult_sReadVD;
  wire         validSource_5_bits_decodeResult_vtype = laneRequestSourceWire_5_bits_decodeResult_vtype;
  wire         validSource_5_bits_decodeResult_sWrite = laneRequestSourceWire_5_bits_decodeResult_sWrite;
  wire         validSource_5_bits_decodeResult_crossRead = laneRequestSourceWire_5_bits_decodeResult_crossRead;
  wire         validSource_5_bits_decodeResult_crossWrite = laneRequestSourceWire_5_bits_decodeResult_crossWrite;
  wire         validSource_5_bits_decodeResult_maskUnit = laneRequestSourceWire_5_bits_decodeResult_maskUnit;
  wire         validSource_5_bits_decodeResult_special = laneRequestSourceWire_5_bits_decodeResult_special;
  wire         validSource_5_bits_decodeResult_saturate = laneRequestSourceWire_5_bits_decodeResult_saturate;
  wire         validSource_5_bits_decodeResult_vwmacc = laneRequestSourceWire_5_bits_decodeResult_vwmacc;
  wire         validSource_5_bits_decodeResult_readOnly = laneRequestSourceWire_5_bits_decodeResult_readOnly;
  wire         validSource_5_bits_decodeResult_maskSource = laneRequestSourceWire_5_bits_decodeResult_maskSource;
  wire         validSource_5_bits_decodeResult_maskDestination = laneRequestSourceWire_5_bits_decodeResult_maskDestination;
  wire         validSource_5_bits_decodeResult_maskLogic = laneRequestSourceWire_5_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_5_bits_decodeResult_uop = laneRequestSourceWire_5_bits_decodeResult_uop;
  wire         validSource_5_bits_decodeResult_iota = laneRequestSourceWire_5_bits_decodeResult_iota;
  wire         validSource_5_bits_decodeResult_mv = laneRequestSourceWire_5_bits_decodeResult_mv;
  wire         validSource_5_bits_decodeResult_extend = laneRequestSourceWire_5_bits_decodeResult_extend;
  wire         validSource_5_bits_decodeResult_unOrderWrite = laneRequestSourceWire_5_bits_decodeResult_unOrderWrite;
  wire         validSource_5_bits_decodeResult_compress = laneRequestSourceWire_5_bits_decodeResult_compress;
  wire         validSource_5_bits_decodeResult_gather16 = laneRequestSourceWire_5_bits_decodeResult_gather16;
  wire         validSource_5_bits_decodeResult_gather = laneRequestSourceWire_5_bits_decodeResult_gather;
  wire         validSource_5_bits_decodeResult_slid = laneRequestSourceWire_5_bits_decodeResult_slid;
  wire         validSource_5_bits_decodeResult_targetRd = laneRequestSourceWire_5_bits_decodeResult_targetRd;
  wire         validSource_5_bits_decodeResult_widenReduce = laneRequestSourceWire_5_bits_decodeResult_widenReduce;
  wire         validSource_5_bits_decodeResult_red = laneRequestSourceWire_5_bits_decodeResult_red;
  wire         validSource_5_bits_decodeResult_nr = laneRequestSourceWire_5_bits_decodeResult_nr;
  wire         validSource_5_bits_decodeResult_itype = laneRequestSourceWire_5_bits_decodeResult_itype;
  wire         validSource_5_bits_decodeResult_unsigned1 = laneRequestSourceWire_5_bits_decodeResult_unsigned1;
  wire         validSource_5_bits_decodeResult_unsigned0 = laneRequestSourceWire_5_bits_decodeResult_unsigned0;
  wire         validSource_5_bits_decodeResult_other = laneRequestSourceWire_5_bits_decodeResult_other;
  wire         validSource_5_bits_decodeResult_multiCycle = laneRequestSourceWire_5_bits_decodeResult_multiCycle;
  wire         validSource_5_bits_decodeResult_divider = laneRequestSourceWire_5_bits_decodeResult_divider;
  wire         validSource_5_bits_decodeResult_multiplier = laneRequestSourceWire_5_bits_decodeResult_multiplier;
  wire         validSource_5_bits_decodeResult_shift = laneRequestSourceWire_5_bits_decodeResult_shift;
  wire         validSource_5_bits_decodeResult_adder = laneRequestSourceWire_5_bits_decodeResult_adder;
  wire         validSource_5_bits_decodeResult_logic = laneRequestSourceWire_5_bits_decodeResult_logic;
  wire         validSource_5_bits_loadStore = laneRequestSourceWire_5_bits_loadStore;
  wire         validSource_5_bits_issueInst = laneRequestSourceWire_5_bits_issueInst;
  wire         validSource_5_bits_store = laneRequestSourceWire_5_bits_store;
  wire         validSource_5_bits_special = laneRequestSourceWire_5_bits_special;
  wire         validSource_5_bits_lsWholeReg = laneRequestSourceWire_5_bits_lsWholeReg;
  wire [4:0]   validSource_5_bits_vs1 = laneRequestSourceWire_5_bits_vs1;
  wire [4:0]   validSource_5_bits_vs2 = laneRequestSourceWire_5_bits_vs2;
  wire [4:0]   validSource_5_bits_vd = laneRequestSourceWire_5_bits_vd;
  wire [1:0]   validSource_5_bits_loadStoreEEW = laneRequestSourceWire_5_bits_loadStoreEEW;
  wire         validSource_5_bits_mask = laneRequestSourceWire_5_bits_mask;
  wire [2:0]   validSource_5_bits_segment = laneRequestSourceWire_5_bits_segment;
  wire [31:0]  validSource_5_bits_readFromScalar = laneRequestSourceWire_5_bits_readFromScalar;
  wire [11:0]  validSource_5_bits_csrInterface_vl = laneRequestSourceWire_5_bits_csrInterface_vl;
  wire [11:0]  validSource_5_bits_csrInterface_vStart = laneRequestSourceWire_5_bits_csrInterface_vStart;
  wire [2:0]   validSource_5_bits_csrInterface_vlmul = laneRequestSourceWire_5_bits_csrInterface_vlmul;
  wire [1:0]   validSource_5_bits_csrInterface_vSew = laneRequestSourceWire_5_bits_csrInterface_vSew;
  wire [1:0]   validSource_5_bits_csrInterface_vxrm = laneRequestSourceWire_5_bits_csrInterface_vxrm;
  wire         validSource_5_bits_csrInterface_vta = laneRequestSourceWire_5_bits_csrInterface_vta;
  wire         validSource_5_bits_csrInterface_vma = laneRequestSourceWire_5_bits_csrInterface_vma;
  wire         tokenCheck_6;
  wire [2:0]   validSource_6_bits_instructionIndex = laneRequestSourceWire_6_bits_instructionIndex;
  wire         validSource_6_bits_decodeResult_orderReduce = laneRequestSourceWire_6_bits_decodeResult_orderReduce;
  wire         validSource_6_bits_decodeResult_floatMul = laneRequestSourceWire_6_bits_decodeResult_floatMul;
  wire [1:0]   validSource_6_bits_decodeResult_fpExecutionType = laneRequestSourceWire_6_bits_decodeResult_fpExecutionType;
  wire         validSource_6_bits_decodeResult_float = laneRequestSourceWire_6_bits_decodeResult_float;
  wire         validSource_6_bits_decodeResult_specialSlot = laneRequestSourceWire_6_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_6_bits_decodeResult_topUop = laneRequestSourceWire_6_bits_decodeResult_topUop;
  wire         validSource_6_bits_decodeResult_popCount = laneRequestSourceWire_6_bits_decodeResult_popCount;
  wire         validSource_6_bits_decodeResult_ffo = laneRequestSourceWire_6_bits_decodeResult_ffo;
  wire         validSource_6_bits_decodeResult_average = laneRequestSourceWire_6_bits_decodeResult_average;
  wire         validSource_6_bits_decodeResult_reverse = laneRequestSourceWire_6_bits_decodeResult_reverse;
  wire         validSource_6_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_6_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_6_bits_decodeResult_scheduler = laneRequestSourceWire_6_bits_decodeResult_scheduler;
  wire         validSource_6_bits_decodeResult_sReadVD = laneRequestSourceWire_6_bits_decodeResult_sReadVD;
  wire         validSource_6_bits_decodeResult_vtype = laneRequestSourceWire_6_bits_decodeResult_vtype;
  wire         validSource_6_bits_decodeResult_sWrite = laneRequestSourceWire_6_bits_decodeResult_sWrite;
  wire         validSource_6_bits_decodeResult_crossRead = laneRequestSourceWire_6_bits_decodeResult_crossRead;
  wire         validSource_6_bits_decodeResult_crossWrite = laneRequestSourceWire_6_bits_decodeResult_crossWrite;
  wire         validSource_6_bits_decodeResult_maskUnit = laneRequestSourceWire_6_bits_decodeResult_maskUnit;
  wire         validSource_6_bits_decodeResult_special = laneRequestSourceWire_6_bits_decodeResult_special;
  wire         validSource_6_bits_decodeResult_saturate = laneRequestSourceWire_6_bits_decodeResult_saturate;
  wire         validSource_6_bits_decodeResult_vwmacc = laneRequestSourceWire_6_bits_decodeResult_vwmacc;
  wire         validSource_6_bits_decodeResult_readOnly = laneRequestSourceWire_6_bits_decodeResult_readOnly;
  wire         validSource_6_bits_decodeResult_maskSource = laneRequestSourceWire_6_bits_decodeResult_maskSource;
  wire         validSource_6_bits_decodeResult_maskDestination = laneRequestSourceWire_6_bits_decodeResult_maskDestination;
  wire         validSource_6_bits_decodeResult_maskLogic = laneRequestSourceWire_6_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_6_bits_decodeResult_uop = laneRequestSourceWire_6_bits_decodeResult_uop;
  wire         validSource_6_bits_decodeResult_iota = laneRequestSourceWire_6_bits_decodeResult_iota;
  wire         validSource_6_bits_decodeResult_mv = laneRequestSourceWire_6_bits_decodeResult_mv;
  wire         validSource_6_bits_decodeResult_extend = laneRequestSourceWire_6_bits_decodeResult_extend;
  wire         validSource_6_bits_decodeResult_unOrderWrite = laneRequestSourceWire_6_bits_decodeResult_unOrderWrite;
  wire         validSource_6_bits_decodeResult_compress = laneRequestSourceWire_6_bits_decodeResult_compress;
  wire         validSource_6_bits_decodeResult_gather16 = laneRequestSourceWire_6_bits_decodeResult_gather16;
  wire         validSource_6_bits_decodeResult_gather = laneRequestSourceWire_6_bits_decodeResult_gather;
  wire         validSource_6_bits_decodeResult_slid = laneRequestSourceWire_6_bits_decodeResult_slid;
  wire         validSource_6_bits_decodeResult_targetRd = laneRequestSourceWire_6_bits_decodeResult_targetRd;
  wire         validSource_6_bits_decodeResult_widenReduce = laneRequestSourceWire_6_bits_decodeResult_widenReduce;
  wire         validSource_6_bits_decodeResult_red = laneRequestSourceWire_6_bits_decodeResult_red;
  wire         validSource_6_bits_decodeResult_nr = laneRequestSourceWire_6_bits_decodeResult_nr;
  wire         validSource_6_bits_decodeResult_itype = laneRequestSourceWire_6_bits_decodeResult_itype;
  wire         validSource_6_bits_decodeResult_unsigned1 = laneRequestSourceWire_6_bits_decodeResult_unsigned1;
  wire         validSource_6_bits_decodeResult_unsigned0 = laneRequestSourceWire_6_bits_decodeResult_unsigned0;
  wire         validSource_6_bits_decodeResult_other = laneRequestSourceWire_6_bits_decodeResult_other;
  wire         validSource_6_bits_decodeResult_multiCycle = laneRequestSourceWire_6_bits_decodeResult_multiCycle;
  wire         validSource_6_bits_decodeResult_divider = laneRequestSourceWire_6_bits_decodeResult_divider;
  wire         validSource_6_bits_decodeResult_multiplier = laneRequestSourceWire_6_bits_decodeResult_multiplier;
  wire         validSource_6_bits_decodeResult_shift = laneRequestSourceWire_6_bits_decodeResult_shift;
  wire         validSource_6_bits_decodeResult_adder = laneRequestSourceWire_6_bits_decodeResult_adder;
  wire         validSource_6_bits_decodeResult_logic = laneRequestSourceWire_6_bits_decodeResult_logic;
  wire         validSource_6_bits_loadStore = laneRequestSourceWire_6_bits_loadStore;
  wire         validSource_6_bits_issueInst = laneRequestSourceWire_6_bits_issueInst;
  wire         validSource_6_bits_store = laneRequestSourceWire_6_bits_store;
  wire         validSource_6_bits_special = laneRequestSourceWire_6_bits_special;
  wire         validSource_6_bits_lsWholeReg = laneRequestSourceWire_6_bits_lsWholeReg;
  wire [4:0]   validSource_6_bits_vs1 = laneRequestSourceWire_6_bits_vs1;
  wire [4:0]   validSource_6_bits_vs2 = laneRequestSourceWire_6_bits_vs2;
  wire [4:0]   validSource_6_bits_vd = laneRequestSourceWire_6_bits_vd;
  wire [1:0]   validSource_6_bits_loadStoreEEW = laneRequestSourceWire_6_bits_loadStoreEEW;
  wire         validSource_6_bits_mask = laneRequestSourceWire_6_bits_mask;
  wire [2:0]   validSource_6_bits_segment = laneRequestSourceWire_6_bits_segment;
  wire [31:0]  validSource_6_bits_readFromScalar = laneRequestSourceWire_6_bits_readFromScalar;
  wire [11:0]  validSource_6_bits_csrInterface_vl = laneRequestSourceWire_6_bits_csrInterface_vl;
  wire [11:0]  validSource_6_bits_csrInterface_vStart = laneRequestSourceWire_6_bits_csrInterface_vStart;
  wire [2:0]   validSource_6_bits_csrInterface_vlmul = laneRequestSourceWire_6_bits_csrInterface_vlmul;
  wire [1:0]   validSource_6_bits_csrInterface_vSew = laneRequestSourceWire_6_bits_csrInterface_vSew;
  wire [1:0]   validSource_6_bits_csrInterface_vxrm = laneRequestSourceWire_6_bits_csrInterface_vxrm;
  wire         validSource_6_bits_csrInterface_vta = laneRequestSourceWire_6_bits_csrInterface_vta;
  wire         validSource_6_bits_csrInterface_vma = laneRequestSourceWire_6_bits_csrInterface_vma;
  wire         tokenCheck_7;
  wire [2:0]   validSource_7_bits_instructionIndex = laneRequestSourceWire_7_bits_instructionIndex;
  wire         validSource_7_bits_decodeResult_orderReduce = laneRequestSourceWire_7_bits_decodeResult_orderReduce;
  wire         validSource_7_bits_decodeResult_floatMul = laneRequestSourceWire_7_bits_decodeResult_floatMul;
  wire [1:0]   validSource_7_bits_decodeResult_fpExecutionType = laneRequestSourceWire_7_bits_decodeResult_fpExecutionType;
  wire         validSource_7_bits_decodeResult_float = laneRequestSourceWire_7_bits_decodeResult_float;
  wire         validSource_7_bits_decodeResult_specialSlot = laneRequestSourceWire_7_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_7_bits_decodeResult_topUop = laneRequestSourceWire_7_bits_decodeResult_topUop;
  wire         validSource_7_bits_decodeResult_popCount = laneRequestSourceWire_7_bits_decodeResult_popCount;
  wire         validSource_7_bits_decodeResult_ffo = laneRequestSourceWire_7_bits_decodeResult_ffo;
  wire         validSource_7_bits_decodeResult_average = laneRequestSourceWire_7_bits_decodeResult_average;
  wire         validSource_7_bits_decodeResult_reverse = laneRequestSourceWire_7_bits_decodeResult_reverse;
  wire         validSource_7_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_7_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_7_bits_decodeResult_scheduler = laneRequestSourceWire_7_bits_decodeResult_scheduler;
  wire         validSource_7_bits_decodeResult_sReadVD = laneRequestSourceWire_7_bits_decodeResult_sReadVD;
  wire         validSource_7_bits_decodeResult_vtype = laneRequestSourceWire_7_bits_decodeResult_vtype;
  wire         validSource_7_bits_decodeResult_sWrite = laneRequestSourceWire_7_bits_decodeResult_sWrite;
  wire         validSource_7_bits_decodeResult_crossRead = laneRequestSourceWire_7_bits_decodeResult_crossRead;
  wire         validSource_7_bits_decodeResult_crossWrite = laneRequestSourceWire_7_bits_decodeResult_crossWrite;
  wire         validSource_7_bits_decodeResult_maskUnit = laneRequestSourceWire_7_bits_decodeResult_maskUnit;
  wire         validSource_7_bits_decodeResult_special = laneRequestSourceWire_7_bits_decodeResult_special;
  wire         validSource_7_bits_decodeResult_saturate = laneRequestSourceWire_7_bits_decodeResult_saturate;
  wire         validSource_7_bits_decodeResult_vwmacc = laneRequestSourceWire_7_bits_decodeResult_vwmacc;
  wire         validSource_7_bits_decodeResult_readOnly = laneRequestSourceWire_7_bits_decodeResult_readOnly;
  wire         validSource_7_bits_decodeResult_maskSource = laneRequestSourceWire_7_bits_decodeResult_maskSource;
  wire         validSource_7_bits_decodeResult_maskDestination = laneRequestSourceWire_7_bits_decodeResult_maskDestination;
  wire         validSource_7_bits_decodeResult_maskLogic = laneRequestSourceWire_7_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_7_bits_decodeResult_uop = laneRequestSourceWire_7_bits_decodeResult_uop;
  wire         validSource_7_bits_decodeResult_iota = laneRequestSourceWire_7_bits_decodeResult_iota;
  wire         validSource_7_bits_decodeResult_mv = laneRequestSourceWire_7_bits_decodeResult_mv;
  wire         validSource_7_bits_decodeResult_extend = laneRequestSourceWire_7_bits_decodeResult_extend;
  wire         validSource_7_bits_decodeResult_unOrderWrite = laneRequestSourceWire_7_bits_decodeResult_unOrderWrite;
  wire         validSource_7_bits_decodeResult_compress = laneRequestSourceWire_7_bits_decodeResult_compress;
  wire         validSource_7_bits_decodeResult_gather16 = laneRequestSourceWire_7_bits_decodeResult_gather16;
  wire         validSource_7_bits_decodeResult_gather = laneRequestSourceWire_7_bits_decodeResult_gather;
  wire         validSource_7_bits_decodeResult_slid = laneRequestSourceWire_7_bits_decodeResult_slid;
  wire         validSource_7_bits_decodeResult_targetRd = laneRequestSourceWire_7_bits_decodeResult_targetRd;
  wire         validSource_7_bits_decodeResult_widenReduce = laneRequestSourceWire_7_bits_decodeResult_widenReduce;
  wire         validSource_7_bits_decodeResult_red = laneRequestSourceWire_7_bits_decodeResult_red;
  wire         validSource_7_bits_decodeResult_nr = laneRequestSourceWire_7_bits_decodeResult_nr;
  wire         validSource_7_bits_decodeResult_itype = laneRequestSourceWire_7_bits_decodeResult_itype;
  wire         validSource_7_bits_decodeResult_unsigned1 = laneRequestSourceWire_7_bits_decodeResult_unsigned1;
  wire         validSource_7_bits_decodeResult_unsigned0 = laneRequestSourceWire_7_bits_decodeResult_unsigned0;
  wire         validSource_7_bits_decodeResult_other = laneRequestSourceWire_7_bits_decodeResult_other;
  wire         validSource_7_bits_decodeResult_multiCycle = laneRequestSourceWire_7_bits_decodeResult_multiCycle;
  wire         validSource_7_bits_decodeResult_divider = laneRequestSourceWire_7_bits_decodeResult_divider;
  wire         validSource_7_bits_decodeResult_multiplier = laneRequestSourceWire_7_bits_decodeResult_multiplier;
  wire         validSource_7_bits_decodeResult_shift = laneRequestSourceWire_7_bits_decodeResult_shift;
  wire         validSource_7_bits_decodeResult_adder = laneRequestSourceWire_7_bits_decodeResult_adder;
  wire         validSource_7_bits_decodeResult_logic = laneRequestSourceWire_7_bits_decodeResult_logic;
  wire         validSource_7_bits_loadStore = laneRequestSourceWire_7_bits_loadStore;
  wire         validSource_7_bits_issueInst = laneRequestSourceWire_7_bits_issueInst;
  wire         validSource_7_bits_store = laneRequestSourceWire_7_bits_store;
  wire         validSource_7_bits_special = laneRequestSourceWire_7_bits_special;
  wire         validSource_7_bits_lsWholeReg = laneRequestSourceWire_7_bits_lsWholeReg;
  wire [4:0]   validSource_7_bits_vs1 = laneRequestSourceWire_7_bits_vs1;
  wire [4:0]   validSource_7_bits_vs2 = laneRequestSourceWire_7_bits_vs2;
  wire [4:0]   validSource_7_bits_vd = laneRequestSourceWire_7_bits_vd;
  wire [1:0]   validSource_7_bits_loadStoreEEW = laneRequestSourceWire_7_bits_loadStoreEEW;
  wire         validSource_7_bits_mask = laneRequestSourceWire_7_bits_mask;
  wire [2:0]   validSource_7_bits_segment = laneRequestSourceWire_7_bits_segment;
  wire [31:0]  validSource_7_bits_readFromScalar = laneRequestSourceWire_7_bits_readFromScalar;
  wire [11:0]  validSource_7_bits_csrInterface_vl = laneRequestSourceWire_7_bits_csrInterface_vl;
  wire [11:0]  validSource_7_bits_csrInterface_vStart = laneRequestSourceWire_7_bits_csrInterface_vStart;
  wire [2:0]   validSource_7_bits_csrInterface_vlmul = laneRequestSourceWire_7_bits_csrInterface_vlmul;
  wire [1:0]   validSource_7_bits_csrInterface_vSew = laneRequestSourceWire_7_bits_csrInterface_vSew;
  wire [1:0]   validSource_7_bits_csrInterface_vxrm = laneRequestSourceWire_7_bits_csrInterface_vxrm;
  wire         validSource_7_bits_csrInterface_vta = laneRequestSourceWire_7_bits_csrInterface_vta;
  wire         validSource_7_bits_csrInterface_vma = laneRequestSourceWire_7_bits_csrInterface_vma;
  wire         tokenCheck_8;
  wire [2:0]   validSource_8_bits_instructionIndex = laneRequestSourceWire_8_bits_instructionIndex;
  wire         validSource_8_bits_decodeResult_orderReduce = laneRequestSourceWire_8_bits_decodeResult_orderReduce;
  wire         validSource_8_bits_decodeResult_floatMul = laneRequestSourceWire_8_bits_decodeResult_floatMul;
  wire [1:0]   validSource_8_bits_decodeResult_fpExecutionType = laneRequestSourceWire_8_bits_decodeResult_fpExecutionType;
  wire         validSource_8_bits_decodeResult_float = laneRequestSourceWire_8_bits_decodeResult_float;
  wire         validSource_8_bits_decodeResult_specialSlot = laneRequestSourceWire_8_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_8_bits_decodeResult_topUop = laneRequestSourceWire_8_bits_decodeResult_topUop;
  wire         validSource_8_bits_decodeResult_popCount = laneRequestSourceWire_8_bits_decodeResult_popCount;
  wire         validSource_8_bits_decodeResult_ffo = laneRequestSourceWire_8_bits_decodeResult_ffo;
  wire         validSource_8_bits_decodeResult_average = laneRequestSourceWire_8_bits_decodeResult_average;
  wire         validSource_8_bits_decodeResult_reverse = laneRequestSourceWire_8_bits_decodeResult_reverse;
  wire         validSource_8_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_8_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_8_bits_decodeResult_scheduler = laneRequestSourceWire_8_bits_decodeResult_scheduler;
  wire         validSource_8_bits_decodeResult_sReadVD = laneRequestSourceWire_8_bits_decodeResult_sReadVD;
  wire         validSource_8_bits_decodeResult_vtype = laneRequestSourceWire_8_bits_decodeResult_vtype;
  wire         validSource_8_bits_decodeResult_sWrite = laneRequestSourceWire_8_bits_decodeResult_sWrite;
  wire         validSource_8_bits_decodeResult_crossRead = laneRequestSourceWire_8_bits_decodeResult_crossRead;
  wire         validSource_8_bits_decodeResult_crossWrite = laneRequestSourceWire_8_bits_decodeResult_crossWrite;
  wire         validSource_8_bits_decodeResult_maskUnit = laneRequestSourceWire_8_bits_decodeResult_maskUnit;
  wire         validSource_8_bits_decodeResult_special = laneRequestSourceWire_8_bits_decodeResult_special;
  wire         validSource_8_bits_decodeResult_saturate = laneRequestSourceWire_8_bits_decodeResult_saturate;
  wire         validSource_8_bits_decodeResult_vwmacc = laneRequestSourceWire_8_bits_decodeResult_vwmacc;
  wire         validSource_8_bits_decodeResult_readOnly = laneRequestSourceWire_8_bits_decodeResult_readOnly;
  wire         validSource_8_bits_decodeResult_maskSource = laneRequestSourceWire_8_bits_decodeResult_maskSource;
  wire         validSource_8_bits_decodeResult_maskDestination = laneRequestSourceWire_8_bits_decodeResult_maskDestination;
  wire         validSource_8_bits_decodeResult_maskLogic = laneRequestSourceWire_8_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_8_bits_decodeResult_uop = laneRequestSourceWire_8_bits_decodeResult_uop;
  wire         validSource_8_bits_decodeResult_iota = laneRequestSourceWire_8_bits_decodeResult_iota;
  wire         validSource_8_bits_decodeResult_mv = laneRequestSourceWire_8_bits_decodeResult_mv;
  wire         validSource_8_bits_decodeResult_extend = laneRequestSourceWire_8_bits_decodeResult_extend;
  wire         validSource_8_bits_decodeResult_unOrderWrite = laneRequestSourceWire_8_bits_decodeResult_unOrderWrite;
  wire         validSource_8_bits_decodeResult_compress = laneRequestSourceWire_8_bits_decodeResult_compress;
  wire         validSource_8_bits_decodeResult_gather16 = laneRequestSourceWire_8_bits_decodeResult_gather16;
  wire         validSource_8_bits_decodeResult_gather = laneRequestSourceWire_8_bits_decodeResult_gather;
  wire         validSource_8_bits_decodeResult_slid = laneRequestSourceWire_8_bits_decodeResult_slid;
  wire         validSource_8_bits_decodeResult_targetRd = laneRequestSourceWire_8_bits_decodeResult_targetRd;
  wire         validSource_8_bits_decodeResult_widenReduce = laneRequestSourceWire_8_bits_decodeResult_widenReduce;
  wire         validSource_8_bits_decodeResult_red = laneRequestSourceWire_8_bits_decodeResult_red;
  wire         validSource_8_bits_decodeResult_nr = laneRequestSourceWire_8_bits_decodeResult_nr;
  wire         validSource_8_bits_decodeResult_itype = laneRequestSourceWire_8_bits_decodeResult_itype;
  wire         validSource_8_bits_decodeResult_unsigned1 = laneRequestSourceWire_8_bits_decodeResult_unsigned1;
  wire         validSource_8_bits_decodeResult_unsigned0 = laneRequestSourceWire_8_bits_decodeResult_unsigned0;
  wire         validSource_8_bits_decodeResult_other = laneRequestSourceWire_8_bits_decodeResult_other;
  wire         validSource_8_bits_decodeResult_multiCycle = laneRequestSourceWire_8_bits_decodeResult_multiCycle;
  wire         validSource_8_bits_decodeResult_divider = laneRequestSourceWire_8_bits_decodeResult_divider;
  wire         validSource_8_bits_decodeResult_multiplier = laneRequestSourceWire_8_bits_decodeResult_multiplier;
  wire         validSource_8_bits_decodeResult_shift = laneRequestSourceWire_8_bits_decodeResult_shift;
  wire         validSource_8_bits_decodeResult_adder = laneRequestSourceWire_8_bits_decodeResult_adder;
  wire         validSource_8_bits_decodeResult_logic = laneRequestSourceWire_8_bits_decodeResult_logic;
  wire         validSource_8_bits_loadStore = laneRequestSourceWire_8_bits_loadStore;
  wire         validSource_8_bits_issueInst = laneRequestSourceWire_8_bits_issueInst;
  wire         validSource_8_bits_store = laneRequestSourceWire_8_bits_store;
  wire         validSource_8_bits_special = laneRequestSourceWire_8_bits_special;
  wire         validSource_8_bits_lsWholeReg = laneRequestSourceWire_8_bits_lsWholeReg;
  wire [4:0]   validSource_8_bits_vs1 = laneRequestSourceWire_8_bits_vs1;
  wire [4:0]   validSource_8_bits_vs2 = laneRequestSourceWire_8_bits_vs2;
  wire [4:0]   validSource_8_bits_vd = laneRequestSourceWire_8_bits_vd;
  wire [1:0]   validSource_8_bits_loadStoreEEW = laneRequestSourceWire_8_bits_loadStoreEEW;
  wire         validSource_8_bits_mask = laneRequestSourceWire_8_bits_mask;
  wire [2:0]   validSource_8_bits_segment = laneRequestSourceWire_8_bits_segment;
  wire [31:0]  validSource_8_bits_readFromScalar = laneRequestSourceWire_8_bits_readFromScalar;
  wire [11:0]  validSource_8_bits_csrInterface_vl = laneRequestSourceWire_8_bits_csrInterface_vl;
  wire [11:0]  validSource_8_bits_csrInterface_vStart = laneRequestSourceWire_8_bits_csrInterface_vStart;
  wire [2:0]   validSource_8_bits_csrInterface_vlmul = laneRequestSourceWire_8_bits_csrInterface_vlmul;
  wire [1:0]   validSource_8_bits_csrInterface_vSew = laneRequestSourceWire_8_bits_csrInterface_vSew;
  wire [1:0]   validSource_8_bits_csrInterface_vxrm = laneRequestSourceWire_8_bits_csrInterface_vxrm;
  wire         validSource_8_bits_csrInterface_vta = laneRequestSourceWire_8_bits_csrInterface_vta;
  wire         validSource_8_bits_csrInterface_vma = laneRequestSourceWire_8_bits_csrInterface_vma;
  wire         tokenCheck_9;
  wire [2:0]   validSource_9_bits_instructionIndex = laneRequestSourceWire_9_bits_instructionIndex;
  wire         validSource_9_bits_decodeResult_orderReduce = laneRequestSourceWire_9_bits_decodeResult_orderReduce;
  wire         validSource_9_bits_decodeResult_floatMul = laneRequestSourceWire_9_bits_decodeResult_floatMul;
  wire [1:0]   validSource_9_bits_decodeResult_fpExecutionType = laneRequestSourceWire_9_bits_decodeResult_fpExecutionType;
  wire         validSource_9_bits_decodeResult_float = laneRequestSourceWire_9_bits_decodeResult_float;
  wire         validSource_9_bits_decodeResult_specialSlot = laneRequestSourceWire_9_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_9_bits_decodeResult_topUop = laneRequestSourceWire_9_bits_decodeResult_topUop;
  wire         validSource_9_bits_decodeResult_popCount = laneRequestSourceWire_9_bits_decodeResult_popCount;
  wire         validSource_9_bits_decodeResult_ffo = laneRequestSourceWire_9_bits_decodeResult_ffo;
  wire         validSource_9_bits_decodeResult_average = laneRequestSourceWire_9_bits_decodeResult_average;
  wire         validSource_9_bits_decodeResult_reverse = laneRequestSourceWire_9_bits_decodeResult_reverse;
  wire         validSource_9_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_9_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_9_bits_decodeResult_scheduler = laneRequestSourceWire_9_bits_decodeResult_scheduler;
  wire         validSource_9_bits_decodeResult_sReadVD = laneRequestSourceWire_9_bits_decodeResult_sReadVD;
  wire         validSource_9_bits_decodeResult_vtype = laneRequestSourceWire_9_bits_decodeResult_vtype;
  wire         validSource_9_bits_decodeResult_sWrite = laneRequestSourceWire_9_bits_decodeResult_sWrite;
  wire         validSource_9_bits_decodeResult_crossRead = laneRequestSourceWire_9_bits_decodeResult_crossRead;
  wire         validSource_9_bits_decodeResult_crossWrite = laneRequestSourceWire_9_bits_decodeResult_crossWrite;
  wire         validSource_9_bits_decodeResult_maskUnit = laneRequestSourceWire_9_bits_decodeResult_maskUnit;
  wire         validSource_9_bits_decodeResult_special = laneRequestSourceWire_9_bits_decodeResult_special;
  wire         validSource_9_bits_decodeResult_saturate = laneRequestSourceWire_9_bits_decodeResult_saturate;
  wire         validSource_9_bits_decodeResult_vwmacc = laneRequestSourceWire_9_bits_decodeResult_vwmacc;
  wire         validSource_9_bits_decodeResult_readOnly = laneRequestSourceWire_9_bits_decodeResult_readOnly;
  wire         validSource_9_bits_decodeResult_maskSource = laneRequestSourceWire_9_bits_decodeResult_maskSource;
  wire         validSource_9_bits_decodeResult_maskDestination = laneRequestSourceWire_9_bits_decodeResult_maskDestination;
  wire         validSource_9_bits_decodeResult_maskLogic = laneRequestSourceWire_9_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_9_bits_decodeResult_uop = laneRequestSourceWire_9_bits_decodeResult_uop;
  wire         validSource_9_bits_decodeResult_iota = laneRequestSourceWire_9_bits_decodeResult_iota;
  wire         validSource_9_bits_decodeResult_mv = laneRequestSourceWire_9_bits_decodeResult_mv;
  wire         validSource_9_bits_decodeResult_extend = laneRequestSourceWire_9_bits_decodeResult_extend;
  wire         validSource_9_bits_decodeResult_unOrderWrite = laneRequestSourceWire_9_bits_decodeResult_unOrderWrite;
  wire         validSource_9_bits_decodeResult_compress = laneRequestSourceWire_9_bits_decodeResult_compress;
  wire         validSource_9_bits_decodeResult_gather16 = laneRequestSourceWire_9_bits_decodeResult_gather16;
  wire         validSource_9_bits_decodeResult_gather = laneRequestSourceWire_9_bits_decodeResult_gather;
  wire         validSource_9_bits_decodeResult_slid = laneRequestSourceWire_9_bits_decodeResult_slid;
  wire         validSource_9_bits_decodeResult_targetRd = laneRequestSourceWire_9_bits_decodeResult_targetRd;
  wire         validSource_9_bits_decodeResult_widenReduce = laneRequestSourceWire_9_bits_decodeResult_widenReduce;
  wire         validSource_9_bits_decodeResult_red = laneRequestSourceWire_9_bits_decodeResult_red;
  wire         validSource_9_bits_decodeResult_nr = laneRequestSourceWire_9_bits_decodeResult_nr;
  wire         validSource_9_bits_decodeResult_itype = laneRequestSourceWire_9_bits_decodeResult_itype;
  wire         validSource_9_bits_decodeResult_unsigned1 = laneRequestSourceWire_9_bits_decodeResult_unsigned1;
  wire         validSource_9_bits_decodeResult_unsigned0 = laneRequestSourceWire_9_bits_decodeResult_unsigned0;
  wire         validSource_9_bits_decodeResult_other = laneRequestSourceWire_9_bits_decodeResult_other;
  wire         validSource_9_bits_decodeResult_multiCycle = laneRequestSourceWire_9_bits_decodeResult_multiCycle;
  wire         validSource_9_bits_decodeResult_divider = laneRequestSourceWire_9_bits_decodeResult_divider;
  wire         validSource_9_bits_decodeResult_multiplier = laneRequestSourceWire_9_bits_decodeResult_multiplier;
  wire         validSource_9_bits_decodeResult_shift = laneRequestSourceWire_9_bits_decodeResult_shift;
  wire         validSource_9_bits_decodeResult_adder = laneRequestSourceWire_9_bits_decodeResult_adder;
  wire         validSource_9_bits_decodeResult_logic = laneRequestSourceWire_9_bits_decodeResult_logic;
  wire         validSource_9_bits_loadStore = laneRequestSourceWire_9_bits_loadStore;
  wire         validSource_9_bits_issueInst = laneRequestSourceWire_9_bits_issueInst;
  wire         validSource_9_bits_store = laneRequestSourceWire_9_bits_store;
  wire         validSource_9_bits_special = laneRequestSourceWire_9_bits_special;
  wire         validSource_9_bits_lsWholeReg = laneRequestSourceWire_9_bits_lsWholeReg;
  wire [4:0]   validSource_9_bits_vs1 = laneRequestSourceWire_9_bits_vs1;
  wire [4:0]   validSource_9_bits_vs2 = laneRequestSourceWire_9_bits_vs2;
  wire [4:0]   validSource_9_bits_vd = laneRequestSourceWire_9_bits_vd;
  wire [1:0]   validSource_9_bits_loadStoreEEW = laneRequestSourceWire_9_bits_loadStoreEEW;
  wire         validSource_9_bits_mask = laneRequestSourceWire_9_bits_mask;
  wire [2:0]   validSource_9_bits_segment = laneRequestSourceWire_9_bits_segment;
  wire [31:0]  validSource_9_bits_readFromScalar = laneRequestSourceWire_9_bits_readFromScalar;
  wire [11:0]  validSource_9_bits_csrInterface_vl = laneRequestSourceWire_9_bits_csrInterface_vl;
  wire [11:0]  validSource_9_bits_csrInterface_vStart = laneRequestSourceWire_9_bits_csrInterface_vStart;
  wire [2:0]   validSource_9_bits_csrInterface_vlmul = laneRequestSourceWire_9_bits_csrInterface_vlmul;
  wire [1:0]   validSource_9_bits_csrInterface_vSew = laneRequestSourceWire_9_bits_csrInterface_vSew;
  wire [1:0]   validSource_9_bits_csrInterface_vxrm = laneRequestSourceWire_9_bits_csrInterface_vxrm;
  wire         validSource_9_bits_csrInterface_vta = laneRequestSourceWire_9_bits_csrInterface_vta;
  wire         validSource_9_bits_csrInterface_vma = laneRequestSourceWire_9_bits_csrInterface_vma;
  wire         tokenCheck_10;
  wire [2:0]   validSource_10_bits_instructionIndex = laneRequestSourceWire_10_bits_instructionIndex;
  wire         validSource_10_bits_decodeResult_orderReduce = laneRequestSourceWire_10_bits_decodeResult_orderReduce;
  wire         validSource_10_bits_decodeResult_floatMul = laneRequestSourceWire_10_bits_decodeResult_floatMul;
  wire [1:0]   validSource_10_bits_decodeResult_fpExecutionType = laneRequestSourceWire_10_bits_decodeResult_fpExecutionType;
  wire         validSource_10_bits_decodeResult_float = laneRequestSourceWire_10_bits_decodeResult_float;
  wire         validSource_10_bits_decodeResult_specialSlot = laneRequestSourceWire_10_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_10_bits_decodeResult_topUop = laneRequestSourceWire_10_bits_decodeResult_topUop;
  wire         validSource_10_bits_decodeResult_popCount = laneRequestSourceWire_10_bits_decodeResult_popCount;
  wire         validSource_10_bits_decodeResult_ffo = laneRequestSourceWire_10_bits_decodeResult_ffo;
  wire         validSource_10_bits_decodeResult_average = laneRequestSourceWire_10_bits_decodeResult_average;
  wire         validSource_10_bits_decodeResult_reverse = laneRequestSourceWire_10_bits_decodeResult_reverse;
  wire         validSource_10_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_10_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_10_bits_decodeResult_scheduler = laneRequestSourceWire_10_bits_decodeResult_scheduler;
  wire         validSource_10_bits_decodeResult_sReadVD = laneRequestSourceWire_10_bits_decodeResult_sReadVD;
  wire         validSource_10_bits_decodeResult_vtype = laneRequestSourceWire_10_bits_decodeResult_vtype;
  wire         validSource_10_bits_decodeResult_sWrite = laneRequestSourceWire_10_bits_decodeResult_sWrite;
  wire         validSource_10_bits_decodeResult_crossRead = laneRequestSourceWire_10_bits_decodeResult_crossRead;
  wire         validSource_10_bits_decodeResult_crossWrite = laneRequestSourceWire_10_bits_decodeResult_crossWrite;
  wire         validSource_10_bits_decodeResult_maskUnit = laneRequestSourceWire_10_bits_decodeResult_maskUnit;
  wire         validSource_10_bits_decodeResult_special = laneRequestSourceWire_10_bits_decodeResult_special;
  wire         validSource_10_bits_decodeResult_saturate = laneRequestSourceWire_10_bits_decodeResult_saturate;
  wire         validSource_10_bits_decodeResult_vwmacc = laneRequestSourceWire_10_bits_decodeResult_vwmacc;
  wire         validSource_10_bits_decodeResult_readOnly = laneRequestSourceWire_10_bits_decodeResult_readOnly;
  wire         validSource_10_bits_decodeResult_maskSource = laneRequestSourceWire_10_bits_decodeResult_maskSource;
  wire         validSource_10_bits_decodeResult_maskDestination = laneRequestSourceWire_10_bits_decodeResult_maskDestination;
  wire         validSource_10_bits_decodeResult_maskLogic = laneRequestSourceWire_10_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_10_bits_decodeResult_uop = laneRequestSourceWire_10_bits_decodeResult_uop;
  wire         validSource_10_bits_decodeResult_iota = laneRequestSourceWire_10_bits_decodeResult_iota;
  wire         validSource_10_bits_decodeResult_mv = laneRequestSourceWire_10_bits_decodeResult_mv;
  wire         validSource_10_bits_decodeResult_extend = laneRequestSourceWire_10_bits_decodeResult_extend;
  wire         validSource_10_bits_decodeResult_unOrderWrite = laneRequestSourceWire_10_bits_decodeResult_unOrderWrite;
  wire         validSource_10_bits_decodeResult_compress = laneRequestSourceWire_10_bits_decodeResult_compress;
  wire         validSource_10_bits_decodeResult_gather16 = laneRequestSourceWire_10_bits_decodeResult_gather16;
  wire         validSource_10_bits_decodeResult_gather = laneRequestSourceWire_10_bits_decodeResult_gather;
  wire         validSource_10_bits_decodeResult_slid = laneRequestSourceWire_10_bits_decodeResult_slid;
  wire         validSource_10_bits_decodeResult_targetRd = laneRequestSourceWire_10_bits_decodeResult_targetRd;
  wire         validSource_10_bits_decodeResult_widenReduce = laneRequestSourceWire_10_bits_decodeResult_widenReduce;
  wire         validSource_10_bits_decodeResult_red = laneRequestSourceWire_10_bits_decodeResult_red;
  wire         validSource_10_bits_decodeResult_nr = laneRequestSourceWire_10_bits_decodeResult_nr;
  wire         validSource_10_bits_decodeResult_itype = laneRequestSourceWire_10_bits_decodeResult_itype;
  wire         validSource_10_bits_decodeResult_unsigned1 = laneRequestSourceWire_10_bits_decodeResult_unsigned1;
  wire         validSource_10_bits_decodeResult_unsigned0 = laneRequestSourceWire_10_bits_decodeResult_unsigned0;
  wire         validSource_10_bits_decodeResult_other = laneRequestSourceWire_10_bits_decodeResult_other;
  wire         validSource_10_bits_decodeResult_multiCycle = laneRequestSourceWire_10_bits_decodeResult_multiCycle;
  wire         validSource_10_bits_decodeResult_divider = laneRequestSourceWire_10_bits_decodeResult_divider;
  wire         validSource_10_bits_decodeResult_multiplier = laneRequestSourceWire_10_bits_decodeResult_multiplier;
  wire         validSource_10_bits_decodeResult_shift = laneRequestSourceWire_10_bits_decodeResult_shift;
  wire         validSource_10_bits_decodeResult_adder = laneRequestSourceWire_10_bits_decodeResult_adder;
  wire         validSource_10_bits_decodeResult_logic = laneRequestSourceWire_10_bits_decodeResult_logic;
  wire         validSource_10_bits_loadStore = laneRequestSourceWire_10_bits_loadStore;
  wire         validSource_10_bits_issueInst = laneRequestSourceWire_10_bits_issueInst;
  wire         validSource_10_bits_store = laneRequestSourceWire_10_bits_store;
  wire         validSource_10_bits_special = laneRequestSourceWire_10_bits_special;
  wire         validSource_10_bits_lsWholeReg = laneRequestSourceWire_10_bits_lsWholeReg;
  wire [4:0]   validSource_10_bits_vs1 = laneRequestSourceWire_10_bits_vs1;
  wire [4:0]   validSource_10_bits_vs2 = laneRequestSourceWire_10_bits_vs2;
  wire [4:0]   validSource_10_bits_vd = laneRequestSourceWire_10_bits_vd;
  wire [1:0]   validSource_10_bits_loadStoreEEW = laneRequestSourceWire_10_bits_loadStoreEEW;
  wire         validSource_10_bits_mask = laneRequestSourceWire_10_bits_mask;
  wire [2:0]   validSource_10_bits_segment = laneRequestSourceWire_10_bits_segment;
  wire [31:0]  validSource_10_bits_readFromScalar = laneRequestSourceWire_10_bits_readFromScalar;
  wire [11:0]  validSource_10_bits_csrInterface_vl = laneRequestSourceWire_10_bits_csrInterface_vl;
  wire [11:0]  validSource_10_bits_csrInterface_vStart = laneRequestSourceWire_10_bits_csrInterface_vStart;
  wire [2:0]   validSource_10_bits_csrInterface_vlmul = laneRequestSourceWire_10_bits_csrInterface_vlmul;
  wire [1:0]   validSource_10_bits_csrInterface_vSew = laneRequestSourceWire_10_bits_csrInterface_vSew;
  wire [1:0]   validSource_10_bits_csrInterface_vxrm = laneRequestSourceWire_10_bits_csrInterface_vxrm;
  wire         validSource_10_bits_csrInterface_vta = laneRequestSourceWire_10_bits_csrInterface_vta;
  wire         validSource_10_bits_csrInterface_vma = laneRequestSourceWire_10_bits_csrInterface_vma;
  wire         tokenCheck_11;
  wire [2:0]   validSource_11_bits_instructionIndex = laneRequestSourceWire_11_bits_instructionIndex;
  wire         validSource_11_bits_decodeResult_orderReduce = laneRequestSourceWire_11_bits_decodeResult_orderReduce;
  wire         validSource_11_bits_decodeResult_floatMul = laneRequestSourceWire_11_bits_decodeResult_floatMul;
  wire [1:0]   validSource_11_bits_decodeResult_fpExecutionType = laneRequestSourceWire_11_bits_decodeResult_fpExecutionType;
  wire         validSource_11_bits_decodeResult_float = laneRequestSourceWire_11_bits_decodeResult_float;
  wire         validSource_11_bits_decodeResult_specialSlot = laneRequestSourceWire_11_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_11_bits_decodeResult_topUop = laneRequestSourceWire_11_bits_decodeResult_topUop;
  wire         validSource_11_bits_decodeResult_popCount = laneRequestSourceWire_11_bits_decodeResult_popCount;
  wire         validSource_11_bits_decodeResult_ffo = laneRequestSourceWire_11_bits_decodeResult_ffo;
  wire         validSource_11_bits_decodeResult_average = laneRequestSourceWire_11_bits_decodeResult_average;
  wire         validSource_11_bits_decodeResult_reverse = laneRequestSourceWire_11_bits_decodeResult_reverse;
  wire         validSource_11_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_11_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_11_bits_decodeResult_scheduler = laneRequestSourceWire_11_bits_decodeResult_scheduler;
  wire         validSource_11_bits_decodeResult_sReadVD = laneRequestSourceWire_11_bits_decodeResult_sReadVD;
  wire         validSource_11_bits_decodeResult_vtype = laneRequestSourceWire_11_bits_decodeResult_vtype;
  wire         validSource_11_bits_decodeResult_sWrite = laneRequestSourceWire_11_bits_decodeResult_sWrite;
  wire         validSource_11_bits_decodeResult_crossRead = laneRequestSourceWire_11_bits_decodeResult_crossRead;
  wire         validSource_11_bits_decodeResult_crossWrite = laneRequestSourceWire_11_bits_decodeResult_crossWrite;
  wire         validSource_11_bits_decodeResult_maskUnit = laneRequestSourceWire_11_bits_decodeResult_maskUnit;
  wire         validSource_11_bits_decodeResult_special = laneRequestSourceWire_11_bits_decodeResult_special;
  wire         validSource_11_bits_decodeResult_saturate = laneRequestSourceWire_11_bits_decodeResult_saturate;
  wire         validSource_11_bits_decodeResult_vwmacc = laneRequestSourceWire_11_bits_decodeResult_vwmacc;
  wire         validSource_11_bits_decodeResult_readOnly = laneRequestSourceWire_11_bits_decodeResult_readOnly;
  wire         validSource_11_bits_decodeResult_maskSource = laneRequestSourceWire_11_bits_decodeResult_maskSource;
  wire         validSource_11_bits_decodeResult_maskDestination = laneRequestSourceWire_11_bits_decodeResult_maskDestination;
  wire         validSource_11_bits_decodeResult_maskLogic = laneRequestSourceWire_11_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_11_bits_decodeResult_uop = laneRequestSourceWire_11_bits_decodeResult_uop;
  wire         validSource_11_bits_decodeResult_iota = laneRequestSourceWire_11_bits_decodeResult_iota;
  wire         validSource_11_bits_decodeResult_mv = laneRequestSourceWire_11_bits_decodeResult_mv;
  wire         validSource_11_bits_decodeResult_extend = laneRequestSourceWire_11_bits_decodeResult_extend;
  wire         validSource_11_bits_decodeResult_unOrderWrite = laneRequestSourceWire_11_bits_decodeResult_unOrderWrite;
  wire         validSource_11_bits_decodeResult_compress = laneRequestSourceWire_11_bits_decodeResult_compress;
  wire         validSource_11_bits_decodeResult_gather16 = laneRequestSourceWire_11_bits_decodeResult_gather16;
  wire         validSource_11_bits_decodeResult_gather = laneRequestSourceWire_11_bits_decodeResult_gather;
  wire         validSource_11_bits_decodeResult_slid = laneRequestSourceWire_11_bits_decodeResult_slid;
  wire         validSource_11_bits_decodeResult_targetRd = laneRequestSourceWire_11_bits_decodeResult_targetRd;
  wire         validSource_11_bits_decodeResult_widenReduce = laneRequestSourceWire_11_bits_decodeResult_widenReduce;
  wire         validSource_11_bits_decodeResult_red = laneRequestSourceWire_11_bits_decodeResult_red;
  wire         validSource_11_bits_decodeResult_nr = laneRequestSourceWire_11_bits_decodeResult_nr;
  wire         validSource_11_bits_decodeResult_itype = laneRequestSourceWire_11_bits_decodeResult_itype;
  wire         validSource_11_bits_decodeResult_unsigned1 = laneRequestSourceWire_11_bits_decodeResult_unsigned1;
  wire         validSource_11_bits_decodeResult_unsigned0 = laneRequestSourceWire_11_bits_decodeResult_unsigned0;
  wire         validSource_11_bits_decodeResult_other = laneRequestSourceWire_11_bits_decodeResult_other;
  wire         validSource_11_bits_decodeResult_multiCycle = laneRequestSourceWire_11_bits_decodeResult_multiCycle;
  wire         validSource_11_bits_decodeResult_divider = laneRequestSourceWire_11_bits_decodeResult_divider;
  wire         validSource_11_bits_decodeResult_multiplier = laneRequestSourceWire_11_bits_decodeResult_multiplier;
  wire         validSource_11_bits_decodeResult_shift = laneRequestSourceWire_11_bits_decodeResult_shift;
  wire         validSource_11_bits_decodeResult_adder = laneRequestSourceWire_11_bits_decodeResult_adder;
  wire         validSource_11_bits_decodeResult_logic = laneRequestSourceWire_11_bits_decodeResult_logic;
  wire         validSource_11_bits_loadStore = laneRequestSourceWire_11_bits_loadStore;
  wire         validSource_11_bits_issueInst = laneRequestSourceWire_11_bits_issueInst;
  wire         validSource_11_bits_store = laneRequestSourceWire_11_bits_store;
  wire         validSource_11_bits_special = laneRequestSourceWire_11_bits_special;
  wire         validSource_11_bits_lsWholeReg = laneRequestSourceWire_11_bits_lsWholeReg;
  wire [4:0]   validSource_11_bits_vs1 = laneRequestSourceWire_11_bits_vs1;
  wire [4:0]   validSource_11_bits_vs2 = laneRequestSourceWire_11_bits_vs2;
  wire [4:0]   validSource_11_bits_vd = laneRequestSourceWire_11_bits_vd;
  wire [1:0]   validSource_11_bits_loadStoreEEW = laneRequestSourceWire_11_bits_loadStoreEEW;
  wire         validSource_11_bits_mask = laneRequestSourceWire_11_bits_mask;
  wire [2:0]   validSource_11_bits_segment = laneRequestSourceWire_11_bits_segment;
  wire [31:0]  validSource_11_bits_readFromScalar = laneRequestSourceWire_11_bits_readFromScalar;
  wire [11:0]  validSource_11_bits_csrInterface_vl = laneRequestSourceWire_11_bits_csrInterface_vl;
  wire [11:0]  validSource_11_bits_csrInterface_vStart = laneRequestSourceWire_11_bits_csrInterface_vStart;
  wire [2:0]   validSource_11_bits_csrInterface_vlmul = laneRequestSourceWire_11_bits_csrInterface_vlmul;
  wire [1:0]   validSource_11_bits_csrInterface_vSew = laneRequestSourceWire_11_bits_csrInterface_vSew;
  wire [1:0]   validSource_11_bits_csrInterface_vxrm = laneRequestSourceWire_11_bits_csrInterface_vxrm;
  wire         validSource_11_bits_csrInterface_vta = laneRequestSourceWire_11_bits_csrInterface_vta;
  wire         validSource_11_bits_csrInterface_vma = laneRequestSourceWire_11_bits_csrInterface_vma;
  wire         tokenCheck_12;
  wire [2:0]   validSource_12_bits_instructionIndex = laneRequestSourceWire_12_bits_instructionIndex;
  wire         validSource_12_bits_decodeResult_orderReduce = laneRequestSourceWire_12_bits_decodeResult_orderReduce;
  wire         validSource_12_bits_decodeResult_floatMul = laneRequestSourceWire_12_bits_decodeResult_floatMul;
  wire [1:0]   validSource_12_bits_decodeResult_fpExecutionType = laneRequestSourceWire_12_bits_decodeResult_fpExecutionType;
  wire         validSource_12_bits_decodeResult_float = laneRequestSourceWire_12_bits_decodeResult_float;
  wire         validSource_12_bits_decodeResult_specialSlot = laneRequestSourceWire_12_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_12_bits_decodeResult_topUop = laneRequestSourceWire_12_bits_decodeResult_topUop;
  wire         validSource_12_bits_decodeResult_popCount = laneRequestSourceWire_12_bits_decodeResult_popCount;
  wire         validSource_12_bits_decodeResult_ffo = laneRequestSourceWire_12_bits_decodeResult_ffo;
  wire         validSource_12_bits_decodeResult_average = laneRequestSourceWire_12_bits_decodeResult_average;
  wire         validSource_12_bits_decodeResult_reverse = laneRequestSourceWire_12_bits_decodeResult_reverse;
  wire         validSource_12_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_12_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_12_bits_decodeResult_scheduler = laneRequestSourceWire_12_bits_decodeResult_scheduler;
  wire         validSource_12_bits_decodeResult_sReadVD = laneRequestSourceWire_12_bits_decodeResult_sReadVD;
  wire         validSource_12_bits_decodeResult_vtype = laneRequestSourceWire_12_bits_decodeResult_vtype;
  wire         validSource_12_bits_decodeResult_sWrite = laneRequestSourceWire_12_bits_decodeResult_sWrite;
  wire         validSource_12_bits_decodeResult_crossRead = laneRequestSourceWire_12_bits_decodeResult_crossRead;
  wire         validSource_12_bits_decodeResult_crossWrite = laneRequestSourceWire_12_bits_decodeResult_crossWrite;
  wire         validSource_12_bits_decodeResult_maskUnit = laneRequestSourceWire_12_bits_decodeResult_maskUnit;
  wire         validSource_12_bits_decodeResult_special = laneRequestSourceWire_12_bits_decodeResult_special;
  wire         validSource_12_bits_decodeResult_saturate = laneRequestSourceWire_12_bits_decodeResult_saturate;
  wire         validSource_12_bits_decodeResult_vwmacc = laneRequestSourceWire_12_bits_decodeResult_vwmacc;
  wire         validSource_12_bits_decodeResult_readOnly = laneRequestSourceWire_12_bits_decodeResult_readOnly;
  wire         validSource_12_bits_decodeResult_maskSource = laneRequestSourceWire_12_bits_decodeResult_maskSource;
  wire         validSource_12_bits_decodeResult_maskDestination = laneRequestSourceWire_12_bits_decodeResult_maskDestination;
  wire         validSource_12_bits_decodeResult_maskLogic = laneRequestSourceWire_12_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_12_bits_decodeResult_uop = laneRequestSourceWire_12_bits_decodeResult_uop;
  wire         validSource_12_bits_decodeResult_iota = laneRequestSourceWire_12_bits_decodeResult_iota;
  wire         validSource_12_bits_decodeResult_mv = laneRequestSourceWire_12_bits_decodeResult_mv;
  wire         validSource_12_bits_decodeResult_extend = laneRequestSourceWire_12_bits_decodeResult_extend;
  wire         validSource_12_bits_decodeResult_unOrderWrite = laneRequestSourceWire_12_bits_decodeResult_unOrderWrite;
  wire         validSource_12_bits_decodeResult_compress = laneRequestSourceWire_12_bits_decodeResult_compress;
  wire         validSource_12_bits_decodeResult_gather16 = laneRequestSourceWire_12_bits_decodeResult_gather16;
  wire         validSource_12_bits_decodeResult_gather = laneRequestSourceWire_12_bits_decodeResult_gather;
  wire         validSource_12_bits_decodeResult_slid = laneRequestSourceWire_12_bits_decodeResult_slid;
  wire         validSource_12_bits_decodeResult_targetRd = laneRequestSourceWire_12_bits_decodeResult_targetRd;
  wire         validSource_12_bits_decodeResult_widenReduce = laneRequestSourceWire_12_bits_decodeResult_widenReduce;
  wire         validSource_12_bits_decodeResult_red = laneRequestSourceWire_12_bits_decodeResult_red;
  wire         validSource_12_bits_decodeResult_nr = laneRequestSourceWire_12_bits_decodeResult_nr;
  wire         validSource_12_bits_decodeResult_itype = laneRequestSourceWire_12_bits_decodeResult_itype;
  wire         validSource_12_bits_decodeResult_unsigned1 = laneRequestSourceWire_12_bits_decodeResult_unsigned1;
  wire         validSource_12_bits_decodeResult_unsigned0 = laneRequestSourceWire_12_bits_decodeResult_unsigned0;
  wire         validSource_12_bits_decodeResult_other = laneRequestSourceWire_12_bits_decodeResult_other;
  wire         validSource_12_bits_decodeResult_multiCycle = laneRequestSourceWire_12_bits_decodeResult_multiCycle;
  wire         validSource_12_bits_decodeResult_divider = laneRequestSourceWire_12_bits_decodeResult_divider;
  wire         validSource_12_bits_decodeResult_multiplier = laneRequestSourceWire_12_bits_decodeResult_multiplier;
  wire         validSource_12_bits_decodeResult_shift = laneRequestSourceWire_12_bits_decodeResult_shift;
  wire         validSource_12_bits_decodeResult_adder = laneRequestSourceWire_12_bits_decodeResult_adder;
  wire         validSource_12_bits_decodeResult_logic = laneRequestSourceWire_12_bits_decodeResult_logic;
  wire         validSource_12_bits_loadStore = laneRequestSourceWire_12_bits_loadStore;
  wire         validSource_12_bits_issueInst = laneRequestSourceWire_12_bits_issueInst;
  wire         validSource_12_bits_store = laneRequestSourceWire_12_bits_store;
  wire         validSource_12_bits_special = laneRequestSourceWire_12_bits_special;
  wire         validSource_12_bits_lsWholeReg = laneRequestSourceWire_12_bits_lsWholeReg;
  wire [4:0]   validSource_12_bits_vs1 = laneRequestSourceWire_12_bits_vs1;
  wire [4:0]   validSource_12_bits_vs2 = laneRequestSourceWire_12_bits_vs2;
  wire [4:0]   validSource_12_bits_vd = laneRequestSourceWire_12_bits_vd;
  wire [1:0]   validSource_12_bits_loadStoreEEW = laneRequestSourceWire_12_bits_loadStoreEEW;
  wire         validSource_12_bits_mask = laneRequestSourceWire_12_bits_mask;
  wire [2:0]   validSource_12_bits_segment = laneRequestSourceWire_12_bits_segment;
  wire [31:0]  validSource_12_bits_readFromScalar = laneRequestSourceWire_12_bits_readFromScalar;
  wire [11:0]  validSource_12_bits_csrInterface_vl = laneRequestSourceWire_12_bits_csrInterface_vl;
  wire [11:0]  validSource_12_bits_csrInterface_vStart = laneRequestSourceWire_12_bits_csrInterface_vStart;
  wire [2:0]   validSource_12_bits_csrInterface_vlmul = laneRequestSourceWire_12_bits_csrInterface_vlmul;
  wire [1:0]   validSource_12_bits_csrInterface_vSew = laneRequestSourceWire_12_bits_csrInterface_vSew;
  wire [1:0]   validSource_12_bits_csrInterface_vxrm = laneRequestSourceWire_12_bits_csrInterface_vxrm;
  wire         validSource_12_bits_csrInterface_vta = laneRequestSourceWire_12_bits_csrInterface_vta;
  wire         validSource_12_bits_csrInterface_vma = laneRequestSourceWire_12_bits_csrInterface_vma;
  wire         tokenCheck_13;
  wire [2:0]   validSource_13_bits_instructionIndex = laneRequestSourceWire_13_bits_instructionIndex;
  wire         validSource_13_bits_decodeResult_orderReduce = laneRequestSourceWire_13_bits_decodeResult_orderReduce;
  wire         validSource_13_bits_decodeResult_floatMul = laneRequestSourceWire_13_bits_decodeResult_floatMul;
  wire [1:0]   validSource_13_bits_decodeResult_fpExecutionType = laneRequestSourceWire_13_bits_decodeResult_fpExecutionType;
  wire         validSource_13_bits_decodeResult_float = laneRequestSourceWire_13_bits_decodeResult_float;
  wire         validSource_13_bits_decodeResult_specialSlot = laneRequestSourceWire_13_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_13_bits_decodeResult_topUop = laneRequestSourceWire_13_bits_decodeResult_topUop;
  wire         validSource_13_bits_decodeResult_popCount = laneRequestSourceWire_13_bits_decodeResult_popCount;
  wire         validSource_13_bits_decodeResult_ffo = laneRequestSourceWire_13_bits_decodeResult_ffo;
  wire         validSource_13_bits_decodeResult_average = laneRequestSourceWire_13_bits_decodeResult_average;
  wire         validSource_13_bits_decodeResult_reverse = laneRequestSourceWire_13_bits_decodeResult_reverse;
  wire         validSource_13_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_13_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_13_bits_decodeResult_scheduler = laneRequestSourceWire_13_bits_decodeResult_scheduler;
  wire         validSource_13_bits_decodeResult_sReadVD = laneRequestSourceWire_13_bits_decodeResult_sReadVD;
  wire         validSource_13_bits_decodeResult_vtype = laneRequestSourceWire_13_bits_decodeResult_vtype;
  wire         validSource_13_bits_decodeResult_sWrite = laneRequestSourceWire_13_bits_decodeResult_sWrite;
  wire         validSource_13_bits_decodeResult_crossRead = laneRequestSourceWire_13_bits_decodeResult_crossRead;
  wire         validSource_13_bits_decodeResult_crossWrite = laneRequestSourceWire_13_bits_decodeResult_crossWrite;
  wire         validSource_13_bits_decodeResult_maskUnit = laneRequestSourceWire_13_bits_decodeResult_maskUnit;
  wire         validSource_13_bits_decodeResult_special = laneRequestSourceWire_13_bits_decodeResult_special;
  wire         validSource_13_bits_decodeResult_saturate = laneRequestSourceWire_13_bits_decodeResult_saturate;
  wire         validSource_13_bits_decodeResult_vwmacc = laneRequestSourceWire_13_bits_decodeResult_vwmacc;
  wire         validSource_13_bits_decodeResult_readOnly = laneRequestSourceWire_13_bits_decodeResult_readOnly;
  wire         validSource_13_bits_decodeResult_maskSource = laneRequestSourceWire_13_bits_decodeResult_maskSource;
  wire         validSource_13_bits_decodeResult_maskDestination = laneRequestSourceWire_13_bits_decodeResult_maskDestination;
  wire         validSource_13_bits_decodeResult_maskLogic = laneRequestSourceWire_13_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_13_bits_decodeResult_uop = laneRequestSourceWire_13_bits_decodeResult_uop;
  wire         validSource_13_bits_decodeResult_iota = laneRequestSourceWire_13_bits_decodeResult_iota;
  wire         validSource_13_bits_decodeResult_mv = laneRequestSourceWire_13_bits_decodeResult_mv;
  wire         validSource_13_bits_decodeResult_extend = laneRequestSourceWire_13_bits_decodeResult_extend;
  wire         validSource_13_bits_decodeResult_unOrderWrite = laneRequestSourceWire_13_bits_decodeResult_unOrderWrite;
  wire         validSource_13_bits_decodeResult_compress = laneRequestSourceWire_13_bits_decodeResult_compress;
  wire         validSource_13_bits_decodeResult_gather16 = laneRequestSourceWire_13_bits_decodeResult_gather16;
  wire         validSource_13_bits_decodeResult_gather = laneRequestSourceWire_13_bits_decodeResult_gather;
  wire         validSource_13_bits_decodeResult_slid = laneRequestSourceWire_13_bits_decodeResult_slid;
  wire         validSource_13_bits_decodeResult_targetRd = laneRequestSourceWire_13_bits_decodeResult_targetRd;
  wire         validSource_13_bits_decodeResult_widenReduce = laneRequestSourceWire_13_bits_decodeResult_widenReduce;
  wire         validSource_13_bits_decodeResult_red = laneRequestSourceWire_13_bits_decodeResult_red;
  wire         validSource_13_bits_decodeResult_nr = laneRequestSourceWire_13_bits_decodeResult_nr;
  wire         validSource_13_bits_decodeResult_itype = laneRequestSourceWire_13_bits_decodeResult_itype;
  wire         validSource_13_bits_decodeResult_unsigned1 = laneRequestSourceWire_13_bits_decodeResult_unsigned1;
  wire         validSource_13_bits_decodeResult_unsigned0 = laneRequestSourceWire_13_bits_decodeResult_unsigned0;
  wire         validSource_13_bits_decodeResult_other = laneRequestSourceWire_13_bits_decodeResult_other;
  wire         validSource_13_bits_decodeResult_multiCycle = laneRequestSourceWire_13_bits_decodeResult_multiCycle;
  wire         validSource_13_bits_decodeResult_divider = laneRequestSourceWire_13_bits_decodeResult_divider;
  wire         validSource_13_bits_decodeResult_multiplier = laneRequestSourceWire_13_bits_decodeResult_multiplier;
  wire         validSource_13_bits_decodeResult_shift = laneRequestSourceWire_13_bits_decodeResult_shift;
  wire         validSource_13_bits_decodeResult_adder = laneRequestSourceWire_13_bits_decodeResult_adder;
  wire         validSource_13_bits_decodeResult_logic = laneRequestSourceWire_13_bits_decodeResult_logic;
  wire         validSource_13_bits_loadStore = laneRequestSourceWire_13_bits_loadStore;
  wire         validSource_13_bits_issueInst = laneRequestSourceWire_13_bits_issueInst;
  wire         validSource_13_bits_store = laneRequestSourceWire_13_bits_store;
  wire         validSource_13_bits_special = laneRequestSourceWire_13_bits_special;
  wire         validSource_13_bits_lsWholeReg = laneRequestSourceWire_13_bits_lsWholeReg;
  wire [4:0]   validSource_13_bits_vs1 = laneRequestSourceWire_13_bits_vs1;
  wire [4:0]   validSource_13_bits_vs2 = laneRequestSourceWire_13_bits_vs2;
  wire [4:0]   validSource_13_bits_vd = laneRequestSourceWire_13_bits_vd;
  wire [1:0]   validSource_13_bits_loadStoreEEW = laneRequestSourceWire_13_bits_loadStoreEEW;
  wire         validSource_13_bits_mask = laneRequestSourceWire_13_bits_mask;
  wire [2:0]   validSource_13_bits_segment = laneRequestSourceWire_13_bits_segment;
  wire [31:0]  validSource_13_bits_readFromScalar = laneRequestSourceWire_13_bits_readFromScalar;
  wire [11:0]  validSource_13_bits_csrInterface_vl = laneRequestSourceWire_13_bits_csrInterface_vl;
  wire [11:0]  validSource_13_bits_csrInterface_vStart = laneRequestSourceWire_13_bits_csrInterface_vStart;
  wire [2:0]   validSource_13_bits_csrInterface_vlmul = laneRequestSourceWire_13_bits_csrInterface_vlmul;
  wire [1:0]   validSource_13_bits_csrInterface_vSew = laneRequestSourceWire_13_bits_csrInterface_vSew;
  wire [1:0]   validSource_13_bits_csrInterface_vxrm = laneRequestSourceWire_13_bits_csrInterface_vxrm;
  wire         validSource_13_bits_csrInterface_vta = laneRequestSourceWire_13_bits_csrInterface_vta;
  wire         validSource_13_bits_csrInterface_vma = laneRequestSourceWire_13_bits_csrInterface_vma;
  wire         tokenCheck_14;
  wire [2:0]   validSource_14_bits_instructionIndex = laneRequestSourceWire_14_bits_instructionIndex;
  wire         validSource_14_bits_decodeResult_orderReduce = laneRequestSourceWire_14_bits_decodeResult_orderReduce;
  wire         validSource_14_bits_decodeResult_floatMul = laneRequestSourceWire_14_bits_decodeResult_floatMul;
  wire [1:0]   validSource_14_bits_decodeResult_fpExecutionType = laneRequestSourceWire_14_bits_decodeResult_fpExecutionType;
  wire         validSource_14_bits_decodeResult_float = laneRequestSourceWire_14_bits_decodeResult_float;
  wire         validSource_14_bits_decodeResult_specialSlot = laneRequestSourceWire_14_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_14_bits_decodeResult_topUop = laneRequestSourceWire_14_bits_decodeResult_topUop;
  wire         validSource_14_bits_decodeResult_popCount = laneRequestSourceWire_14_bits_decodeResult_popCount;
  wire         validSource_14_bits_decodeResult_ffo = laneRequestSourceWire_14_bits_decodeResult_ffo;
  wire         validSource_14_bits_decodeResult_average = laneRequestSourceWire_14_bits_decodeResult_average;
  wire         validSource_14_bits_decodeResult_reverse = laneRequestSourceWire_14_bits_decodeResult_reverse;
  wire         validSource_14_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_14_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_14_bits_decodeResult_scheduler = laneRequestSourceWire_14_bits_decodeResult_scheduler;
  wire         validSource_14_bits_decodeResult_sReadVD = laneRequestSourceWire_14_bits_decodeResult_sReadVD;
  wire         validSource_14_bits_decodeResult_vtype = laneRequestSourceWire_14_bits_decodeResult_vtype;
  wire         validSource_14_bits_decodeResult_sWrite = laneRequestSourceWire_14_bits_decodeResult_sWrite;
  wire         validSource_14_bits_decodeResult_crossRead = laneRequestSourceWire_14_bits_decodeResult_crossRead;
  wire         validSource_14_bits_decodeResult_crossWrite = laneRequestSourceWire_14_bits_decodeResult_crossWrite;
  wire         validSource_14_bits_decodeResult_maskUnit = laneRequestSourceWire_14_bits_decodeResult_maskUnit;
  wire         validSource_14_bits_decodeResult_special = laneRequestSourceWire_14_bits_decodeResult_special;
  wire         validSource_14_bits_decodeResult_saturate = laneRequestSourceWire_14_bits_decodeResult_saturate;
  wire         validSource_14_bits_decodeResult_vwmacc = laneRequestSourceWire_14_bits_decodeResult_vwmacc;
  wire         validSource_14_bits_decodeResult_readOnly = laneRequestSourceWire_14_bits_decodeResult_readOnly;
  wire         validSource_14_bits_decodeResult_maskSource = laneRequestSourceWire_14_bits_decodeResult_maskSource;
  wire         validSource_14_bits_decodeResult_maskDestination = laneRequestSourceWire_14_bits_decodeResult_maskDestination;
  wire         validSource_14_bits_decodeResult_maskLogic = laneRequestSourceWire_14_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_14_bits_decodeResult_uop = laneRequestSourceWire_14_bits_decodeResult_uop;
  wire         validSource_14_bits_decodeResult_iota = laneRequestSourceWire_14_bits_decodeResult_iota;
  wire         validSource_14_bits_decodeResult_mv = laneRequestSourceWire_14_bits_decodeResult_mv;
  wire         validSource_14_bits_decodeResult_extend = laneRequestSourceWire_14_bits_decodeResult_extend;
  wire         validSource_14_bits_decodeResult_unOrderWrite = laneRequestSourceWire_14_bits_decodeResult_unOrderWrite;
  wire         validSource_14_bits_decodeResult_compress = laneRequestSourceWire_14_bits_decodeResult_compress;
  wire         validSource_14_bits_decodeResult_gather16 = laneRequestSourceWire_14_bits_decodeResult_gather16;
  wire         validSource_14_bits_decodeResult_gather = laneRequestSourceWire_14_bits_decodeResult_gather;
  wire         validSource_14_bits_decodeResult_slid = laneRequestSourceWire_14_bits_decodeResult_slid;
  wire         validSource_14_bits_decodeResult_targetRd = laneRequestSourceWire_14_bits_decodeResult_targetRd;
  wire         validSource_14_bits_decodeResult_widenReduce = laneRequestSourceWire_14_bits_decodeResult_widenReduce;
  wire         validSource_14_bits_decodeResult_red = laneRequestSourceWire_14_bits_decodeResult_red;
  wire         validSource_14_bits_decodeResult_nr = laneRequestSourceWire_14_bits_decodeResult_nr;
  wire         validSource_14_bits_decodeResult_itype = laneRequestSourceWire_14_bits_decodeResult_itype;
  wire         validSource_14_bits_decodeResult_unsigned1 = laneRequestSourceWire_14_bits_decodeResult_unsigned1;
  wire         validSource_14_bits_decodeResult_unsigned0 = laneRequestSourceWire_14_bits_decodeResult_unsigned0;
  wire         validSource_14_bits_decodeResult_other = laneRequestSourceWire_14_bits_decodeResult_other;
  wire         validSource_14_bits_decodeResult_multiCycle = laneRequestSourceWire_14_bits_decodeResult_multiCycle;
  wire         validSource_14_bits_decodeResult_divider = laneRequestSourceWire_14_bits_decodeResult_divider;
  wire         validSource_14_bits_decodeResult_multiplier = laneRequestSourceWire_14_bits_decodeResult_multiplier;
  wire         validSource_14_bits_decodeResult_shift = laneRequestSourceWire_14_bits_decodeResult_shift;
  wire         validSource_14_bits_decodeResult_adder = laneRequestSourceWire_14_bits_decodeResult_adder;
  wire         validSource_14_bits_decodeResult_logic = laneRequestSourceWire_14_bits_decodeResult_logic;
  wire         validSource_14_bits_loadStore = laneRequestSourceWire_14_bits_loadStore;
  wire         validSource_14_bits_issueInst = laneRequestSourceWire_14_bits_issueInst;
  wire         validSource_14_bits_store = laneRequestSourceWire_14_bits_store;
  wire         validSource_14_bits_special = laneRequestSourceWire_14_bits_special;
  wire         validSource_14_bits_lsWholeReg = laneRequestSourceWire_14_bits_lsWholeReg;
  wire [4:0]   validSource_14_bits_vs1 = laneRequestSourceWire_14_bits_vs1;
  wire [4:0]   validSource_14_bits_vs2 = laneRequestSourceWire_14_bits_vs2;
  wire [4:0]   validSource_14_bits_vd = laneRequestSourceWire_14_bits_vd;
  wire [1:0]   validSource_14_bits_loadStoreEEW = laneRequestSourceWire_14_bits_loadStoreEEW;
  wire         validSource_14_bits_mask = laneRequestSourceWire_14_bits_mask;
  wire [2:0]   validSource_14_bits_segment = laneRequestSourceWire_14_bits_segment;
  wire [31:0]  validSource_14_bits_readFromScalar = laneRequestSourceWire_14_bits_readFromScalar;
  wire [11:0]  validSource_14_bits_csrInterface_vl = laneRequestSourceWire_14_bits_csrInterface_vl;
  wire [11:0]  validSource_14_bits_csrInterface_vStart = laneRequestSourceWire_14_bits_csrInterface_vStart;
  wire [2:0]   validSource_14_bits_csrInterface_vlmul = laneRequestSourceWire_14_bits_csrInterface_vlmul;
  wire [1:0]   validSource_14_bits_csrInterface_vSew = laneRequestSourceWire_14_bits_csrInterface_vSew;
  wire [1:0]   validSource_14_bits_csrInterface_vxrm = laneRequestSourceWire_14_bits_csrInterface_vxrm;
  wire         validSource_14_bits_csrInterface_vta = laneRequestSourceWire_14_bits_csrInterface_vta;
  wire         validSource_14_bits_csrInterface_vma = laneRequestSourceWire_14_bits_csrInterface_vma;
  wire         tokenCheck_15;
  wire [2:0]   validSource_15_bits_instructionIndex = laneRequestSourceWire_15_bits_instructionIndex;
  wire         validSource_15_bits_decodeResult_orderReduce = laneRequestSourceWire_15_bits_decodeResult_orderReduce;
  wire         validSource_15_bits_decodeResult_floatMul = laneRequestSourceWire_15_bits_decodeResult_floatMul;
  wire [1:0]   validSource_15_bits_decodeResult_fpExecutionType = laneRequestSourceWire_15_bits_decodeResult_fpExecutionType;
  wire         validSource_15_bits_decodeResult_float = laneRequestSourceWire_15_bits_decodeResult_float;
  wire         validSource_15_bits_decodeResult_specialSlot = laneRequestSourceWire_15_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_15_bits_decodeResult_topUop = laneRequestSourceWire_15_bits_decodeResult_topUop;
  wire         validSource_15_bits_decodeResult_popCount = laneRequestSourceWire_15_bits_decodeResult_popCount;
  wire         validSource_15_bits_decodeResult_ffo = laneRequestSourceWire_15_bits_decodeResult_ffo;
  wire         validSource_15_bits_decodeResult_average = laneRequestSourceWire_15_bits_decodeResult_average;
  wire         validSource_15_bits_decodeResult_reverse = laneRequestSourceWire_15_bits_decodeResult_reverse;
  wire         validSource_15_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_15_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_15_bits_decodeResult_scheduler = laneRequestSourceWire_15_bits_decodeResult_scheduler;
  wire         validSource_15_bits_decodeResult_sReadVD = laneRequestSourceWire_15_bits_decodeResult_sReadVD;
  wire         validSource_15_bits_decodeResult_vtype = laneRequestSourceWire_15_bits_decodeResult_vtype;
  wire         validSource_15_bits_decodeResult_sWrite = laneRequestSourceWire_15_bits_decodeResult_sWrite;
  wire         validSource_15_bits_decodeResult_crossRead = laneRequestSourceWire_15_bits_decodeResult_crossRead;
  wire         validSource_15_bits_decodeResult_crossWrite = laneRequestSourceWire_15_bits_decodeResult_crossWrite;
  wire         validSource_15_bits_decodeResult_maskUnit = laneRequestSourceWire_15_bits_decodeResult_maskUnit;
  wire         validSource_15_bits_decodeResult_special = laneRequestSourceWire_15_bits_decodeResult_special;
  wire         validSource_15_bits_decodeResult_saturate = laneRequestSourceWire_15_bits_decodeResult_saturate;
  wire         validSource_15_bits_decodeResult_vwmacc = laneRequestSourceWire_15_bits_decodeResult_vwmacc;
  wire         validSource_15_bits_decodeResult_readOnly = laneRequestSourceWire_15_bits_decodeResult_readOnly;
  wire         validSource_15_bits_decodeResult_maskSource = laneRequestSourceWire_15_bits_decodeResult_maskSource;
  wire         validSource_15_bits_decodeResult_maskDestination = laneRequestSourceWire_15_bits_decodeResult_maskDestination;
  wire         validSource_15_bits_decodeResult_maskLogic = laneRequestSourceWire_15_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_15_bits_decodeResult_uop = laneRequestSourceWire_15_bits_decodeResult_uop;
  wire         validSource_15_bits_decodeResult_iota = laneRequestSourceWire_15_bits_decodeResult_iota;
  wire         validSource_15_bits_decodeResult_mv = laneRequestSourceWire_15_bits_decodeResult_mv;
  wire         validSource_15_bits_decodeResult_extend = laneRequestSourceWire_15_bits_decodeResult_extend;
  wire         validSource_15_bits_decodeResult_unOrderWrite = laneRequestSourceWire_15_bits_decodeResult_unOrderWrite;
  wire         validSource_15_bits_decodeResult_compress = laneRequestSourceWire_15_bits_decodeResult_compress;
  wire         validSource_15_bits_decodeResult_gather16 = laneRequestSourceWire_15_bits_decodeResult_gather16;
  wire         validSource_15_bits_decodeResult_gather = laneRequestSourceWire_15_bits_decodeResult_gather;
  wire         validSource_15_bits_decodeResult_slid = laneRequestSourceWire_15_bits_decodeResult_slid;
  wire         validSource_15_bits_decodeResult_targetRd = laneRequestSourceWire_15_bits_decodeResult_targetRd;
  wire         validSource_15_bits_decodeResult_widenReduce = laneRequestSourceWire_15_bits_decodeResult_widenReduce;
  wire         validSource_15_bits_decodeResult_red = laneRequestSourceWire_15_bits_decodeResult_red;
  wire         validSource_15_bits_decodeResult_nr = laneRequestSourceWire_15_bits_decodeResult_nr;
  wire         validSource_15_bits_decodeResult_itype = laneRequestSourceWire_15_bits_decodeResult_itype;
  wire         validSource_15_bits_decodeResult_unsigned1 = laneRequestSourceWire_15_bits_decodeResult_unsigned1;
  wire         validSource_15_bits_decodeResult_unsigned0 = laneRequestSourceWire_15_bits_decodeResult_unsigned0;
  wire         validSource_15_bits_decodeResult_other = laneRequestSourceWire_15_bits_decodeResult_other;
  wire         validSource_15_bits_decodeResult_multiCycle = laneRequestSourceWire_15_bits_decodeResult_multiCycle;
  wire         validSource_15_bits_decodeResult_divider = laneRequestSourceWire_15_bits_decodeResult_divider;
  wire         validSource_15_bits_decodeResult_multiplier = laneRequestSourceWire_15_bits_decodeResult_multiplier;
  wire         validSource_15_bits_decodeResult_shift = laneRequestSourceWire_15_bits_decodeResult_shift;
  wire         validSource_15_bits_decodeResult_adder = laneRequestSourceWire_15_bits_decodeResult_adder;
  wire         validSource_15_bits_decodeResult_logic = laneRequestSourceWire_15_bits_decodeResult_logic;
  wire         validSource_15_bits_loadStore = laneRequestSourceWire_15_bits_loadStore;
  wire         validSource_15_bits_issueInst = laneRequestSourceWire_15_bits_issueInst;
  wire         validSource_15_bits_store = laneRequestSourceWire_15_bits_store;
  wire         validSource_15_bits_special = laneRequestSourceWire_15_bits_special;
  wire         validSource_15_bits_lsWholeReg = laneRequestSourceWire_15_bits_lsWholeReg;
  wire [4:0]   validSource_15_bits_vs1 = laneRequestSourceWire_15_bits_vs1;
  wire [4:0]   validSource_15_bits_vs2 = laneRequestSourceWire_15_bits_vs2;
  wire [4:0]   validSource_15_bits_vd = laneRequestSourceWire_15_bits_vd;
  wire [1:0]   validSource_15_bits_loadStoreEEW = laneRequestSourceWire_15_bits_loadStoreEEW;
  wire         validSource_15_bits_mask = laneRequestSourceWire_15_bits_mask;
  wire [2:0]   validSource_15_bits_segment = laneRequestSourceWire_15_bits_segment;
  wire [31:0]  validSource_15_bits_readFromScalar = laneRequestSourceWire_15_bits_readFromScalar;
  wire [11:0]  validSource_15_bits_csrInterface_vl = laneRequestSourceWire_15_bits_csrInterface_vl;
  wire [11:0]  validSource_15_bits_csrInterface_vStart = laneRequestSourceWire_15_bits_csrInterface_vStart;
  wire [2:0]   validSource_15_bits_csrInterface_vlmul = laneRequestSourceWire_15_bits_csrInterface_vlmul;
  wire [1:0]   validSource_15_bits_csrInterface_vSew = laneRequestSourceWire_15_bits_csrInterface_vSew;
  wire [1:0]   validSource_15_bits_csrInterface_vxrm = laneRequestSourceWire_15_bits_csrInterface_vxrm;
  wire         validSource_15_bits_csrInterface_vta = laneRequestSourceWire_15_bits_csrInterface_vta;
  wire         validSource_15_bits_csrInterface_vma = laneRequestSourceWire_15_bits_csrInterface_vma;
  wire         queue_deq_ready = laneRequestSinkWire_0_ready;
  wire         queue_deq_valid;
  wire [2:0]   queue_deq_bits_instructionIndex;
  wire         queue_deq_bits_decodeResult_orderReduce;
  wire         queue_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_deq_bits_decodeResult_fpExecutionType;
  wire         queue_deq_bits_decodeResult_float;
  wire         queue_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_deq_bits_decodeResult_topUop;
  wire         queue_deq_bits_decodeResult_popCount;
  wire         queue_deq_bits_decodeResult_ffo;
  wire         queue_deq_bits_decodeResult_average;
  wire         queue_deq_bits_decodeResult_reverse;
  wire         queue_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_deq_bits_decodeResult_scheduler;
  wire         queue_deq_bits_decodeResult_sReadVD;
  wire         queue_deq_bits_decodeResult_vtype;
  wire         queue_deq_bits_decodeResult_sWrite;
  wire         queue_deq_bits_decodeResult_crossRead;
  wire         queue_deq_bits_decodeResult_crossWrite;
  wire         queue_deq_bits_decodeResult_maskUnit;
  wire         queue_deq_bits_decodeResult_special;
  wire         queue_deq_bits_decodeResult_saturate;
  wire         queue_deq_bits_decodeResult_vwmacc;
  wire         queue_deq_bits_decodeResult_readOnly;
  wire         queue_deq_bits_decodeResult_maskSource;
  wire         queue_deq_bits_decodeResult_maskDestination;
  wire         queue_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_deq_bits_decodeResult_uop;
  wire         queue_deq_bits_decodeResult_iota;
  wire         queue_deq_bits_decodeResult_mv;
  wire         queue_deq_bits_decodeResult_extend;
  wire         queue_deq_bits_decodeResult_unOrderWrite;
  wire         queue_deq_bits_decodeResult_compress;
  wire         queue_deq_bits_decodeResult_gather16;
  wire         queue_deq_bits_decodeResult_gather;
  wire         queue_deq_bits_decodeResult_slid;
  wire         queue_deq_bits_decodeResult_targetRd;
  wire         queue_deq_bits_decodeResult_widenReduce;
  wire         queue_deq_bits_decodeResult_red;
  wire         queue_deq_bits_decodeResult_nr;
  wire         queue_deq_bits_decodeResult_itype;
  wire         queue_deq_bits_decodeResult_unsigned1;
  wire         queue_deq_bits_decodeResult_unsigned0;
  wire         queue_deq_bits_decodeResult_other;
  wire         queue_deq_bits_decodeResult_multiCycle;
  wire         queue_deq_bits_decodeResult_divider;
  wire         queue_deq_bits_decodeResult_multiplier;
  wire         queue_deq_bits_decodeResult_shift;
  wire         queue_deq_bits_decodeResult_adder;
  wire         queue_deq_bits_decodeResult_logic;
  wire         queue_deq_bits_loadStore;
  wire         queue_deq_bits_issueInst;
  wire         queue_deq_bits_store;
  wire         queue_deq_bits_special;
  wire         queue_deq_bits_lsWholeReg;
  wire [4:0]   queue_deq_bits_vs1;
  wire [4:0]   queue_deq_bits_vs2;
  wire [4:0]   queue_deq_bits_vd;
  wire [1:0]   queue_deq_bits_loadStoreEEW;
  wire         queue_deq_bits_mask;
  wire [2:0]   queue_deq_bits_segment;
  wire [31:0]  queue_deq_bits_readFromScalar;
  wire [11:0]  queue_deq_bits_csrInterface_vl;
  wire [11:0]  queue_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_deq_bits_csrInterface_vxrm;
  wire         queue_deq_bits_csrInterface_vta;
  wire         queue_deq_bits_csrInterface_vma;
  wire         queue_1_deq_ready = laneRequestSinkWire_1_ready;
  wire         queue_1_deq_valid;
  wire [2:0]   queue_1_deq_bits_instructionIndex;
  wire         queue_1_deq_bits_decodeResult_orderReduce;
  wire         queue_1_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_1_deq_bits_decodeResult_fpExecutionType;
  wire         queue_1_deq_bits_decodeResult_float;
  wire         queue_1_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_1_deq_bits_decodeResult_topUop;
  wire         queue_1_deq_bits_decodeResult_popCount;
  wire         queue_1_deq_bits_decodeResult_ffo;
  wire         queue_1_deq_bits_decodeResult_average;
  wire         queue_1_deq_bits_decodeResult_reverse;
  wire         queue_1_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_1_deq_bits_decodeResult_scheduler;
  wire         queue_1_deq_bits_decodeResult_sReadVD;
  wire         queue_1_deq_bits_decodeResult_vtype;
  wire         queue_1_deq_bits_decodeResult_sWrite;
  wire         queue_1_deq_bits_decodeResult_crossRead;
  wire         queue_1_deq_bits_decodeResult_crossWrite;
  wire         queue_1_deq_bits_decodeResult_maskUnit;
  wire         queue_1_deq_bits_decodeResult_special;
  wire         queue_1_deq_bits_decodeResult_saturate;
  wire         queue_1_deq_bits_decodeResult_vwmacc;
  wire         queue_1_deq_bits_decodeResult_readOnly;
  wire         queue_1_deq_bits_decodeResult_maskSource;
  wire         queue_1_deq_bits_decodeResult_maskDestination;
  wire         queue_1_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_1_deq_bits_decodeResult_uop;
  wire         queue_1_deq_bits_decodeResult_iota;
  wire         queue_1_deq_bits_decodeResult_mv;
  wire         queue_1_deq_bits_decodeResult_extend;
  wire         queue_1_deq_bits_decodeResult_unOrderWrite;
  wire         queue_1_deq_bits_decodeResult_compress;
  wire         queue_1_deq_bits_decodeResult_gather16;
  wire         queue_1_deq_bits_decodeResult_gather;
  wire         queue_1_deq_bits_decodeResult_slid;
  wire         queue_1_deq_bits_decodeResult_targetRd;
  wire         queue_1_deq_bits_decodeResult_widenReduce;
  wire         queue_1_deq_bits_decodeResult_red;
  wire         queue_1_deq_bits_decodeResult_nr;
  wire         queue_1_deq_bits_decodeResult_itype;
  wire         queue_1_deq_bits_decodeResult_unsigned1;
  wire         queue_1_deq_bits_decodeResult_unsigned0;
  wire         queue_1_deq_bits_decodeResult_other;
  wire         queue_1_deq_bits_decodeResult_multiCycle;
  wire         queue_1_deq_bits_decodeResult_divider;
  wire         queue_1_deq_bits_decodeResult_multiplier;
  wire         queue_1_deq_bits_decodeResult_shift;
  wire         queue_1_deq_bits_decodeResult_adder;
  wire         queue_1_deq_bits_decodeResult_logic;
  wire         queue_1_deq_bits_loadStore;
  wire         queue_1_deq_bits_issueInst;
  wire         queue_1_deq_bits_store;
  wire         queue_1_deq_bits_special;
  wire         queue_1_deq_bits_lsWholeReg;
  wire [4:0]   queue_1_deq_bits_vs1;
  wire [4:0]   queue_1_deq_bits_vs2;
  wire [4:0]   queue_1_deq_bits_vd;
  wire [1:0]   queue_1_deq_bits_loadStoreEEW;
  wire         queue_1_deq_bits_mask;
  wire [2:0]   queue_1_deq_bits_segment;
  wire [31:0]  queue_1_deq_bits_readFromScalar;
  wire [11:0]  queue_1_deq_bits_csrInterface_vl;
  wire [11:0]  queue_1_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_1_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_1_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_1_deq_bits_csrInterface_vxrm;
  wire         queue_1_deq_bits_csrInterface_vta;
  wire         queue_1_deq_bits_csrInterface_vma;
  wire         queue_2_deq_ready = laneRequestSinkWire_2_ready;
  wire         queue_2_deq_valid;
  wire [2:0]   queue_2_deq_bits_instructionIndex;
  wire         queue_2_deq_bits_decodeResult_orderReduce;
  wire         queue_2_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_2_deq_bits_decodeResult_fpExecutionType;
  wire         queue_2_deq_bits_decodeResult_float;
  wire         queue_2_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_2_deq_bits_decodeResult_topUop;
  wire         queue_2_deq_bits_decodeResult_popCount;
  wire         queue_2_deq_bits_decodeResult_ffo;
  wire         queue_2_deq_bits_decodeResult_average;
  wire         queue_2_deq_bits_decodeResult_reverse;
  wire         queue_2_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_2_deq_bits_decodeResult_scheduler;
  wire         queue_2_deq_bits_decodeResult_sReadVD;
  wire         queue_2_deq_bits_decodeResult_vtype;
  wire         queue_2_deq_bits_decodeResult_sWrite;
  wire         queue_2_deq_bits_decodeResult_crossRead;
  wire         queue_2_deq_bits_decodeResult_crossWrite;
  wire         queue_2_deq_bits_decodeResult_maskUnit;
  wire         queue_2_deq_bits_decodeResult_special;
  wire         queue_2_deq_bits_decodeResult_saturate;
  wire         queue_2_deq_bits_decodeResult_vwmacc;
  wire         queue_2_deq_bits_decodeResult_readOnly;
  wire         queue_2_deq_bits_decodeResult_maskSource;
  wire         queue_2_deq_bits_decodeResult_maskDestination;
  wire         queue_2_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_2_deq_bits_decodeResult_uop;
  wire         queue_2_deq_bits_decodeResult_iota;
  wire         queue_2_deq_bits_decodeResult_mv;
  wire         queue_2_deq_bits_decodeResult_extend;
  wire         queue_2_deq_bits_decodeResult_unOrderWrite;
  wire         queue_2_deq_bits_decodeResult_compress;
  wire         queue_2_deq_bits_decodeResult_gather16;
  wire         queue_2_deq_bits_decodeResult_gather;
  wire         queue_2_deq_bits_decodeResult_slid;
  wire         queue_2_deq_bits_decodeResult_targetRd;
  wire         queue_2_deq_bits_decodeResult_widenReduce;
  wire         queue_2_deq_bits_decodeResult_red;
  wire         queue_2_deq_bits_decodeResult_nr;
  wire         queue_2_deq_bits_decodeResult_itype;
  wire         queue_2_deq_bits_decodeResult_unsigned1;
  wire         queue_2_deq_bits_decodeResult_unsigned0;
  wire         queue_2_deq_bits_decodeResult_other;
  wire         queue_2_deq_bits_decodeResult_multiCycle;
  wire         queue_2_deq_bits_decodeResult_divider;
  wire         queue_2_deq_bits_decodeResult_multiplier;
  wire         queue_2_deq_bits_decodeResult_shift;
  wire         queue_2_deq_bits_decodeResult_adder;
  wire         queue_2_deq_bits_decodeResult_logic;
  wire         queue_2_deq_bits_loadStore;
  wire         queue_2_deq_bits_issueInst;
  wire         queue_2_deq_bits_store;
  wire         queue_2_deq_bits_special;
  wire         queue_2_deq_bits_lsWholeReg;
  wire [4:0]   queue_2_deq_bits_vs1;
  wire [4:0]   queue_2_deq_bits_vs2;
  wire [4:0]   queue_2_deq_bits_vd;
  wire [1:0]   queue_2_deq_bits_loadStoreEEW;
  wire         queue_2_deq_bits_mask;
  wire [2:0]   queue_2_deq_bits_segment;
  wire [31:0]  queue_2_deq_bits_readFromScalar;
  wire [11:0]  queue_2_deq_bits_csrInterface_vl;
  wire [11:0]  queue_2_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_2_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_2_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_2_deq_bits_csrInterface_vxrm;
  wire         queue_2_deq_bits_csrInterface_vta;
  wire         queue_2_deq_bits_csrInterface_vma;
  wire         queue_3_deq_ready = laneRequestSinkWire_3_ready;
  wire         queue_3_deq_valid;
  wire [2:0]   queue_3_deq_bits_instructionIndex;
  wire         queue_3_deq_bits_decodeResult_orderReduce;
  wire         queue_3_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_3_deq_bits_decodeResult_fpExecutionType;
  wire         queue_3_deq_bits_decodeResult_float;
  wire         queue_3_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_3_deq_bits_decodeResult_topUop;
  wire         queue_3_deq_bits_decodeResult_popCount;
  wire         queue_3_deq_bits_decodeResult_ffo;
  wire         queue_3_deq_bits_decodeResult_average;
  wire         queue_3_deq_bits_decodeResult_reverse;
  wire         queue_3_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_3_deq_bits_decodeResult_scheduler;
  wire         queue_3_deq_bits_decodeResult_sReadVD;
  wire         queue_3_deq_bits_decodeResult_vtype;
  wire         queue_3_deq_bits_decodeResult_sWrite;
  wire         queue_3_deq_bits_decodeResult_crossRead;
  wire         queue_3_deq_bits_decodeResult_crossWrite;
  wire         queue_3_deq_bits_decodeResult_maskUnit;
  wire         queue_3_deq_bits_decodeResult_special;
  wire         queue_3_deq_bits_decodeResult_saturate;
  wire         queue_3_deq_bits_decodeResult_vwmacc;
  wire         queue_3_deq_bits_decodeResult_readOnly;
  wire         queue_3_deq_bits_decodeResult_maskSource;
  wire         queue_3_deq_bits_decodeResult_maskDestination;
  wire         queue_3_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_3_deq_bits_decodeResult_uop;
  wire         queue_3_deq_bits_decodeResult_iota;
  wire         queue_3_deq_bits_decodeResult_mv;
  wire         queue_3_deq_bits_decodeResult_extend;
  wire         queue_3_deq_bits_decodeResult_unOrderWrite;
  wire         queue_3_deq_bits_decodeResult_compress;
  wire         queue_3_deq_bits_decodeResult_gather16;
  wire         queue_3_deq_bits_decodeResult_gather;
  wire         queue_3_deq_bits_decodeResult_slid;
  wire         queue_3_deq_bits_decodeResult_targetRd;
  wire         queue_3_deq_bits_decodeResult_widenReduce;
  wire         queue_3_deq_bits_decodeResult_red;
  wire         queue_3_deq_bits_decodeResult_nr;
  wire         queue_3_deq_bits_decodeResult_itype;
  wire         queue_3_deq_bits_decodeResult_unsigned1;
  wire         queue_3_deq_bits_decodeResult_unsigned0;
  wire         queue_3_deq_bits_decodeResult_other;
  wire         queue_3_deq_bits_decodeResult_multiCycle;
  wire         queue_3_deq_bits_decodeResult_divider;
  wire         queue_3_deq_bits_decodeResult_multiplier;
  wire         queue_3_deq_bits_decodeResult_shift;
  wire         queue_3_deq_bits_decodeResult_adder;
  wire         queue_3_deq_bits_decodeResult_logic;
  wire         queue_3_deq_bits_loadStore;
  wire         queue_3_deq_bits_issueInst;
  wire         queue_3_deq_bits_store;
  wire         queue_3_deq_bits_special;
  wire         queue_3_deq_bits_lsWholeReg;
  wire [4:0]   queue_3_deq_bits_vs1;
  wire [4:0]   queue_3_deq_bits_vs2;
  wire [4:0]   queue_3_deq_bits_vd;
  wire [1:0]   queue_3_deq_bits_loadStoreEEW;
  wire         queue_3_deq_bits_mask;
  wire [2:0]   queue_3_deq_bits_segment;
  wire [31:0]  queue_3_deq_bits_readFromScalar;
  wire [11:0]  queue_3_deq_bits_csrInterface_vl;
  wire [11:0]  queue_3_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_3_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_3_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_3_deq_bits_csrInterface_vxrm;
  wire         queue_3_deq_bits_csrInterface_vta;
  wire         queue_3_deq_bits_csrInterface_vma;
  wire         queue_4_deq_ready = laneRequestSinkWire_4_ready;
  wire         queue_4_deq_valid;
  wire [2:0]   queue_4_deq_bits_instructionIndex;
  wire         queue_4_deq_bits_decodeResult_orderReduce;
  wire         queue_4_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_4_deq_bits_decodeResult_fpExecutionType;
  wire         queue_4_deq_bits_decodeResult_float;
  wire         queue_4_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_4_deq_bits_decodeResult_topUop;
  wire         queue_4_deq_bits_decodeResult_popCount;
  wire         queue_4_deq_bits_decodeResult_ffo;
  wire         queue_4_deq_bits_decodeResult_average;
  wire         queue_4_deq_bits_decodeResult_reverse;
  wire         queue_4_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_4_deq_bits_decodeResult_scheduler;
  wire         queue_4_deq_bits_decodeResult_sReadVD;
  wire         queue_4_deq_bits_decodeResult_vtype;
  wire         queue_4_deq_bits_decodeResult_sWrite;
  wire         queue_4_deq_bits_decodeResult_crossRead;
  wire         queue_4_deq_bits_decodeResult_crossWrite;
  wire         queue_4_deq_bits_decodeResult_maskUnit;
  wire         queue_4_deq_bits_decodeResult_special;
  wire         queue_4_deq_bits_decodeResult_saturate;
  wire         queue_4_deq_bits_decodeResult_vwmacc;
  wire         queue_4_deq_bits_decodeResult_readOnly;
  wire         queue_4_deq_bits_decodeResult_maskSource;
  wire         queue_4_deq_bits_decodeResult_maskDestination;
  wire         queue_4_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_4_deq_bits_decodeResult_uop;
  wire         queue_4_deq_bits_decodeResult_iota;
  wire         queue_4_deq_bits_decodeResult_mv;
  wire         queue_4_deq_bits_decodeResult_extend;
  wire         queue_4_deq_bits_decodeResult_unOrderWrite;
  wire         queue_4_deq_bits_decodeResult_compress;
  wire         queue_4_deq_bits_decodeResult_gather16;
  wire         queue_4_deq_bits_decodeResult_gather;
  wire         queue_4_deq_bits_decodeResult_slid;
  wire         queue_4_deq_bits_decodeResult_targetRd;
  wire         queue_4_deq_bits_decodeResult_widenReduce;
  wire         queue_4_deq_bits_decodeResult_red;
  wire         queue_4_deq_bits_decodeResult_nr;
  wire         queue_4_deq_bits_decodeResult_itype;
  wire         queue_4_deq_bits_decodeResult_unsigned1;
  wire         queue_4_deq_bits_decodeResult_unsigned0;
  wire         queue_4_deq_bits_decodeResult_other;
  wire         queue_4_deq_bits_decodeResult_multiCycle;
  wire         queue_4_deq_bits_decodeResult_divider;
  wire         queue_4_deq_bits_decodeResult_multiplier;
  wire         queue_4_deq_bits_decodeResult_shift;
  wire         queue_4_deq_bits_decodeResult_adder;
  wire         queue_4_deq_bits_decodeResult_logic;
  wire         queue_4_deq_bits_loadStore;
  wire         queue_4_deq_bits_issueInst;
  wire         queue_4_deq_bits_store;
  wire         queue_4_deq_bits_special;
  wire         queue_4_deq_bits_lsWholeReg;
  wire [4:0]   queue_4_deq_bits_vs1;
  wire [4:0]   queue_4_deq_bits_vs2;
  wire [4:0]   queue_4_deq_bits_vd;
  wire [1:0]   queue_4_deq_bits_loadStoreEEW;
  wire         queue_4_deq_bits_mask;
  wire [2:0]   queue_4_deq_bits_segment;
  wire [31:0]  queue_4_deq_bits_readFromScalar;
  wire [11:0]  queue_4_deq_bits_csrInterface_vl;
  wire [11:0]  queue_4_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_4_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_4_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_4_deq_bits_csrInterface_vxrm;
  wire         queue_4_deq_bits_csrInterface_vta;
  wire         queue_4_deq_bits_csrInterface_vma;
  wire         queue_5_deq_ready = laneRequestSinkWire_5_ready;
  wire         queue_5_deq_valid;
  wire [2:0]   queue_5_deq_bits_instructionIndex;
  wire         queue_5_deq_bits_decodeResult_orderReduce;
  wire         queue_5_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_5_deq_bits_decodeResult_fpExecutionType;
  wire         queue_5_deq_bits_decodeResult_float;
  wire         queue_5_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_5_deq_bits_decodeResult_topUop;
  wire         queue_5_deq_bits_decodeResult_popCount;
  wire         queue_5_deq_bits_decodeResult_ffo;
  wire         queue_5_deq_bits_decodeResult_average;
  wire         queue_5_deq_bits_decodeResult_reverse;
  wire         queue_5_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_5_deq_bits_decodeResult_scheduler;
  wire         queue_5_deq_bits_decodeResult_sReadVD;
  wire         queue_5_deq_bits_decodeResult_vtype;
  wire         queue_5_deq_bits_decodeResult_sWrite;
  wire         queue_5_deq_bits_decodeResult_crossRead;
  wire         queue_5_deq_bits_decodeResult_crossWrite;
  wire         queue_5_deq_bits_decodeResult_maskUnit;
  wire         queue_5_deq_bits_decodeResult_special;
  wire         queue_5_deq_bits_decodeResult_saturate;
  wire         queue_5_deq_bits_decodeResult_vwmacc;
  wire         queue_5_deq_bits_decodeResult_readOnly;
  wire         queue_5_deq_bits_decodeResult_maskSource;
  wire         queue_5_deq_bits_decodeResult_maskDestination;
  wire         queue_5_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_5_deq_bits_decodeResult_uop;
  wire         queue_5_deq_bits_decodeResult_iota;
  wire         queue_5_deq_bits_decodeResult_mv;
  wire         queue_5_deq_bits_decodeResult_extend;
  wire         queue_5_deq_bits_decodeResult_unOrderWrite;
  wire         queue_5_deq_bits_decodeResult_compress;
  wire         queue_5_deq_bits_decodeResult_gather16;
  wire         queue_5_deq_bits_decodeResult_gather;
  wire         queue_5_deq_bits_decodeResult_slid;
  wire         queue_5_deq_bits_decodeResult_targetRd;
  wire         queue_5_deq_bits_decodeResult_widenReduce;
  wire         queue_5_deq_bits_decodeResult_red;
  wire         queue_5_deq_bits_decodeResult_nr;
  wire         queue_5_deq_bits_decodeResult_itype;
  wire         queue_5_deq_bits_decodeResult_unsigned1;
  wire         queue_5_deq_bits_decodeResult_unsigned0;
  wire         queue_5_deq_bits_decodeResult_other;
  wire         queue_5_deq_bits_decodeResult_multiCycle;
  wire         queue_5_deq_bits_decodeResult_divider;
  wire         queue_5_deq_bits_decodeResult_multiplier;
  wire         queue_5_deq_bits_decodeResult_shift;
  wire         queue_5_deq_bits_decodeResult_adder;
  wire         queue_5_deq_bits_decodeResult_logic;
  wire         queue_5_deq_bits_loadStore;
  wire         queue_5_deq_bits_issueInst;
  wire         queue_5_deq_bits_store;
  wire         queue_5_deq_bits_special;
  wire         queue_5_deq_bits_lsWholeReg;
  wire [4:0]   queue_5_deq_bits_vs1;
  wire [4:0]   queue_5_deq_bits_vs2;
  wire [4:0]   queue_5_deq_bits_vd;
  wire [1:0]   queue_5_deq_bits_loadStoreEEW;
  wire         queue_5_deq_bits_mask;
  wire [2:0]   queue_5_deq_bits_segment;
  wire [31:0]  queue_5_deq_bits_readFromScalar;
  wire [11:0]  queue_5_deq_bits_csrInterface_vl;
  wire [11:0]  queue_5_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_5_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_5_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_5_deq_bits_csrInterface_vxrm;
  wire         queue_5_deq_bits_csrInterface_vta;
  wire         queue_5_deq_bits_csrInterface_vma;
  wire         queue_6_deq_ready = laneRequestSinkWire_6_ready;
  wire         queue_6_deq_valid;
  wire [2:0]   queue_6_deq_bits_instructionIndex;
  wire         queue_6_deq_bits_decodeResult_orderReduce;
  wire         queue_6_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_6_deq_bits_decodeResult_fpExecutionType;
  wire         queue_6_deq_bits_decodeResult_float;
  wire         queue_6_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_6_deq_bits_decodeResult_topUop;
  wire         queue_6_deq_bits_decodeResult_popCount;
  wire         queue_6_deq_bits_decodeResult_ffo;
  wire         queue_6_deq_bits_decodeResult_average;
  wire         queue_6_deq_bits_decodeResult_reverse;
  wire         queue_6_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_6_deq_bits_decodeResult_scheduler;
  wire         queue_6_deq_bits_decodeResult_sReadVD;
  wire         queue_6_deq_bits_decodeResult_vtype;
  wire         queue_6_deq_bits_decodeResult_sWrite;
  wire         queue_6_deq_bits_decodeResult_crossRead;
  wire         queue_6_deq_bits_decodeResult_crossWrite;
  wire         queue_6_deq_bits_decodeResult_maskUnit;
  wire         queue_6_deq_bits_decodeResult_special;
  wire         queue_6_deq_bits_decodeResult_saturate;
  wire         queue_6_deq_bits_decodeResult_vwmacc;
  wire         queue_6_deq_bits_decodeResult_readOnly;
  wire         queue_6_deq_bits_decodeResult_maskSource;
  wire         queue_6_deq_bits_decodeResult_maskDestination;
  wire         queue_6_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_6_deq_bits_decodeResult_uop;
  wire         queue_6_deq_bits_decodeResult_iota;
  wire         queue_6_deq_bits_decodeResult_mv;
  wire         queue_6_deq_bits_decodeResult_extend;
  wire         queue_6_deq_bits_decodeResult_unOrderWrite;
  wire         queue_6_deq_bits_decodeResult_compress;
  wire         queue_6_deq_bits_decodeResult_gather16;
  wire         queue_6_deq_bits_decodeResult_gather;
  wire         queue_6_deq_bits_decodeResult_slid;
  wire         queue_6_deq_bits_decodeResult_targetRd;
  wire         queue_6_deq_bits_decodeResult_widenReduce;
  wire         queue_6_deq_bits_decodeResult_red;
  wire         queue_6_deq_bits_decodeResult_nr;
  wire         queue_6_deq_bits_decodeResult_itype;
  wire         queue_6_deq_bits_decodeResult_unsigned1;
  wire         queue_6_deq_bits_decodeResult_unsigned0;
  wire         queue_6_deq_bits_decodeResult_other;
  wire         queue_6_deq_bits_decodeResult_multiCycle;
  wire         queue_6_deq_bits_decodeResult_divider;
  wire         queue_6_deq_bits_decodeResult_multiplier;
  wire         queue_6_deq_bits_decodeResult_shift;
  wire         queue_6_deq_bits_decodeResult_adder;
  wire         queue_6_deq_bits_decodeResult_logic;
  wire         queue_6_deq_bits_loadStore;
  wire         queue_6_deq_bits_issueInst;
  wire         queue_6_deq_bits_store;
  wire         queue_6_deq_bits_special;
  wire         queue_6_deq_bits_lsWholeReg;
  wire [4:0]   queue_6_deq_bits_vs1;
  wire [4:0]   queue_6_deq_bits_vs2;
  wire [4:0]   queue_6_deq_bits_vd;
  wire [1:0]   queue_6_deq_bits_loadStoreEEW;
  wire         queue_6_deq_bits_mask;
  wire [2:0]   queue_6_deq_bits_segment;
  wire [31:0]  queue_6_deq_bits_readFromScalar;
  wire [11:0]  queue_6_deq_bits_csrInterface_vl;
  wire [11:0]  queue_6_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_6_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_6_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_6_deq_bits_csrInterface_vxrm;
  wire         queue_6_deq_bits_csrInterface_vta;
  wire         queue_6_deq_bits_csrInterface_vma;
  wire         queue_7_deq_ready = laneRequestSinkWire_7_ready;
  wire         queue_7_deq_valid;
  wire [2:0]   queue_7_deq_bits_instructionIndex;
  wire         queue_7_deq_bits_decodeResult_orderReduce;
  wire         queue_7_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_7_deq_bits_decodeResult_fpExecutionType;
  wire         queue_7_deq_bits_decodeResult_float;
  wire         queue_7_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_7_deq_bits_decodeResult_topUop;
  wire         queue_7_deq_bits_decodeResult_popCount;
  wire         queue_7_deq_bits_decodeResult_ffo;
  wire         queue_7_deq_bits_decodeResult_average;
  wire         queue_7_deq_bits_decodeResult_reverse;
  wire         queue_7_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_7_deq_bits_decodeResult_scheduler;
  wire         queue_7_deq_bits_decodeResult_sReadVD;
  wire         queue_7_deq_bits_decodeResult_vtype;
  wire         queue_7_deq_bits_decodeResult_sWrite;
  wire         queue_7_deq_bits_decodeResult_crossRead;
  wire         queue_7_deq_bits_decodeResult_crossWrite;
  wire         queue_7_deq_bits_decodeResult_maskUnit;
  wire         queue_7_deq_bits_decodeResult_special;
  wire         queue_7_deq_bits_decodeResult_saturate;
  wire         queue_7_deq_bits_decodeResult_vwmacc;
  wire         queue_7_deq_bits_decodeResult_readOnly;
  wire         queue_7_deq_bits_decodeResult_maskSource;
  wire         queue_7_deq_bits_decodeResult_maskDestination;
  wire         queue_7_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_7_deq_bits_decodeResult_uop;
  wire         queue_7_deq_bits_decodeResult_iota;
  wire         queue_7_deq_bits_decodeResult_mv;
  wire         queue_7_deq_bits_decodeResult_extend;
  wire         queue_7_deq_bits_decodeResult_unOrderWrite;
  wire         queue_7_deq_bits_decodeResult_compress;
  wire         queue_7_deq_bits_decodeResult_gather16;
  wire         queue_7_deq_bits_decodeResult_gather;
  wire         queue_7_deq_bits_decodeResult_slid;
  wire         queue_7_deq_bits_decodeResult_targetRd;
  wire         queue_7_deq_bits_decodeResult_widenReduce;
  wire         queue_7_deq_bits_decodeResult_red;
  wire         queue_7_deq_bits_decodeResult_nr;
  wire         queue_7_deq_bits_decodeResult_itype;
  wire         queue_7_deq_bits_decodeResult_unsigned1;
  wire         queue_7_deq_bits_decodeResult_unsigned0;
  wire         queue_7_deq_bits_decodeResult_other;
  wire         queue_7_deq_bits_decodeResult_multiCycle;
  wire         queue_7_deq_bits_decodeResult_divider;
  wire         queue_7_deq_bits_decodeResult_multiplier;
  wire         queue_7_deq_bits_decodeResult_shift;
  wire         queue_7_deq_bits_decodeResult_adder;
  wire         queue_7_deq_bits_decodeResult_logic;
  wire         queue_7_deq_bits_loadStore;
  wire         queue_7_deq_bits_issueInst;
  wire         queue_7_deq_bits_store;
  wire         queue_7_deq_bits_special;
  wire         queue_7_deq_bits_lsWholeReg;
  wire [4:0]   queue_7_deq_bits_vs1;
  wire [4:0]   queue_7_deq_bits_vs2;
  wire [4:0]   queue_7_deq_bits_vd;
  wire [1:0]   queue_7_deq_bits_loadStoreEEW;
  wire         queue_7_deq_bits_mask;
  wire [2:0]   queue_7_deq_bits_segment;
  wire [31:0]  queue_7_deq_bits_readFromScalar;
  wire [11:0]  queue_7_deq_bits_csrInterface_vl;
  wire [11:0]  queue_7_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_7_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_7_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_7_deq_bits_csrInterface_vxrm;
  wire         queue_7_deq_bits_csrInterface_vta;
  wire         queue_7_deq_bits_csrInterface_vma;
  wire         queue_8_deq_ready = laneRequestSinkWire_8_ready;
  wire         queue_8_deq_valid;
  wire [2:0]   queue_8_deq_bits_instructionIndex;
  wire         queue_8_deq_bits_decodeResult_orderReduce;
  wire         queue_8_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_8_deq_bits_decodeResult_fpExecutionType;
  wire         queue_8_deq_bits_decodeResult_float;
  wire         queue_8_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_8_deq_bits_decodeResult_topUop;
  wire         queue_8_deq_bits_decodeResult_popCount;
  wire         queue_8_deq_bits_decodeResult_ffo;
  wire         queue_8_deq_bits_decodeResult_average;
  wire         queue_8_deq_bits_decodeResult_reverse;
  wire         queue_8_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_8_deq_bits_decodeResult_scheduler;
  wire         queue_8_deq_bits_decodeResult_sReadVD;
  wire         queue_8_deq_bits_decodeResult_vtype;
  wire         queue_8_deq_bits_decodeResult_sWrite;
  wire         queue_8_deq_bits_decodeResult_crossRead;
  wire         queue_8_deq_bits_decodeResult_crossWrite;
  wire         queue_8_deq_bits_decodeResult_maskUnit;
  wire         queue_8_deq_bits_decodeResult_special;
  wire         queue_8_deq_bits_decodeResult_saturate;
  wire         queue_8_deq_bits_decodeResult_vwmacc;
  wire         queue_8_deq_bits_decodeResult_readOnly;
  wire         queue_8_deq_bits_decodeResult_maskSource;
  wire         queue_8_deq_bits_decodeResult_maskDestination;
  wire         queue_8_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_8_deq_bits_decodeResult_uop;
  wire         queue_8_deq_bits_decodeResult_iota;
  wire         queue_8_deq_bits_decodeResult_mv;
  wire         queue_8_deq_bits_decodeResult_extend;
  wire         queue_8_deq_bits_decodeResult_unOrderWrite;
  wire         queue_8_deq_bits_decodeResult_compress;
  wire         queue_8_deq_bits_decodeResult_gather16;
  wire         queue_8_deq_bits_decodeResult_gather;
  wire         queue_8_deq_bits_decodeResult_slid;
  wire         queue_8_deq_bits_decodeResult_targetRd;
  wire         queue_8_deq_bits_decodeResult_widenReduce;
  wire         queue_8_deq_bits_decodeResult_red;
  wire         queue_8_deq_bits_decodeResult_nr;
  wire         queue_8_deq_bits_decodeResult_itype;
  wire         queue_8_deq_bits_decodeResult_unsigned1;
  wire         queue_8_deq_bits_decodeResult_unsigned0;
  wire         queue_8_deq_bits_decodeResult_other;
  wire         queue_8_deq_bits_decodeResult_multiCycle;
  wire         queue_8_deq_bits_decodeResult_divider;
  wire         queue_8_deq_bits_decodeResult_multiplier;
  wire         queue_8_deq_bits_decodeResult_shift;
  wire         queue_8_deq_bits_decodeResult_adder;
  wire         queue_8_deq_bits_decodeResult_logic;
  wire         queue_8_deq_bits_loadStore;
  wire         queue_8_deq_bits_issueInst;
  wire         queue_8_deq_bits_store;
  wire         queue_8_deq_bits_special;
  wire         queue_8_deq_bits_lsWholeReg;
  wire [4:0]   queue_8_deq_bits_vs1;
  wire [4:0]   queue_8_deq_bits_vs2;
  wire [4:0]   queue_8_deq_bits_vd;
  wire [1:0]   queue_8_deq_bits_loadStoreEEW;
  wire         queue_8_deq_bits_mask;
  wire [2:0]   queue_8_deq_bits_segment;
  wire [31:0]  queue_8_deq_bits_readFromScalar;
  wire [11:0]  queue_8_deq_bits_csrInterface_vl;
  wire [11:0]  queue_8_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_8_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_8_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_8_deq_bits_csrInterface_vxrm;
  wire         queue_8_deq_bits_csrInterface_vta;
  wire         queue_8_deq_bits_csrInterface_vma;
  wire         queue_9_deq_ready = laneRequestSinkWire_9_ready;
  wire         queue_9_deq_valid;
  wire [2:0]   queue_9_deq_bits_instructionIndex;
  wire         queue_9_deq_bits_decodeResult_orderReduce;
  wire         queue_9_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_9_deq_bits_decodeResult_fpExecutionType;
  wire         queue_9_deq_bits_decodeResult_float;
  wire         queue_9_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_9_deq_bits_decodeResult_topUop;
  wire         queue_9_deq_bits_decodeResult_popCount;
  wire         queue_9_deq_bits_decodeResult_ffo;
  wire         queue_9_deq_bits_decodeResult_average;
  wire         queue_9_deq_bits_decodeResult_reverse;
  wire         queue_9_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_9_deq_bits_decodeResult_scheduler;
  wire         queue_9_deq_bits_decodeResult_sReadVD;
  wire         queue_9_deq_bits_decodeResult_vtype;
  wire         queue_9_deq_bits_decodeResult_sWrite;
  wire         queue_9_deq_bits_decodeResult_crossRead;
  wire         queue_9_deq_bits_decodeResult_crossWrite;
  wire         queue_9_deq_bits_decodeResult_maskUnit;
  wire         queue_9_deq_bits_decodeResult_special;
  wire         queue_9_deq_bits_decodeResult_saturate;
  wire         queue_9_deq_bits_decodeResult_vwmacc;
  wire         queue_9_deq_bits_decodeResult_readOnly;
  wire         queue_9_deq_bits_decodeResult_maskSource;
  wire         queue_9_deq_bits_decodeResult_maskDestination;
  wire         queue_9_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_9_deq_bits_decodeResult_uop;
  wire         queue_9_deq_bits_decodeResult_iota;
  wire         queue_9_deq_bits_decodeResult_mv;
  wire         queue_9_deq_bits_decodeResult_extend;
  wire         queue_9_deq_bits_decodeResult_unOrderWrite;
  wire         queue_9_deq_bits_decodeResult_compress;
  wire         queue_9_deq_bits_decodeResult_gather16;
  wire         queue_9_deq_bits_decodeResult_gather;
  wire         queue_9_deq_bits_decodeResult_slid;
  wire         queue_9_deq_bits_decodeResult_targetRd;
  wire         queue_9_deq_bits_decodeResult_widenReduce;
  wire         queue_9_deq_bits_decodeResult_red;
  wire         queue_9_deq_bits_decodeResult_nr;
  wire         queue_9_deq_bits_decodeResult_itype;
  wire         queue_9_deq_bits_decodeResult_unsigned1;
  wire         queue_9_deq_bits_decodeResult_unsigned0;
  wire         queue_9_deq_bits_decodeResult_other;
  wire         queue_9_deq_bits_decodeResult_multiCycle;
  wire         queue_9_deq_bits_decodeResult_divider;
  wire         queue_9_deq_bits_decodeResult_multiplier;
  wire         queue_9_deq_bits_decodeResult_shift;
  wire         queue_9_deq_bits_decodeResult_adder;
  wire         queue_9_deq_bits_decodeResult_logic;
  wire         queue_9_deq_bits_loadStore;
  wire         queue_9_deq_bits_issueInst;
  wire         queue_9_deq_bits_store;
  wire         queue_9_deq_bits_special;
  wire         queue_9_deq_bits_lsWholeReg;
  wire [4:0]   queue_9_deq_bits_vs1;
  wire [4:0]   queue_9_deq_bits_vs2;
  wire [4:0]   queue_9_deq_bits_vd;
  wire [1:0]   queue_9_deq_bits_loadStoreEEW;
  wire         queue_9_deq_bits_mask;
  wire [2:0]   queue_9_deq_bits_segment;
  wire [31:0]  queue_9_deq_bits_readFromScalar;
  wire [11:0]  queue_9_deq_bits_csrInterface_vl;
  wire [11:0]  queue_9_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_9_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_9_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_9_deq_bits_csrInterface_vxrm;
  wire         queue_9_deq_bits_csrInterface_vta;
  wire         queue_9_deq_bits_csrInterface_vma;
  wire         queue_10_deq_ready = laneRequestSinkWire_10_ready;
  wire         queue_10_deq_valid;
  wire [2:0]   queue_10_deq_bits_instructionIndex;
  wire         queue_10_deq_bits_decodeResult_orderReduce;
  wire         queue_10_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_10_deq_bits_decodeResult_fpExecutionType;
  wire         queue_10_deq_bits_decodeResult_float;
  wire         queue_10_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_10_deq_bits_decodeResult_topUop;
  wire         queue_10_deq_bits_decodeResult_popCount;
  wire         queue_10_deq_bits_decodeResult_ffo;
  wire         queue_10_deq_bits_decodeResult_average;
  wire         queue_10_deq_bits_decodeResult_reverse;
  wire         queue_10_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_10_deq_bits_decodeResult_scheduler;
  wire         queue_10_deq_bits_decodeResult_sReadVD;
  wire         queue_10_deq_bits_decodeResult_vtype;
  wire         queue_10_deq_bits_decodeResult_sWrite;
  wire         queue_10_deq_bits_decodeResult_crossRead;
  wire         queue_10_deq_bits_decodeResult_crossWrite;
  wire         queue_10_deq_bits_decodeResult_maskUnit;
  wire         queue_10_deq_bits_decodeResult_special;
  wire         queue_10_deq_bits_decodeResult_saturate;
  wire         queue_10_deq_bits_decodeResult_vwmacc;
  wire         queue_10_deq_bits_decodeResult_readOnly;
  wire         queue_10_deq_bits_decodeResult_maskSource;
  wire         queue_10_deq_bits_decodeResult_maskDestination;
  wire         queue_10_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_10_deq_bits_decodeResult_uop;
  wire         queue_10_deq_bits_decodeResult_iota;
  wire         queue_10_deq_bits_decodeResult_mv;
  wire         queue_10_deq_bits_decodeResult_extend;
  wire         queue_10_deq_bits_decodeResult_unOrderWrite;
  wire         queue_10_deq_bits_decodeResult_compress;
  wire         queue_10_deq_bits_decodeResult_gather16;
  wire         queue_10_deq_bits_decodeResult_gather;
  wire         queue_10_deq_bits_decodeResult_slid;
  wire         queue_10_deq_bits_decodeResult_targetRd;
  wire         queue_10_deq_bits_decodeResult_widenReduce;
  wire         queue_10_deq_bits_decodeResult_red;
  wire         queue_10_deq_bits_decodeResult_nr;
  wire         queue_10_deq_bits_decodeResult_itype;
  wire         queue_10_deq_bits_decodeResult_unsigned1;
  wire         queue_10_deq_bits_decodeResult_unsigned0;
  wire         queue_10_deq_bits_decodeResult_other;
  wire         queue_10_deq_bits_decodeResult_multiCycle;
  wire         queue_10_deq_bits_decodeResult_divider;
  wire         queue_10_deq_bits_decodeResult_multiplier;
  wire         queue_10_deq_bits_decodeResult_shift;
  wire         queue_10_deq_bits_decodeResult_adder;
  wire         queue_10_deq_bits_decodeResult_logic;
  wire         queue_10_deq_bits_loadStore;
  wire         queue_10_deq_bits_issueInst;
  wire         queue_10_deq_bits_store;
  wire         queue_10_deq_bits_special;
  wire         queue_10_deq_bits_lsWholeReg;
  wire [4:0]   queue_10_deq_bits_vs1;
  wire [4:0]   queue_10_deq_bits_vs2;
  wire [4:0]   queue_10_deq_bits_vd;
  wire [1:0]   queue_10_deq_bits_loadStoreEEW;
  wire         queue_10_deq_bits_mask;
  wire [2:0]   queue_10_deq_bits_segment;
  wire [31:0]  queue_10_deq_bits_readFromScalar;
  wire [11:0]  queue_10_deq_bits_csrInterface_vl;
  wire [11:0]  queue_10_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_10_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_10_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_10_deq_bits_csrInterface_vxrm;
  wire         queue_10_deq_bits_csrInterface_vta;
  wire         queue_10_deq_bits_csrInterface_vma;
  wire         queue_11_deq_ready = laneRequestSinkWire_11_ready;
  wire         queue_11_deq_valid;
  wire [2:0]   queue_11_deq_bits_instructionIndex;
  wire         queue_11_deq_bits_decodeResult_orderReduce;
  wire         queue_11_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_11_deq_bits_decodeResult_fpExecutionType;
  wire         queue_11_deq_bits_decodeResult_float;
  wire         queue_11_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_11_deq_bits_decodeResult_topUop;
  wire         queue_11_deq_bits_decodeResult_popCount;
  wire         queue_11_deq_bits_decodeResult_ffo;
  wire         queue_11_deq_bits_decodeResult_average;
  wire         queue_11_deq_bits_decodeResult_reverse;
  wire         queue_11_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_11_deq_bits_decodeResult_scheduler;
  wire         queue_11_deq_bits_decodeResult_sReadVD;
  wire         queue_11_deq_bits_decodeResult_vtype;
  wire         queue_11_deq_bits_decodeResult_sWrite;
  wire         queue_11_deq_bits_decodeResult_crossRead;
  wire         queue_11_deq_bits_decodeResult_crossWrite;
  wire         queue_11_deq_bits_decodeResult_maskUnit;
  wire         queue_11_deq_bits_decodeResult_special;
  wire         queue_11_deq_bits_decodeResult_saturate;
  wire         queue_11_deq_bits_decodeResult_vwmacc;
  wire         queue_11_deq_bits_decodeResult_readOnly;
  wire         queue_11_deq_bits_decodeResult_maskSource;
  wire         queue_11_deq_bits_decodeResult_maskDestination;
  wire         queue_11_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_11_deq_bits_decodeResult_uop;
  wire         queue_11_deq_bits_decodeResult_iota;
  wire         queue_11_deq_bits_decodeResult_mv;
  wire         queue_11_deq_bits_decodeResult_extend;
  wire         queue_11_deq_bits_decodeResult_unOrderWrite;
  wire         queue_11_deq_bits_decodeResult_compress;
  wire         queue_11_deq_bits_decodeResult_gather16;
  wire         queue_11_deq_bits_decodeResult_gather;
  wire         queue_11_deq_bits_decodeResult_slid;
  wire         queue_11_deq_bits_decodeResult_targetRd;
  wire         queue_11_deq_bits_decodeResult_widenReduce;
  wire         queue_11_deq_bits_decodeResult_red;
  wire         queue_11_deq_bits_decodeResult_nr;
  wire         queue_11_deq_bits_decodeResult_itype;
  wire         queue_11_deq_bits_decodeResult_unsigned1;
  wire         queue_11_deq_bits_decodeResult_unsigned0;
  wire         queue_11_deq_bits_decodeResult_other;
  wire         queue_11_deq_bits_decodeResult_multiCycle;
  wire         queue_11_deq_bits_decodeResult_divider;
  wire         queue_11_deq_bits_decodeResult_multiplier;
  wire         queue_11_deq_bits_decodeResult_shift;
  wire         queue_11_deq_bits_decodeResult_adder;
  wire         queue_11_deq_bits_decodeResult_logic;
  wire         queue_11_deq_bits_loadStore;
  wire         queue_11_deq_bits_issueInst;
  wire         queue_11_deq_bits_store;
  wire         queue_11_deq_bits_special;
  wire         queue_11_deq_bits_lsWholeReg;
  wire [4:0]   queue_11_deq_bits_vs1;
  wire [4:0]   queue_11_deq_bits_vs2;
  wire [4:0]   queue_11_deq_bits_vd;
  wire [1:0]   queue_11_deq_bits_loadStoreEEW;
  wire         queue_11_deq_bits_mask;
  wire [2:0]   queue_11_deq_bits_segment;
  wire [31:0]  queue_11_deq_bits_readFromScalar;
  wire [11:0]  queue_11_deq_bits_csrInterface_vl;
  wire [11:0]  queue_11_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_11_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_11_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_11_deq_bits_csrInterface_vxrm;
  wire         queue_11_deq_bits_csrInterface_vta;
  wire         queue_11_deq_bits_csrInterface_vma;
  wire         queue_12_deq_ready = laneRequestSinkWire_12_ready;
  wire         queue_12_deq_valid;
  wire [2:0]   queue_12_deq_bits_instructionIndex;
  wire         queue_12_deq_bits_decodeResult_orderReduce;
  wire         queue_12_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_12_deq_bits_decodeResult_fpExecutionType;
  wire         queue_12_deq_bits_decodeResult_float;
  wire         queue_12_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_12_deq_bits_decodeResult_topUop;
  wire         queue_12_deq_bits_decodeResult_popCount;
  wire         queue_12_deq_bits_decodeResult_ffo;
  wire         queue_12_deq_bits_decodeResult_average;
  wire         queue_12_deq_bits_decodeResult_reverse;
  wire         queue_12_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_12_deq_bits_decodeResult_scheduler;
  wire         queue_12_deq_bits_decodeResult_sReadVD;
  wire         queue_12_deq_bits_decodeResult_vtype;
  wire         queue_12_deq_bits_decodeResult_sWrite;
  wire         queue_12_deq_bits_decodeResult_crossRead;
  wire         queue_12_deq_bits_decodeResult_crossWrite;
  wire         queue_12_deq_bits_decodeResult_maskUnit;
  wire         queue_12_deq_bits_decodeResult_special;
  wire         queue_12_deq_bits_decodeResult_saturate;
  wire         queue_12_deq_bits_decodeResult_vwmacc;
  wire         queue_12_deq_bits_decodeResult_readOnly;
  wire         queue_12_deq_bits_decodeResult_maskSource;
  wire         queue_12_deq_bits_decodeResult_maskDestination;
  wire         queue_12_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_12_deq_bits_decodeResult_uop;
  wire         queue_12_deq_bits_decodeResult_iota;
  wire         queue_12_deq_bits_decodeResult_mv;
  wire         queue_12_deq_bits_decodeResult_extend;
  wire         queue_12_deq_bits_decodeResult_unOrderWrite;
  wire         queue_12_deq_bits_decodeResult_compress;
  wire         queue_12_deq_bits_decodeResult_gather16;
  wire         queue_12_deq_bits_decodeResult_gather;
  wire         queue_12_deq_bits_decodeResult_slid;
  wire         queue_12_deq_bits_decodeResult_targetRd;
  wire         queue_12_deq_bits_decodeResult_widenReduce;
  wire         queue_12_deq_bits_decodeResult_red;
  wire         queue_12_deq_bits_decodeResult_nr;
  wire         queue_12_deq_bits_decodeResult_itype;
  wire         queue_12_deq_bits_decodeResult_unsigned1;
  wire         queue_12_deq_bits_decodeResult_unsigned0;
  wire         queue_12_deq_bits_decodeResult_other;
  wire         queue_12_deq_bits_decodeResult_multiCycle;
  wire         queue_12_deq_bits_decodeResult_divider;
  wire         queue_12_deq_bits_decodeResult_multiplier;
  wire         queue_12_deq_bits_decodeResult_shift;
  wire         queue_12_deq_bits_decodeResult_adder;
  wire         queue_12_deq_bits_decodeResult_logic;
  wire         queue_12_deq_bits_loadStore;
  wire         queue_12_deq_bits_issueInst;
  wire         queue_12_deq_bits_store;
  wire         queue_12_deq_bits_special;
  wire         queue_12_deq_bits_lsWholeReg;
  wire [4:0]   queue_12_deq_bits_vs1;
  wire [4:0]   queue_12_deq_bits_vs2;
  wire [4:0]   queue_12_deq_bits_vd;
  wire [1:0]   queue_12_deq_bits_loadStoreEEW;
  wire         queue_12_deq_bits_mask;
  wire [2:0]   queue_12_deq_bits_segment;
  wire [31:0]  queue_12_deq_bits_readFromScalar;
  wire [11:0]  queue_12_deq_bits_csrInterface_vl;
  wire [11:0]  queue_12_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_12_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_12_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_12_deq_bits_csrInterface_vxrm;
  wire         queue_12_deq_bits_csrInterface_vta;
  wire         queue_12_deq_bits_csrInterface_vma;
  wire         queue_13_deq_ready = laneRequestSinkWire_13_ready;
  wire         queue_13_deq_valid;
  wire [2:0]   queue_13_deq_bits_instructionIndex;
  wire         queue_13_deq_bits_decodeResult_orderReduce;
  wire         queue_13_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_13_deq_bits_decodeResult_fpExecutionType;
  wire         queue_13_deq_bits_decodeResult_float;
  wire         queue_13_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_13_deq_bits_decodeResult_topUop;
  wire         queue_13_deq_bits_decodeResult_popCount;
  wire         queue_13_deq_bits_decodeResult_ffo;
  wire         queue_13_deq_bits_decodeResult_average;
  wire         queue_13_deq_bits_decodeResult_reverse;
  wire         queue_13_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_13_deq_bits_decodeResult_scheduler;
  wire         queue_13_deq_bits_decodeResult_sReadVD;
  wire         queue_13_deq_bits_decodeResult_vtype;
  wire         queue_13_deq_bits_decodeResult_sWrite;
  wire         queue_13_deq_bits_decodeResult_crossRead;
  wire         queue_13_deq_bits_decodeResult_crossWrite;
  wire         queue_13_deq_bits_decodeResult_maskUnit;
  wire         queue_13_deq_bits_decodeResult_special;
  wire         queue_13_deq_bits_decodeResult_saturate;
  wire         queue_13_deq_bits_decodeResult_vwmacc;
  wire         queue_13_deq_bits_decodeResult_readOnly;
  wire         queue_13_deq_bits_decodeResult_maskSource;
  wire         queue_13_deq_bits_decodeResult_maskDestination;
  wire         queue_13_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_13_deq_bits_decodeResult_uop;
  wire         queue_13_deq_bits_decodeResult_iota;
  wire         queue_13_deq_bits_decodeResult_mv;
  wire         queue_13_deq_bits_decodeResult_extend;
  wire         queue_13_deq_bits_decodeResult_unOrderWrite;
  wire         queue_13_deq_bits_decodeResult_compress;
  wire         queue_13_deq_bits_decodeResult_gather16;
  wire         queue_13_deq_bits_decodeResult_gather;
  wire         queue_13_deq_bits_decodeResult_slid;
  wire         queue_13_deq_bits_decodeResult_targetRd;
  wire         queue_13_deq_bits_decodeResult_widenReduce;
  wire         queue_13_deq_bits_decodeResult_red;
  wire         queue_13_deq_bits_decodeResult_nr;
  wire         queue_13_deq_bits_decodeResult_itype;
  wire         queue_13_deq_bits_decodeResult_unsigned1;
  wire         queue_13_deq_bits_decodeResult_unsigned0;
  wire         queue_13_deq_bits_decodeResult_other;
  wire         queue_13_deq_bits_decodeResult_multiCycle;
  wire         queue_13_deq_bits_decodeResult_divider;
  wire         queue_13_deq_bits_decodeResult_multiplier;
  wire         queue_13_deq_bits_decodeResult_shift;
  wire         queue_13_deq_bits_decodeResult_adder;
  wire         queue_13_deq_bits_decodeResult_logic;
  wire         queue_13_deq_bits_loadStore;
  wire         queue_13_deq_bits_issueInst;
  wire         queue_13_deq_bits_store;
  wire         queue_13_deq_bits_special;
  wire         queue_13_deq_bits_lsWholeReg;
  wire [4:0]   queue_13_deq_bits_vs1;
  wire [4:0]   queue_13_deq_bits_vs2;
  wire [4:0]   queue_13_deq_bits_vd;
  wire [1:0]   queue_13_deq_bits_loadStoreEEW;
  wire         queue_13_deq_bits_mask;
  wire [2:0]   queue_13_deq_bits_segment;
  wire [31:0]  queue_13_deq_bits_readFromScalar;
  wire [11:0]  queue_13_deq_bits_csrInterface_vl;
  wire [11:0]  queue_13_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_13_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_13_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_13_deq_bits_csrInterface_vxrm;
  wire         queue_13_deq_bits_csrInterface_vta;
  wire         queue_13_deq_bits_csrInterface_vma;
  wire         queue_14_deq_ready = laneRequestSinkWire_14_ready;
  wire         queue_14_deq_valid;
  wire [2:0]   queue_14_deq_bits_instructionIndex;
  wire         queue_14_deq_bits_decodeResult_orderReduce;
  wire         queue_14_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_14_deq_bits_decodeResult_fpExecutionType;
  wire         queue_14_deq_bits_decodeResult_float;
  wire         queue_14_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_14_deq_bits_decodeResult_topUop;
  wire         queue_14_deq_bits_decodeResult_popCount;
  wire         queue_14_deq_bits_decodeResult_ffo;
  wire         queue_14_deq_bits_decodeResult_average;
  wire         queue_14_deq_bits_decodeResult_reverse;
  wire         queue_14_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_14_deq_bits_decodeResult_scheduler;
  wire         queue_14_deq_bits_decodeResult_sReadVD;
  wire         queue_14_deq_bits_decodeResult_vtype;
  wire         queue_14_deq_bits_decodeResult_sWrite;
  wire         queue_14_deq_bits_decodeResult_crossRead;
  wire         queue_14_deq_bits_decodeResult_crossWrite;
  wire         queue_14_deq_bits_decodeResult_maskUnit;
  wire         queue_14_deq_bits_decodeResult_special;
  wire         queue_14_deq_bits_decodeResult_saturate;
  wire         queue_14_deq_bits_decodeResult_vwmacc;
  wire         queue_14_deq_bits_decodeResult_readOnly;
  wire         queue_14_deq_bits_decodeResult_maskSource;
  wire         queue_14_deq_bits_decodeResult_maskDestination;
  wire         queue_14_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_14_deq_bits_decodeResult_uop;
  wire         queue_14_deq_bits_decodeResult_iota;
  wire         queue_14_deq_bits_decodeResult_mv;
  wire         queue_14_deq_bits_decodeResult_extend;
  wire         queue_14_deq_bits_decodeResult_unOrderWrite;
  wire         queue_14_deq_bits_decodeResult_compress;
  wire         queue_14_deq_bits_decodeResult_gather16;
  wire         queue_14_deq_bits_decodeResult_gather;
  wire         queue_14_deq_bits_decodeResult_slid;
  wire         queue_14_deq_bits_decodeResult_targetRd;
  wire         queue_14_deq_bits_decodeResult_widenReduce;
  wire         queue_14_deq_bits_decodeResult_red;
  wire         queue_14_deq_bits_decodeResult_nr;
  wire         queue_14_deq_bits_decodeResult_itype;
  wire         queue_14_deq_bits_decodeResult_unsigned1;
  wire         queue_14_deq_bits_decodeResult_unsigned0;
  wire         queue_14_deq_bits_decodeResult_other;
  wire         queue_14_deq_bits_decodeResult_multiCycle;
  wire         queue_14_deq_bits_decodeResult_divider;
  wire         queue_14_deq_bits_decodeResult_multiplier;
  wire         queue_14_deq_bits_decodeResult_shift;
  wire         queue_14_deq_bits_decodeResult_adder;
  wire         queue_14_deq_bits_decodeResult_logic;
  wire         queue_14_deq_bits_loadStore;
  wire         queue_14_deq_bits_issueInst;
  wire         queue_14_deq_bits_store;
  wire         queue_14_deq_bits_special;
  wire         queue_14_deq_bits_lsWholeReg;
  wire [4:0]   queue_14_deq_bits_vs1;
  wire [4:0]   queue_14_deq_bits_vs2;
  wire [4:0]   queue_14_deq_bits_vd;
  wire [1:0]   queue_14_deq_bits_loadStoreEEW;
  wire         queue_14_deq_bits_mask;
  wire [2:0]   queue_14_deq_bits_segment;
  wire [31:0]  queue_14_deq_bits_readFromScalar;
  wire [11:0]  queue_14_deq_bits_csrInterface_vl;
  wire [11:0]  queue_14_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_14_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_14_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_14_deq_bits_csrInterface_vxrm;
  wire         queue_14_deq_bits_csrInterface_vta;
  wire         queue_14_deq_bits_csrInterface_vma;
  wire         queue_15_deq_ready = laneRequestSinkWire_15_ready;
  wire         queue_15_deq_valid;
  wire [2:0]   queue_15_deq_bits_instructionIndex;
  wire         queue_15_deq_bits_decodeResult_orderReduce;
  wire         queue_15_deq_bits_decodeResult_floatMul;
  wire [1:0]   queue_15_deq_bits_decodeResult_fpExecutionType;
  wire         queue_15_deq_bits_decodeResult_float;
  wire         queue_15_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_15_deq_bits_decodeResult_topUop;
  wire         queue_15_deq_bits_decodeResult_popCount;
  wire         queue_15_deq_bits_decodeResult_ffo;
  wire         queue_15_deq_bits_decodeResult_average;
  wire         queue_15_deq_bits_decodeResult_reverse;
  wire         queue_15_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_15_deq_bits_decodeResult_scheduler;
  wire         queue_15_deq_bits_decodeResult_sReadVD;
  wire         queue_15_deq_bits_decodeResult_vtype;
  wire         queue_15_deq_bits_decodeResult_sWrite;
  wire         queue_15_deq_bits_decodeResult_crossRead;
  wire         queue_15_deq_bits_decodeResult_crossWrite;
  wire         queue_15_deq_bits_decodeResult_maskUnit;
  wire         queue_15_deq_bits_decodeResult_special;
  wire         queue_15_deq_bits_decodeResult_saturate;
  wire         queue_15_deq_bits_decodeResult_vwmacc;
  wire         queue_15_deq_bits_decodeResult_readOnly;
  wire         queue_15_deq_bits_decodeResult_maskSource;
  wire         queue_15_deq_bits_decodeResult_maskDestination;
  wire         queue_15_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_15_deq_bits_decodeResult_uop;
  wire         queue_15_deq_bits_decodeResult_iota;
  wire         queue_15_deq_bits_decodeResult_mv;
  wire         queue_15_deq_bits_decodeResult_extend;
  wire         queue_15_deq_bits_decodeResult_unOrderWrite;
  wire         queue_15_deq_bits_decodeResult_compress;
  wire         queue_15_deq_bits_decodeResult_gather16;
  wire         queue_15_deq_bits_decodeResult_gather;
  wire         queue_15_deq_bits_decodeResult_slid;
  wire         queue_15_deq_bits_decodeResult_targetRd;
  wire         queue_15_deq_bits_decodeResult_widenReduce;
  wire         queue_15_deq_bits_decodeResult_red;
  wire         queue_15_deq_bits_decodeResult_nr;
  wire         queue_15_deq_bits_decodeResult_itype;
  wire         queue_15_deq_bits_decodeResult_unsigned1;
  wire         queue_15_deq_bits_decodeResult_unsigned0;
  wire         queue_15_deq_bits_decodeResult_other;
  wire         queue_15_deq_bits_decodeResult_multiCycle;
  wire         queue_15_deq_bits_decodeResult_divider;
  wire         queue_15_deq_bits_decodeResult_multiplier;
  wire         queue_15_deq_bits_decodeResult_shift;
  wire         queue_15_deq_bits_decodeResult_adder;
  wire         queue_15_deq_bits_decodeResult_logic;
  wire         queue_15_deq_bits_loadStore;
  wire         queue_15_deq_bits_issueInst;
  wire         queue_15_deq_bits_store;
  wire         queue_15_deq_bits_special;
  wire         queue_15_deq_bits_lsWholeReg;
  wire [4:0]   queue_15_deq_bits_vs1;
  wire [4:0]   queue_15_deq_bits_vs2;
  wire [4:0]   queue_15_deq_bits_vd;
  wire [1:0]   queue_15_deq_bits_loadStoreEEW;
  wire         queue_15_deq_bits_mask;
  wire [2:0]   queue_15_deq_bits_segment;
  wire [31:0]  queue_15_deq_bits_readFromScalar;
  wire [11:0]  queue_15_deq_bits_csrInterface_vl;
  wire [11:0]  queue_15_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_15_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_15_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_15_deq_bits_csrInterface_vxrm;
  wire         queue_15_deq_bits_csrInterface_vta;
  wire         queue_15_deq_bits_csrInterface_vma;
  wire         validSink_valid;
  wire [2:0]   validSink_bits_instructionIndex;
  wire         validSink_bits_decodeResult_orderReduce;
  wire         validSink_bits_decodeResult_floatMul;
  wire [1:0]   validSink_bits_decodeResult_fpExecutionType;
  wire         validSink_bits_decodeResult_float;
  wire         validSink_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_bits_decodeResult_topUop;
  wire         validSink_bits_decodeResult_popCount;
  wire         validSink_bits_decodeResult_ffo;
  wire         validSink_bits_decodeResult_average;
  wire         validSink_bits_decodeResult_reverse;
  wire         validSink_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_bits_decodeResult_scheduler;
  wire         validSink_bits_decodeResult_sReadVD;
  wire         validSink_bits_decodeResult_vtype;
  wire         validSink_bits_decodeResult_sWrite;
  wire         validSink_bits_decodeResult_crossRead;
  wire         validSink_bits_decodeResult_crossWrite;
  wire         validSink_bits_decodeResult_maskUnit;
  wire         validSink_bits_decodeResult_special;
  wire         validSink_bits_decodeResult_saturate;
  wire         validSink_bits_decodeResult_vwmacc;
  wire         validSink_bits_decodeResult_readOnly;
  wire         validSink_bits_decodeResult_maskSource;
  wire         validSink_bits_decodeResult_maskDestination;
  wire         validSink_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_bits_decodeResult_uop;
  wire         validSink_bits_decodeResult_iota;
  wire         validSink_bits_decodeResult_mv;
  wire         validSink_bits_decodeResult_extend;
  wire         validSink_bits_decodeResult_unOrderWrite;
  wire         validSink_bits_decodeResult_compress;
  wire         validSink_bits_decodeResult_gather16;
  wire         validSink_bits_decodeResult_gather;
  wire         validSink_bits_decodeResult_slid;
  wire         validSink_bits_decodeResult_targetRd;
  wire         validSink_bits_decodeResult_widenReduce;
  wire         validSink_bits_decodeResult_red;
  wire         validSink_bits_decodeResult_nr;
  wire         validSink_bits_decodeResult_itype;
  wire         validSink_bits_decodeResult_unsigned1;
  wire         validSink_bits_decodeResult_unsigned0;
  wire         validSink_bits_decodeResult_other;
  wire         validSink_bits_decodeResult_multiCycle;
  wire         validSink_bits_decodeResult_divider;
  wire         validSink_bits_decodeResult_multiplier;
  wire         validSink_bits_decodeResult_shift;
  wire         validSink_bits_decodeResult_adder;
  wire         validSink_bits_decodeResult_logic;
  wire         validSink_bits_loadStore;
  wire         validSink_bits_issueInst;
  wire         validSink_bits_store;
  wire         validSink_bits_special;
  wire         validSink_bits_lsWholeReg;
  wire [4:0]   validSink_bits_vs1;
  wire [4:0]   validSink_bits_vs2;
  wire [4:0]   validSink_bits_vd;
  wire [1:0]   validSink_bits_loadStoreEEW;
  wire         validSink_bits_mask;
  wire [2:0]   validSink_bits_segment;
  wire [31:0]  validSink_bits_readFromScalar;
  wire [11:0]  validSink_bits_csrInterface_vl;
  wire [11:0]  validSink_bits_csrInterface_vStart;
  wire [2:0]   validSink_bits_csrInterface_vlmul;
  wire [1:0]   validSink_bits_csrInterface_vSew;
  wire [1:0]   validSink_bits_csrInterface_vxrm;
  wire         validSink_bits_csrInterface_vta;
  wire         validSink_bits_csrInterface_vma;
  wire         laneRequestSinkWire_0_valid = queue_deq_valid;
  wire [2:0]   laneRequestSinkWire_0_bits_instructionIndex = queue_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_0_bits_decodeResult_orderReduce = queue_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_0_bits_decodeResult_floatMul = queue_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_0_bits_decodeResult_fpExecutionType = queue_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_0_bits_decodeResult_float = queue_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_0_bits_decodeResult_specialSlot = queue_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_0_bits_decodeResult_topUop = queue_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_0_bits_decodeResult_popCount = queue_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_0_bits_decodeResult_ffo = queue_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_0_bits_decodeResult_average = queue_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_0_bits_decodeResult_reverse = queue_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_0_bits_decodeResult_dontNeedExecuteInLane = queue_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_0_bits_decodeResult_scheduler = queue_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_0_bits_decodeResult_sReadVD = queue_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_0_bits_decodeResult_vtype = queue_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_0_bits_decodeResult_sWrite = queue_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_crossRead = queue_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_0_bits_decodeResult_crossWrite = queue_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskUnit = queue_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_0_bits_decodeResult_special = queue_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_0_bits_decodeResult_saturate = queue_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_0_bits_decodeResult_vwmacc = queue_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_0_bits_decodeResult_readOnly = queue_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskSource = queue_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskDestination = queue_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskLogic = queue_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_0_bits_decodeResult_uop = queue_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_0_bits_decodeResult_iota = queue_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_0_bits_decodeResult_mv = queue_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_0_bits_decodeResult_extend = queue_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_0_bits_decodeResult_unOrderWrite = queue_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_compress = queue_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_0_bits_decodeResult_gather16 = queue_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_0_bits_decodeResult_gather = queue_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_0_bits_decodeResult_slid = queue_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_0_bits_decodeResult_targetRd = queue_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_0_bits_decodeResult_widenReduce = queue_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_0_bits_decodeResult_red = queue_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_0_bits_decodeResult_nr = queue_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_0_bits_decodeResult_itype = queue_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_0_bits_decodeResult_unsigned1 = queue_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_0_bits_decodeResult_unsigned0 = queue_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_0_bits_decodeResult_other = queue_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_0_bits_decodeResult_multiCycle = queue_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_0_bits_decodeResult_divider = queue_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_0_bits_decodeResult_multiplier = queue_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_0_bits_decodeResult_shift = queue_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_0_bits_decodeResult_adder = queue_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_0_bits_decodeResult_logic = queue_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_0_bits_loadStore = queue_deq_bits_loadStore;
  wire         laneRequestSinkWire_0_bits_issueInst = queue_deq_bits_issueInst;
  wire         laneRequestSinkWire_0_bits_store = queue_deq_bits_store;
  wire         laneRequestSinkWire_0_bits_special = queue_deq_bits_special;
  wire         laneRequestSinkWire_0_bits_lsWholeReg = queue_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_0_bits_vs1 = queue_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_0_bits_vs2 = queue_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_0_bits_vd = queue_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_0_bits_loadStoreEEW = queue_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_0_bits_mask = queue_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_0_bits_segment = queue_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_0_bits_readFromScalar = queue_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_0_bits_csrInterface_vl = queue_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_0_bits_csrInterface_vStart = queue_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_0_bits_csrInterface_vlmul = queue_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_0_bits_csrInterface_vSew = queue_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_0_bits_csrInterface_vxrm = queue_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_0_bits_csrInterface_vta = queue_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_0_bits_csrInterface_vma = queue_deq_bits_csrInterface_vma;
  wire [1:0]   queue_enq_bits_csrInterface_vxrm;
  wire         queue_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi = {queue_enq_bits_csrInterface_vxrm, queue_enq_bits_csrInterface_vta};
  wire         queue_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo = {queue_dataIn_lo_hi, queue_enq_bits_csrInterface_vma};
  wire [2:0]   queue_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo = {queue_enq_bits_csrInterface_vlmul, queue_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_enq_bits_csrInterface_vl;
  wire [11:0]  queue_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi = {queue_enq_bits_csrInterface_vl, queue_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi = {queue_dataIn_hi_hi, queue_dataIn_hi_lo};
  wire         queue_enq_bits_decodeResult_shift;
  wire         queue_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi = {queue_enq_bits_decodeResult_shift, queue_enq_bits_decodeResult_adder};
  wire         queue_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo = {queue_dataIn_lo_lo_lo_lo_hi, queue_enq_bits_decodeResult_logic};
  wire         queue_enq_bits_decodeResult_multiCycle;
  wire         queue_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi = {queue_enq_bits_decodeResult_multiCycle, queue_enq_bits_decodeResult_divider};
  wire         queue_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi = {queue_dataIn_lo_lo_lo_hi_hi, queue_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo = {queue_dataIn_lo_lo_lo_hi, queue_dataIn_lo_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_unsigned1;
  wire         queue_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi = {queue_enq_bits_decodeResult_unsigned1, queue_enq_bits_decodeResult_unsigned0};
  wire         queue_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo = {queue_dataIn_lo_lo_hi_lo_hi, queue_enq_bits_decodeResult_other};
  wire         queue_enq_bits_decodeResult_red;
  wire         queue_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi = {queue_enq_bits_decodeResult_red, queue_enq_bits_decodeResult_nr};
  wire         queue_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi = {queue_dataIn_lo_lo_hi_hi_hi, queue_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi = {queue_dataIn_lo_lo_hi_hi, queue_dataIn_lo_lo_hi_lo};
  wire [11:0]  queue_dataIn_lo_lo = {queue_dataIn_lo_lo_hi, queue_dataIn_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_slid;
  wire         queue_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi = {queue_enq_bits_decodeResult_slid, queue_enq_bits_decodeResult_targetRd};
  wire         queue_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo = {queue_dataIn_lo_hi_lo_lo_hi, queue_enq_bits_decodeResult_widenReduce};
  wire         queue_enq_bits_decodeResult_compress;
  wire         queue_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi = {queue_enq_bits_decodeResult_compress, queue_enq_bits_decodeResult_gather16};
  wire         queue_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi = {queue_dataIn_lo_hi_lo_hi_hi, queue_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo = {queue_dataIn_lo_hi_lo_hi, queue_dataIn_lo_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_mv;
  wire         queue_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi = {queue_enq_bits_decodeResult_mv, queue_enq_bits_decodeResult_extend};
  wire         queue_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo = {queue_dataIn_lo_hi_hi_lo_hi, queue_enq_bits_decodeResult_unOrderWrite};
  wire         queue_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi = {queue_enq_bits_decodeResult_maskLogic, queue_enq_bits_decodeResult_uop};
  wire         queue_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi = {queue_dataIn_lo_hi_hi_hi_hi, queue_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi = {queue_dataIn_lo_hi_hi_hi, queue_dataIn_lo_hi_hi_lo};
  wire [14:0]  queue_dataIn_lo_hi_1 = {queue_dataIn_lo_hi_hi, queue_dataIn_lo_hi_lo};
  wire [26:0]  queue_dataIn_lo_1 = {queue_dataIn_lo_hi_1, queue_dataIn_lo_lo};
  wire         queue_enq_bits_decodeResult_readOnly;
  wire         queue_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi = {queue_enq_bits_decodeResult_readOnly, queue_enq_bits_decodeResult_maskSource};
  wire         queue_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo = {queue_dataIn_hi_lo_lo_lo_hi, queue_enq_bits_decodeResult_maskDestination};
  wire         queue_enq_bits_decodeResult_special;
  wire         queue_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi = {queue_enq_bits_decodeResult_special, queue_enq_bits_decodeResult_saturate};
  wire         queue_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi = {queue_dataIn_hi_lo_lo_hi_hi, queue_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo = {queue_dataIn_hi_lo_lo_hi, queue_dataIn_hi_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_crossRead;
  wire         queue_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi = {queue_enq_bits_decodeResult_crossRead, queue_enq_bits_decodeResult_crossWrite};
  wire         queue_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo = {queue_dataIn_hi_lo_hi_lo_hi, queue_enq_bits_decodeResult_maskUnit};
  wire         queue_enq_bits_decodeResult_sReadVD;
  wire         queue_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi = {queue_enq_bits_decodeResult_sReadVD, queue_enq_bits_decodeResult_vtype};
  wire         queue_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi = {queue_dataIn_hi_lo_hi_hi_hi, queue_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi = {queue_dataIn_hi_lo_hi_hi, queue_dataIn_hi_lo_hi_lo};
  wire [11:0]  queue_dataIn_hi_lo_1 = {queue_dataIn_hi_lo_hi, queue_dataIn_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_reverse;
  wire         queue_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi = {queue_enq_bits_decodeResult_reverse, queue_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo = {queue_dataIn_hi_hi_lo_lo_hi, queue_enq_bits_decodeResult_scheduler};
  wire         queue_enq_bits_decodeResult_popCount;
  wire         queue_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi = {queue_enq_bits_decodeResult_popCount, queue_enq_bits_decodeResult_ffo};
  wire         queue_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi = {queue_dataIn_hi_hi_lo_hi_hi, queue_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo = {queue_dataIn_hi_hi_lo_hi, queue_dataIn_hi_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_float;
  wire         queue_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi = {queue_enq_bits_decodeResult_float, queue_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo = {queue_dataIn_hi_hi_hi_lo_hi, queue_enq_bits_decodeResult_topUop};
  wire         queue_enq_bits_decodeResult_orderReduce;
  wire         queue_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi = {queue_enq_bits_decodeResult_orderReduce, queue_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi = {queue_dataIn_hi_hi_hi_hi_hi, queue_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi = {queue_dataIn_hi_hi_hi_hi, queue_dataIn_hi_hi_hi_lo};
  wire [16:0]  queue_dataIn_hi_hi_1 = {queue_dataIn_hi_hi_hi, queue_dataIn_hi_hi_lo};
  wire [28:0]  queue_dataIn_hi_1 = {queue_dataIn_hi_hi_1, queue_dataIn_hi_lo_1};
  wire [2:0]   queue_enq_bits_segment;
  wire [31:0]  queue_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_1 = {queue_enq_bits_segment, queue_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_1 = {queue_dataIn_lo_lo_hi_1, queue_dataIn_hi, queue_dataIn_lo};
  wire [1:0]   queue_enq_bits_loadStoreEEW;
  wire         queue_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_1 = {queue_enq_bits_loadStoreEEW, queue_enq_bits_mask};
  wire [4:0]   queue_enq_bits_vs2;
  wire [4:0]   queue_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_1 = {queue_enq_bits_vs2, queue_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_2 = {queue_dataIn_lo_hi_hi_1, queue_dataIn_lo_hi_lo_1};
  wire [80:0]  queue_dataIn_lo_2 = {queue_dataIn_lo_hi_2, queue_dataIn_lo_lo_1};
  wire         queue_enq_bits_lsWholeReg;
  wire [4:0]   queue_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_1 = {queue_enq_bits_lsWholeReg, queue_enq_bits_vs1};
  wire         queue_enq_bits_store;
  wire         queue_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_1 = {queue_enq_bits_store, queue_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_2 = {queue_dataIn_hi_lo_hi_1, queue_dataIn_hi_lo_lo_1};
  wire         queue_enq_bits_loadStore;
  wire         queue_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_1 = {queue_enq_bits_loadStore, queue_enq_bits_issueInst};
  wire [2:0]   queue_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_1 = {queue_enq_bits_instructionIndex, queue_dataIn_hi_1, queue_dataIn_lo_1};
  wire [60:0]  queue_dataIn_hi_hi_2 = {queue_dataIn_hi_hi_hi_1, queue_dataIn_hi_hi_lo_1};
  wire [68:0]  queue_dataIn_hi_2 = {queue_dataIn_hi_hi_2, queue_dataIn_hi_lo_2};
  wire [149:0] queue_dataIn = {queue_dataIn_hi_2, queue_dataIn_lo_2};
  wire         queue_dataOut_csrInterface_vma = _queue_fifo_data_out[0];
  wire         queue_dataOut_csrInterface_vta = _queue_fifo_data_out[1];
  wire [1:0]   queue_dataOut_csrInterface_vxrm = _queue_fifo_data_out[3:2];
  wire [1:0]   queue_dataOut_csrInterface_vSew = _queue_fifo_data_out[5:4];
  wire [2:0]   queue_dataOut_csrInterface_vlmul = _queue_fifo_data_out[8:6];
  wire [11:0]  queue_dataOut_csrInterface_vStart = _queue_fifo_data_out[20:9];
  wire [11:0]  queue_dataOut_csrInterface_vl = _queue_fifo_data_out[32:21];
  wire [31:0]  queue_dataOut_readFromScalar = _queue_fifo_data_out[64:33];
  wire [2:0]   queue_dataOut_segment = _queue_fifo_data_out[67:65];
  wire         queue_dataOut_mask = _queue_fifo_data_out[68];
  wire [1:0]   queue_dataOut_loadStoreEEW = _queue_fifo_data_out[70:69];
  wire [4:0]   queue_dataOut_vd = _queue_fifo_data_out[75:71];
  wire [4:0]   queue_dataOut_vs2 = _queue_fifo_data_out[80:76];
  wire [4:0]   queue_dataOut_vs1 = _queue_fifo_data_out[85:81];
  wire         queue_dataOut_lsWholeReg = _queue_fifo_data_out[86];
  wire         queue_dataOut_special = _queue_fifo_data_out[87];
  wire         queue_dataOut_store = _queue_fifo_data_out[88];
  wire         queue_dataOut_issueInst = _queue_fifo_data_out[89];
  wire         queue_dataOut_loadStore = _queue_fifo_data_out[90];
  wire         queue_dataOut_decodeResult_logic = _queue_fifo_data_out[91];
  wire         queue_dataOut_decodeResult_adder = _queue_fifo_data_out[92];
  wire         queue_dataOut_decodeResult_shift = _queue_fifo_data_out[93];
  wire         queue_dataOut_decodeResult_multiplier = _queue_fifo_data_out[94];
  wire         queue_dataOut_decodeResult_divider = _queue_fifo_data_out[95];
  wire         queue_dataOut_decodeResult_multiCycle = _queue_fifo_data_out[96];
  wire         queue_dataOut_decodeResult_other = _queue_fifo_data_out[97];
  wire         queue_dataOut_decodeResult_unsigned0 = _queue_fifo_data_out[98];
  wire         queue_dataOut_decodeResult_unsigned1 = _queue_fifo_data_out[99];
  wire         queue_dataOut_decodeResult_itype = _queue_fifo_data_out[100];
  wire         queue_dataOut_decodeResult_nr = _queue_fifo_data_out[101];
  wire         queue_dataOut_decodeResult_red = _queue_fifo_data_out[102];
  wire         queue_dataOut_decodeResult_widenReduce = _queue_fifo_data_out[103];
  wire         queue_dataOut_decodeResult_targetRd = _queue_fifo_data_out[104];
  wire         queue_dataOut_decodeResult_slid = _queue_fifo_data_out[105];
  wire         queue_dataOut_decodeResult_gather = _queue_fifo_data_out[106];
  wire         queue_dataOut_decodeResult_gather16 = _queue_fifo_data_out[107];
  wire         queue_dataOut_decodeResult_compress = _queue_fifo_data_out[108];
  wire         queue_dataOut_decodeResult_unOrderWrite = _queue_fifo_data_out[109];
  wire         queue_dataOut_decodeResult_extend = _queue_fifo_data_out[110];
  wire         queue_dataOut_decodeResult_mv = _queue_fifo_data_out[111];
  wire         queue_dataOut_decodeResult_iota = _queue_fifo_data_out[112];
  wire [3:0]   queue_dataOut_decodeResult_uop = _queue_fifo_data_out[116:113];
  wire         queue_dataOut_decodeResult_maskLogic = _queue_fifo_data_out[117];
  wire         queue_dataOut_decodeResult_maskDestination = _queue_fifo_data_out[118];
  wire         queue_dataOut_decodeResult_maskSource = _queue_fifo_data_out[119];
  wire         queue_dataOut_decodeResult_readOnly = _queue_fifo_data_out[120];
  wire         queue_dataOut_decodeResult_vwmacc = _queue_fifo_data_out[121];
  wire         queue_dataOut_decodeResult_saturate = _queue_fifo_data_out[122];
  wire         queue_dataOut_decodeResult_special = _queue_fifo_data_out[123];
  wire         queue_dataOut_decodeResult_maskUnit = _queue_fifo_data_out[124];
  wire         queue_dataOut_decodeResult_crossWrite = _queue_fifo_data_out[125];
  wire         queue_dataOut_decodeResult_crossRead = _queue_fifo_data_out[126];
  wire         queue_dataOut_decodeResult_sWrite = _queue_fifo_data_out[127];
  wire         queue_dataOut_decodeResult_vtype = _queue_fifo_data_out[128];
  wire         queue_dataOut_decodeResult_sReadVD = _queue_fifo_data_out[129];
  wire         queue_dataOut_decodeResult_scheduler = _queue_fifo_data_out[130];
  wire         queue_dataOut_decodeResult_dontNeedExecuteInLane = _queue_fifo_data_out[131];
  wire         queue_dataOut_decodeResult_reverse = _queue_fifo_data_out[132];
  wire         queue_dataOut_decodeResult_average = _queue_fifo_data_out[133];
  wire         queue_dataOut_decodeResult_ffo = _queue_fifo_data_out[134];
  wire         queue_dataOut_decodeResult_popCount = _queue_fifo_data_out[135];
  wire [4:0]   queue_dataOut_decodeResult_topUop = _queue_fifo_data_out[140:136];
  wire         queue_dataOut_decodeResult_specialSlot = _queue_fifo_data_out[141];
  wire         queue_dataOut_decodeResult_float = _queue_fifo_data_out[142];
  wire [1:0]   queue_dataOut_decodeResult_fpExecutionType = _queue_fifo_data_out[144:143];
  wire         queue_dataOut_decodeResult_floatMul = _queue_fifo_data_out[145];
  wire         queue_dataOut_decodeResult_orderReduce = _queue_fifo_data_out[146];
  wire [2:0]   queue_dataOut_instructionIndex = _queue_fifo_data_out[149:147];
  wire         queue_enq_ready = ~_queue_fifo_full;
  wire         queue_enq_valid;
  assign queue_deq_valid = ~_queue_fifo_empty | queue_enq_valid;
  assign queue_deq_bits_instructionIndex = _queue_fifo_empty ? queue_enq_bits_instructionIndex : queue_dataOut_instructionIndex;
  assign queue_deq_bits_decodeResult_orderReduce = _queue_fifo_empty ? queue_enq_bits_decodeResult_orderReduce : queue_dataOut_decodeResult_orderReduce;
  assign queue_deq_bits_decodeResult_floatMul = _queue_fifo_empty ? queue_enq_bits_decodeResult_floatMul : queue_dataOut_decodeResult_floatMul;
  assign queue_deq_bits_decodeResult_fpExecutionType = _queue_fifo_empty ? queue_enq_bits_decodeResult_fpExecutionType : queue_dataOut_decodeResult_fpExecutionType;
  assign queue_deq_bits_decodeResult_float = _queue_fifo_empty ? queue_enq_bits_decodeResult_float : queue_dataOut_decodeResult_float;
  assign queue_deq_bits_decodeResult_specialSlot = _queue_fifo_empty ? queue_enq_bits_decodeResult_specialSlot : queue_dataOut_decodeResult_specialSlot;
  assign queue_deq_bits_decodeResult_topUop = _queue_fifo_empty ? queue_enq_bits_decodeResult_topUop : queue_dataOut_decodeResult_topUop;
  assign queue_deq_bits_decodeResult_popCount = _queue_fifo_empty ? queue_enq_bits_decodeResult_popCount : queue_dataOut_decodeResult_popCount;
  assign queue_deq_bits_decodeResult_ffo = _queue_fifo_empty ? queue_enq_bits_decodeResult_ffo : queue_dataOut_decodeResult_ffo;
  assign queue_deq_bits_decodeResult_average = _queue_fifo_empty ? queue_enq_bits_decodeResult_average : queue_dataOut_decodeResult_average;
  assign queue_deq_bits_decodeResult_reverse = _queue_fifo_empty ? queue_enq_bits_decodeResult_reverse : queue_dataOut_decodeResult_reverse;
  assign queue_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_empty ? queue_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_decodeResult_dontNeedExecuteInLane;
  assign queue_deq_bits_decodeResult_scheduler = _queue_fifo_empty ? queue_enq_bits_decodeResult_scheduler : queue_dataOut_decodeResult_scheduler;
  assign queue_deq_bits_decodeResult_sReadVD = _queue_fifo_empty ? queue_enq_bits_decodeResult_sReadVD : queue_dataOut_decodeResult_sReadVD;
  assign queue_deq_bits_decodeResult_vtype = _queue_fifo_empty ? queue_enq_bits_decodeResult_vtype : queue_dataOut_decodeResult_vtype;
  assign queue_deq_bits_decodeResult_sWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_sWrite : queue_dataOut_decodeResult_sWrite;
  assign queue_deq_bits_decodeResult_crossRead = _queue_fifo_empty ? queue_enq_bits_decodeResult_crossRead : queue_dataOut_decodeResult_crossRead;
  assign queue_deq_bits_decodeResult_crossWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_crossWrite : queue_dataOut_decodeResult_crossWrite;
  assign queue_deq_bits_decodeResult_maskUnit = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskUnit : queue_dataOut_decodeResult_maskUnit;
  assign queue_deq_bits_decodeResult_special = _queue_fifo_empty ? queue_enq_bits_decodeResult_special : queue_dataOut_decodeResult_special;
  assign queue_deq_bits_decodeResult_saturate = _queue_fifo_empty ? queue_enq_bits_decodeResult_saturate : queue_dataOut_decodeResult_saturate;
  assign queue_deq_bits_decodeResult_vwmacc = _queue_fifo_empty ? queue_enq_bits_decodeResult_vwmacc : queue_dataOut_decodeResult_vwmacc;
  assign queue_deq_bits_decodeResult_readOnly = _queue_fifo_empty ? queue_enq_bits_decodeResult_readOnly : queue_dataOut_decodeResult_readOnly;
  assign queue_deq_bits_decodeResult_maskSource = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskSource : queue_dataOut_decodeResult_maskSource;
  assign queue_deq_bits_decodeResult_maskDestination = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskDestination : queue_dataOut_decodeResult_maskDestination;
  assign queue_deq_bits_decodeResult_maskLogic = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskLogic : queue_dataOut_decodeResult_maskLogic;
  assign queue_deq_bits_decodeResult_uop = _queue_fifo_empty ? queue_enq_bits_decodeResult_uop : queue_dataOut_decodeResult_uop;
  assign queue_deq_bits_decodeResult_iota = _queue_fifo_empty ? queue_enq_bits_decodeResult_iota : queue_dataOut_decodeResult_iota;
  assign queue_deq_bits_decodeResult_mv = _queue_fifo_empty ? queue_enq_bits_decodeResult_mv : queue_dataOut_decodeResult_mv;
  assign queue_deq_bits_decodeResult_extend = _queue_fifo_empty ? queue_enq_bits_decodeResult_extend : queue_dataOut_decodeResult_extend;
  assign queue_deq_bits_decodeResult_unOrderWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_unOrderWrite : queue_dataOut_decodeResult_unOrderWrite;
  assign queue_deq_bits_decodeResult_compress = _queue_fifo_empty ? queue_enq_bits_decodeResult_compress : queue_dataOut_decodeResult_compress;
  assign queue_deq_bits_decodeResult_gather16 = _queue_fifo_empty ? queue_enq_bits_decodeResult_gather16 : queue_dataOut_decodeResult_gather16;
  assign queue_deq_bits_decodeResult_gather = _queue_fifo_empty ? queue_enq_bits_decodeResult_gather : queue_dataOut_decodeResult_gather;
  assign queue_deq_bits_decodeResult_slid = _queue_fifo_empty ? queue_enq_bits_decodeResult_slid : queue_dataOut_decodeResult_slid;
  assign queue_deq_bits_decodeResult_targetRd = _queue_fifo_empty ? queue_enq_bits_decodeResult_targetRd : queue_dataOut_decodeResult_targetRd;
  assign queue_deq_bits_decodeResult_widenReduce = _queue_fifo_empty ? queue_enq_bits_decodeResult_widenReduce : queue_dataOut_decodeResult_widenReduce;
  assign queue_deq_bits_decodeResult_red = _queue_fifo_empty ? queue_enq_bits_decodeResult_red : queue_dataOut_decodeResult_red;
  assign queue_deq_bits_decodeResult_nr = _queue_fifo_empty ? queue_enq_bits_decodeResult_nr : queue_dataOut_decodeResult_nr;
  assign queue_deq_bits_decodeResult_itype = _queue_fifo_empty ? queue_enq_bits_decodeResult_itype : queue_dataOut_decodeResult_itype;
  assign queue_deq_bits_decodeResult_unsigned1 = _queue_fifo_empty ? queue_enq_bits_decodeResult_unsigned1 : queue_dataOut_decodeResult_unsigned1;
  assign queue_deq_bits_decodeResult_unsigned0 = _queue_fifo_empty ? queue_enq_bits_decodeResult_unsigned0 : queue_dataOut_decodeResult_unsigned0;
  assign queue_deq_bits_decodeResult_other = _queue_fifo_empty ? queue_enq_bits_decodeResult_other : queue_dataOut_decodeResult_other;
  assign queue_deq_bits_decodeResult_multiCycle = _queue_fifo_empty ? queue_enq_bits_decodeResult_multiCycle : queue_dataOut_decodeResult_multiCycle;
  assign queue_deq_bits_decodeResult_divider = _queue_fifo_empty ? queue_enq_bits_decodeResult_divider : queue_dataOut_decodeResult_divider;
  assign queue_deq_bits_decodeResult_multiplier = _queue_fifo_empty ? queue_enq_bits_decodeResult_multiplier : queue_dataOut_decodeResult_multiplier;
  assign queue_deq_bits_decodeResult_shift = _queue_fifo_empty ? queue_enq_bits_decodeResult_shift : queue_dataOut_decodeResult_shift;
  assign queue_deq_bits_decodeResult_adder = _queue_fifo_empty ? queue_enq_bits_decodeResult_adder : queue_dataOut_decodeResult_adder;
  assign queue_deq_bits_decodeResult_logic = _queue_fifo_empty ? queue_enq_bits_decodeResult_logic : queue_dataOut_decodeResult_logic;
  assign queue_deq_bits_loadStore = _queue_fifo_empty ? queue_enq_bits_loadStore : queue_dataOut_loadStore;
  assign queue_deq_bits_issueInst = _queue_fifo_empty ? queue_enq_bits_issueInst : queue_dataOut_issueInst;
  assign queue_deq_bits_store = _queue_fifo_empty ? queue_enq_bits_store : queue_dataOut_store;
  assign queue_deq_bits_special = _queue_fifo_empty ? queue_enq_bits_special : queue_dataOut_special;
  assign queue_deq_bits_lsWholeReg = _queue_fifo_empty ? queue_enq_bits_lsWholeReg : queue_dataOut_lsWholeReg;
  assign queue_deq_bits_vs1 = _queue_fifo_empty ? queue_enq_bits_vs1 : queue_dataOut_vs1;
  assign queue_deq_bits_vs2 = _queue_fifo_empty ? queue_enq_bits_vs2 : queue_dataOut_vs2;
  assign queue_deq_bits_vd = _queue_fifo_empty ? queue_enq_bits_vd : queue_dataOut_vd;
  assign queue_deq_bits_loadStoreEEW = _queue_fifo_empty ? queue_enq_bits_loadStoreEEW : queue_dataOut_loadStoreEEW;
  assign queue_deq_bits_mask = _queue_fifo_empty ? queue_enq_bits_mask : queue_dataOut_mask;
  assign queue_deq_bits_segment = _queue_fifo_empty ? queue_enq_bits_segment : queue_dataOut_segment;
  assign queue_deq_bits_readFromScalar = _queue_fifo_empty ? queue_enq_bits_readFromScalar : queue_dataOut_readFromScalar;
  assign queue_deq_bits_csrInterface_vl = _queue_fifo_empty ? queue_enq_bits_csrInterface_vl : queue_dataOut_csrInterface_vl;
  assign queue_deq_bits_csrInterface_vStart = _queue_fifo_empty ? queue_enq_bits_csrInterface_vStart : queue_dataOut_csrInterface_vStart;
  assign queue_deq_bits_csrInterface_vlmul = _queue_fifo_empty ? queue_enq_bits_csrInterface_vlmul : queue_dataOut_csrInterface_vlmul;
  assign queue_deq_bits_csrInterface_vSew = _queue_fifo_empty ? queue_enq_bits_csrInterface_vSew : queue_dataOut_csrInterface_vSew;
  assign queue_deq_bits_csrInterface_vxrm = _queue_fifo_empty ? queue_enq_bits_csrInterface_vxrm : queue_dataOut_csrInterface_vxrm;
  assign queue_deq_bits_csrInterface_vta = _queue_fifo_empty ? queue_enq_bits_csrInterface_vta : queue_dataOut_csrInterface_vta;
  assign queue_deq_bits_csrInterface_vma = _queue_fifo_empty ? queue_enq_bits_csrInterface_vma : queue_dataOut_csrInterface_vma;
  wire         laneVec_0_laneRequest_bits_issueInst = laneRequestSinkWire_0_ready & laneRequestSinkWire_0_valid;
  reg          releasePipe_pipe_v;
  wire         releasePipe_pipe_out_valid = releasePipe_pipe_v;
  wire         laneRequestSourceWire_0_ready;
  wire         validSource_valid = laneRequestSourceWire_0_ready & laneRequestSourceWire_0_valid;
  reg  [2:0]   tokenCheck_counter;
  wire [2:0]   tokenCheck_counterChange = validSource_valid ? 3'h1 : 3'h7;
  assign tokenCheck = ~(tokenCheck_counter[2]);
  assign laneRequestSourceWire_0_ready = tokenCheck;
  assign queue_enq_valid = validSink_valid;
  assign queue_enq_bits_instructionIndex = validSink_bits_instructionIndex;
  assign queue_enq_bits_decodeResult_orderReduce = validSink_bits_decodeResult_orderReduce;
  assign queue_enq_bits_decodeResult_floatMul = validSink_bits_decodeResult_floatMul;
  assign queue_enq_bits_decodeResult_fpExecutionType = validSink_bits_decodeResult_fpExecutionType;
  assign queue_enq_bits_decodeResult_float = validSink_bits_decodeResult_float;
  assign queue_enq_bits_decodeResult_specialSlot = validSink_bits_decodeResult_specialSlot;
  assign queue_enq_bits_decodeResult_topUop = validSink_bits_decodeResult_topUop;
  assign queue_enq_bits_decodeResult_popCount = validSink_bits_decodeResult_popCount;
  assign queue_enq_bits_decodeResult_ffo = validSink_bits_decodeResult_ffo;
  assign queue_enq_bits_decodeResult_average = validSink_bits_decodeResult_average;
  assign queue_enq_bits_decodeResult_reverse = validSink_bits_decodeResult_reverse;
  assign queue_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_enq_bits_decodeResult_scheduler = validSink_bits_decodeResult_scheduler;
  assign queue_enq_bits_decodeResult_sReadVD = validSink_bits_decodeResult_sReadVD;
  assign queue_enq_bits_decodeResult_vtype = validSink_bits_decodeResult_vtype;
  assign queue_enq_bits_decodeResult_sWrite = validSink_bits_decodeResult_sWrite;
  assign queue_enq_bits_decodeResult_crossRead = validSink_bits_decodeResult_crossRead;
  assign queue_enq_bits_decodeResult_crossWrite = validSink_bits_decodeResult_crossWrite;
  assign queue_enq_bits_decodeResult_maskUnit = validSink_bits_decodeResult_maskUnit;
  assign queue_enq_bits_decodeResult_special = validSink_bits_decodeResult_special;
  assign queue_enq_bits_decodeResult_saturate = validSink_bits_decodeResult_saturate;
  assign queue_enq_bits_decodeResult_vwmacc = validSink_bits_decodeResult_vwmacc;
  assign queue_enq_bits_decodeResult_readOnly = validSink_bits_decodeResult_readOnly;
  assign queue_enq_bits_decodeResult_maskSource = validSink_bits_decodeResult_maskSource;
  assign queue_enq_bits_decodeResult_maskDestination = validSink_bits_decodeResult_maskDestination;
  assign queue_enq_bits_decodeResult_maskLogic = validSink_bits_decodeResult_maskLogic;
  assign queue_enq_bits_decodeResult_uop = validSink_bits_decodeResult_uop;
  assign queue_enq_bits_decodeResult_iota = validSink_bits_decodeResult_iota;
  assign queue_enq_bits_decodeResult_mv = validSink_bits_decodeResult_mv;
  assign queue_enq_bits_decodeResult_extend = validSink_bits_decodeResult_extend;
  assign queue_enq_bits_decodeResult_unOrderWrite = validSink_bits_decodeResult_unOrderWrite;
  assign queue_enq_bits_decodeResult_compress = validSink_bits_decodeResult_compress;
  assign queue_enq_bits_decodeResult_gather16 = validSink_bits_decodeResult_gather16;
  assign queue_enq_bits_decodeResult_gather = validSink_bits_decodeResult_gather;
  assign queue_enq_bits_decodeResult_slid = validSink_bits_decodeResult_slid;
  assign queue_enq_bits_decodeResult_targetRd = validSink_bits_decodeResult_targetRd;
  assign queue_enq_bits_decodeResult_widenReduce = validSink_bits_decodeResult_widenReduce;
  assign queue_enq_bits_decodeResult_red = validSink_bits_decodeResult_red;
  assign queue_enq_bits_decodeResult_nr = validSink_bits_decodeResult_nr;
  assign queue_enq_bits_decodeResult_itype = validSink_bits_decodeResult_itype;
  assign queue_enq_bits_decodeResult_unsigned1 = validSink_bits_decodeResult_unsigned1;
  assign queue_enq_bits_decodeResult_unsigned0 = validSink_bits_decodeResult_unsigned0;
  assign queue_enq_bits_decodeResult_other = validSink_bits_decodeResult_other;
  assign queue_enq_bits_decodeResult_multiCycle = validSink_bits_decodeResult_multiCycle;
  assign queue_enq_bits_decodeResult_divider = validSink_bits_decodeResult_divider;
  assign queue_enq_bits_decodeResult_multiplier = validSink_bits_decodeResult_multiplier;
  assign queue_enq_bits_decodeResult_shift = validSink_bits_decodeResult_shift;
  assign queue_enq_bits_decodeResult_adder = validSink_bits_decodeResult_adder;
  assign queue_enq_bits_decodeResult_logic = validSink_bits_decodeResult_logic;
  assign queue_enq_bits_loadStore = validSink_bits_loadStore;
  assign queue_enq_bits_issueInst = validSink_bits_issueInst;
  assign queue_enq_bits_store = validSink_bits_store;
  assign queue_enq_bits_special = validSink_bits_special;
  assign queue_enq_bits_lsWholeReg = validSink_bits_lsWholeReg;
  assign queue_enq_bits_vs1 = validSink_bits_vs1;
  assign queue_enq_bits_vs2 = validSink_bits_vs2;
  assign queue_enq_bits_vd = validSink_bits_vd;
  assign queue_enq_bits_loadStoreEEW = validSink_bits_loadStoreEEW;
  assign queue_enq_bits_mask = validSink_bits_mask;
  assign queue_enq_bits_segment = validSink_bits_segment;
  assign queue_enq_bits_readFromScalar = validSink_bits_readFromScalar;
  assign queue_enq_bits_csrInterface_vl = validSink_bits_csrInterface_vl;
  assign queue_enq_bits_csrInterface_vStart = validSink_bits_csrInterface_vStart;
  assign queue_enq_bits_csrInterface_vlmul = validSink_bits_csrInterface_vlmul;
  assign queue_enq_bits_csrInterface_vSew = validSink_bits_csrInterface_vSew;
  assign queue_enq_bits_csrInterface_vxrm = validSink_bits_csrInterface_vxrm;
  assign queue_enq_bits_csrInterface_vta = validSink_bits_csrInterface_vta;
  assign queue_enq_bits_csrInterface_vma = validSink_bits_csrInterface_vma;
  reg          shifterReg_0_valid;
  assign validSink_valid = shifterReg_0_valid;
  reg  [2:0]   shifterReg_0_bits_instructionIndex;
  assign validSink_bits_instructionIndex = shifterReg_0_bits_instructionIndex;
  reg          shifterReg_0_bits_decodeResult_orderReduce;
  assign validSink_bits_decodeResult_orderReduce = shifterReg_0_bits_decodeResult_orderReduce;
  reg          shifterReg_0_bits_decodeResult_floatMul;
  assign validSink_bits_decodeResult_floatMul = shifterReg_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_0_bits_decodeResult_fpExecutionType;
  assign validSink_bits_decodeResult_fpExecutionType = shifterReg_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_0_bits_decodeResult_float;
  assign validSink_bits_decodeResult_float = shifterReg_0_bits_decodeResult_float;
  reg          shifterReg_0_bits_decodeResult_specialSlot;
  assign validSink_bits_decodeResult_specialSlot = shifterReg_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_0_bits_decodeResult_topUop;
  assign validSink_bits_decodeResult_topUop = shifterReg_0_bits_decodeResult_topUop;
  reg          shifterReg_0_bits_decodeResult_popCount;
  assign validSink_bits_decodeResult_popCount = shifterReg_0_bits_decodeResult_popCount;
  reg          shifterReg_0_bits_decodeResult_ffo;
  assign validSink_bits_decodeResult_ffo = shifterReg_0_bits_decodeResult_ffo;
  reg          shifterReg_0_bits_decodeResult_average;
  assign validSink_bits_decodeResult_average = shifterReg_0_bits_decodeResult_average;
  reg          shifterReg_0_bits_decodeResult_reverse;
  assign validSink_bits_decodeResult_reverse = shifterReg_0_bits_decodeResult_reverse;
  reg          shifterReg_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_bits_decodeResult_dontNeedExecuteInLane = shifterReg_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_0_bits_decodeResult_scheduler;
  assign validSink_bits_decodeResult_scheduler = shifterReg_0_bits_decodeResult_scheduler;
  reg          shifterReg_0_bits_decodeResult_sReadVD;
  assign validSink_bits_decodeResult_sReadVD = shifterReg_0_bits_decodeResult_sReadVD;
  reg          shifterReg_0_bits_decodeResult_vtype;
  assign validSink_bits_decodeResult_vtype = shifterReg_0_bits_decodeResult_vtype;
  reg          shifterReg_0_bits_decodeResult_sWrite;
  assign validSink_bits_decodeResult_sWrite = shifterReg_0_bits_decodeResult_sWrite;
  reg          shifterReg_0_bits_decodeResult_crossRead;
  assign validSink_bits_decodeResult_crossRead = shifterReg_0_bits_decodeResult_crossRead;
  reg          shifterReg_0_bits_decodeResult_crossWrite;
  assign validSink_bits_decodeResult_crossWrite = shifterReg_0_bits_decodeResult_crossWrite;
  reg          shifterReg_0_bits_decodeResult_maskUnit;
  assign validSink_bits_decodeResult_maskUnit = shifterReg_0_bits_decodeResult_maskUnit;
  reg          shifterReg_0_bits_decodeResult_special;
  assign validSink_bits_decodeResult_special = shifterReg_0_bits_decodeResult_special;
  reg          shifterReg_0_bits_decodeResult_saturate;
  assign validSink_bits_decodeResult_saturate = shifterReg_0_bits_decodeResult_saturate;
  reg          shifterReg_0_bits_decodeResult_vwmacc;
  assign validSink_bits_decodeResult_vwmacc = shifterReg_0_bits_decodeResult_vwmacc;
  reg          shifterReg_0_bits_decodeResult_readOnly;
  assign validSink_bits_decodeResult_readOnly = shifterReg_0_bits_decodeResult_readOnly;
  reg          shifterReg_0_bits_decodeResult_maskSource;
  assign validSink_bits_decodeResult_maskSource = shifterReg_0_bits_decodeResult_maskSource;
  reg          shifterReg_0_bits_decodeResult_maskDestination;
  assign validSink_bits_decodeResult_maskDestination = shifterReg_0_bits_decodeResult_maskDestination;
  reg          shifterReg_0_bits_decodeResult_maskLogic;
  assign validSink_bits_decodeResult_maskLogic = shifterReg_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_0_bits_decodeResult_uop;
  assign validSink_bits_decodeResult_uop = shifterReg_0_bits_decodeResult_uop;
  reg          shifterReg_0_bits_decodeResult_iota;
  assign validSink_bits_decodeResult_iota = shifterReg_0_bits_decodeResult_iota;
  reg          shifterReg_0_bits_decodeResult_mv;
  assign validSink_bits_decodeResult_mv = shifterReg_0_bits_decodeResult_mv;
  reg          shifterReg_0_bits_decodeResult_extend;
  assign validSink_bits_decodeResult_extend = shifterReg_0_bits_decodeResult_extend;
  reg          shifterReg_0_bits_decodeResult_unOrderWrite;
  assign validSink_bits_decodeResult_unOrderWrite = shifterReg_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_0_bits_decodeResult_compress;
  assign validSink_bits_decodeResult_compress = shifterReg_0_bits_decodeResult_compress;
  reg          shifterReg_0_bits_decodeResult_gather16;
  assign validSink_bits_decodeResult_gather16 = shifterReg_0_bits_decodeResult_gather16;
  reg          shifterReg_0_bits_decodeResult_gather;
  assign validSink_bits_decodeResult_gather = shifterReg_0_bits_decodeResult_gather;
  reg          shifterReg_0_bits_decodeResult_slid;
  assign validSink_bits_decodeResult_slid = shifterReg_0_bits_decodeResult_slid;
  reg          shifterReg_0_bits_decodeResult_targetRd;
  assign validSink_bits_decodeResult_targetRd = shifterReg_0_bits_decodeResult_targetRd;
  reg          shifterReg_0_bits_decodeResult_widenReduce;
  assign validSink_bits_decodeResult_widenReduce = shifterReg_0_bits_decodeResult_widenReduce;
  reg          shifterReg_0_bits_decodeResult_red;
  assign validSink_bits_decodeResult_red = shifterReg_0_bits_decodeResult_red;
  reg          shifterReg_0_bits_decodeResult_nr;
  assign validSink_bits_decodeResult_nr = shifterReg_0_bits_decodeResult_nr;
  reg          shifterReg_0_bits_decodeResult_itype;
  assign validSink_bits_decodeResult_itype = shifterReg_0_bits_decodeResult_itype;
  reg          shifterReg_0_bits_decodeResult_unsigned1;
  assign validSink_bits_decodeResult_unsigned1 = shifterReg_0_bits_decodeResult_unsigned1;
  reg          shifterReg_0_bits_decodeResult_unsigned0;
  assign validSink_bits_decodeResult_unsigned0 = shifterReg_0_bits_decodeResult_unsigned0;
  reg          shifterReg_0_bits_decodeResult_other;
  assign validSink_bits_decodeResult_other = shifterReg_0_bits_decodeResult_other;
  reg          shifterReg_0_bits_decodeResult_multiCycle;
  assign validSink_bits_decodeResult_multiCycle = shifterReg_0_bits_decodeResult_multiCycle;
  reg          shifterReg_0_bits_decodeResult_divider;
  assign validSink_bits_decodeResult_divider = shifterReg_0_bits_decodeResult_divider;
  reg          shifterReg_0_bits_decodeResult_multiplier;
  assign validSink_bits_decodeResult_multiplier = shifterReg_0_bits_decodeResult_multiplier;
  reg          shifterReg_0_bits_decodeResult_shift;
  assign validSink_bits_decodeResult_shift = shifterReg_0_bits_decodeResult_shift;
  reg          shifterReg_0_bits_decodeResult_adder;
  assign validSink_bits_decodeResult_adder = shifterReg_0_bits_decodeResult_adder;
  reg          shifterReg_0_bits_decodeResult_logic;
  assign validSink_bits_decodeResult_logic = shifterReg_0_bits_decodeResult_logic;
  reg          shifterReg_0_bits_loadStore;
  assign validSink_bits_loadStore = shifterReg_0_bits_loadStore;
  reg          shifterReg_0_bits_issueInst;
  assign validSink_bits_issueInst = shifterReg_0_bits_issueInst;
  reg          shifterReg_0_bits_store;
  assign validSink_bits_store = shifterReg_0_bits_store;
  reg          shifterReg_0_bits_special;
  assign validSink_bits_special = shifterReg_0_bits_special;
  reg          shifterReg_0_bits_lsWholeReg;
  assign validSink_bits_lsWholeReg = shifterReg_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_0_bits_vs1;
  assign validSink_bits_vs1 = shifterReg_0_bits_vs1;
  reg  [4:0]   shifterReg_0_bits_vs2;
  assign validSink_bits_vs2 = shifterReg_0_bits_vs2;
  reg  [4:0]   shifterReg_0_bits_vd;
  assign validSink_bits_vd = shifterReg_0_bits_vd;
  reg  [1:0]   shifterReg_0_bits_loadStoreEEW;
  assign validSink_bits_loadStoreEEW = shifterReg_0_bits_loadStoreEEW;
  reg          shifterReg_0_bits_mask;
  assign validSink_bits_mask = shifterReg_0_bits_mask;
  reg  [2:0]   shifterReg_0_bits_segment;
  assign validSink_bits_segment = shifterReg_0_bits_segment;
  reg  [31:0]  shifterReg_0_bits_readFromScalar;
  assign validSink_bits_readFromScalar = shifterReg_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_0_bits_csrInterface_vl;
  assign validSink_bits_csrInterface_vl = shifterReg_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_0_bits_csrInterface_vStart;
  assign validSink_bits_csrInterface_vStart = shifterReg_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_0_bits_csrInterface_vlmul;
  assign validSink_bits_csrInterface_vlmul = shifterReg_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_0_bits_csrInterface_vSew;
  assign validSink_bits_csrInterface_vSew = shifterReg_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_0_bits_csrInterface_vxrm;
  assign validSink_bits_csrInterface_vxrm = shifterReg_0_bits_csrInterface_vxrm;
  reg          shifterReg_0_bits_csrInterface_vta;
  assign validSink_bits_csrInterface_vta = shifterReg_0_bits_csrInterface_vta;
  reg          shifterReg_0_bits_csrInterface_vma;
  assign validSink_bits_csrInterface_vma = shifterReg_0_bits_csrInterface_vma;
  wire         shifterValid = shifterReg_0_valid | validSource_valid;
  wire         validSink_1_valid;
  wire [2:0]   validSink_1_bits_instructionIndex;
  wire         validSink_1_bits_decodeResult_orderReduce;
  wire         validSink_1_bits_decodeResult_floatMul;
  wire [1:0]   validSink_1_bits_decodeResult_fpExecutionType;
  wire         validSink_1_bits_decodeResult_float;
  wire         validSink_1_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_1_bits_decodeResult_topUop;
  wire         validSink_1_bits_decodeResult_popCount;
  wire         validSink_1_bits_decodeResult_ffo;
  wire         validSink_1_bits_decodeResult_average;
  wire         validSink_1_bits_decodeResult_reverse;
  wire         validSink_1_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_1_bits_decodeResult_scheduler;
  wire         validSink_1_bits_decodeResult_sReadVD;
  wire         validSink_1_bits_decodeResult_vtype;
  wire         validSink_1_bits_decodeResult_sWrite;
  wire         validSink_1_bits_decodeResult_crossRead;
  wire         validSink_1_bits_decodeResult_crossWrite;
  wire         validSink_1_bits_decodeResult_maskUnit;
  wire         validSink_1_bits_decodeResult_special;
  wire         validSink_1_bits_decodeResult_saturate;
  wire         validSink_1_bits_decodeResult_vwmacc;
  wire         validSink_1_bits_decodeResult_readOnly;
  wire         validSink_1_bits_decodeResult_maskSource;
  wire         validSink_1_bits_decodeResult_maskDestination;
  wire         validSink_1_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_1_bits_decodeResult_uop;
  wire         validSink_1_bits_decodeResult_iota;
  wire         validSink_1_bits_decodeResult_mv;
  wire         validSink_1_bits_decodeResult_extend;
  wire         validSink_1_bits_decodeResult_unOrderWrite;
  wire         validSink_1_bits_decodeResult_compress;
  wire         validSink_1_bits_decodeResult_gather16;
  wire         validSink_1_bits_decodeResult_gather;
  wire         validSink_1_bits_decodeResult_slid;
  wire         validSink_1_bits_decodeResult_targetRd;
  wire         validSink_1_bits_decodeResult_widenReduce;
  wire         validSink_1_bits_decodeResult_red;
  wire         validSink_1_bits_decodeResult_nr;
  wire         validSink_1_bits_decodeResult_itype;
  wire         validSink_1_bits_decodeResult_unsigned1;
  wire         validSink_1_bits_decodeResult_unsigned0;
  wire         validSink_1_bits_decodeResult_other;
  wire         validSink_1_bits_decodeResult_multiCycle;
  wire         validSink_1_bits_decodeResult_divider;
  wire         validSink_1_bits_decodeResult_multiplier;
  wire         validSink_1_bits_decodeResult_shift;
  wire         validSink_1_bits_decodeResult_adder;
  wire         validSink_1_bits_decodeResult_logic;
  wire         validSink_1_bits_loadStore;
  wire         validSink_1_bits_issueInst;
  wire         validSink_1_bits_store;
  wire         validSink_1_bits_special;
  wire         validSink_1_bits_lsWholeReg;
  wire [4:0]   validSink_1_bits_vs1;
  wire [4:0]   validSink_1_bits_vs2;
  wire [4:0]   validSink_1_bits_vd;
  wire [1:0]   validSink_1_bits_loadStoreEEW;
  wire         validSink_1_bits_mask;
  wire [2:0]   validSink_1_bits_segment;
  wire [31:0]  validSink_1_bits_readFromScalar;
  wire [11:0]  validSink_1_bits_csrInterface_vl;
  wire [11:0]  validSink_1_bits_csrInterface_vStart;
  wire [2:0]   validSink_1_bits_csrInterface_vlmul;
  wire [1:0]   validSink_1_bits_csrInterface_vSew;
  wire [1:0]   validSink_1_bits_csrInterface_vxrm;
  wire         validSink_1_bits_csrInterface_vta;
  wire         validSink_1_bits_csrInterface_vma;
  wire         laneRequestSinkWire_1_valid = queue_1_deq_valid;
  wire [2:0]   laneRequestSinkWire_1_bits_instructionIndex = queue_1_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_1_bits_decodeResult_orderReduce = queue_1_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_1_bits_decodeResult_floatMul = queue_1_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_1_bits_decodeResult_fpExecutionType = queue_1_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_1_bits_decodeResult_float = queue_1_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_1_bits_decodeResult_specialSlot = queue_1_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_1_bits_decodeResult_topUop = queue_1_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_1_bits_decodeResult_popCount = queue_1_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_1_bits_decodeResult_ffo = queue_1_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_1_bits_decodeResult_average = queue_1_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_1_bits_decodeResult_reverse = queue_1_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_1_bits_decodeResult_dontNeedExecuteInLane = queue_1_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_1_bits_decodeResult_scheduler = queue_1_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_1_bits_decodeResult_sReadVD = queue_1_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_1_bits_decodeResult_vtype = queue_1_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_1_bits_decodeResult_sWrite = queue_1_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_crossRead = queue_1_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_1_bits_decodeResult_crossWrite = queue_1_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskUnit = queue_1_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_1_bits_decodeResult_special = queue_1_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_1_bits_decodeResult_saturate = queue_1_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_1_bits_decodeResult_vwmacc = queue_1_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_1_bits_decodeResult_readOnly = queue_1_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskSource = queue_1_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskDestination = queue_1_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskLogic = queue_1_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_1_bits_decodeResult_uop = queue_1_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_1_bits_decodeResult_iota = queue_1_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_1_bits_decodeResult_mv = queue_1_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_1_bits_decodeResult_extend = queue_1_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_1_bits_decodeResult_unOrderWrite = queue_1_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_compress = queue_1_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_1_bits_decodeResult_gather16 = queue_1_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_1_bits_decodeResult_gather = queue_1_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_1_bits_decodeResult_slid = queue_1_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_1_bits_decodeResult_targetRd = queue_1_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_1_bits_decodeResult_widenReduce = queue_1_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_1_bits_decodeResult_red = queue_1_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_1_bits_decodeResult_nr = queue_1_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_1_bits_decodeResult_itype = queue_1_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_1_bits_decodeResult_unsigned1 = queue_1_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_1_bits_decodeResult_unsigned0 = queue_1_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_1_bits_decodeResult_other = queue_1_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_1_bits_decodeResult_multiCycle = queue_1_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_1_bits_decodeResult_divider = queue_1_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_1_bits_decodeResult_multiplier = queue_1_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_1_bits_decodeResult_shift = queue_1_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_1_bits_decodeResult_adder = queue_1_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_1_bits_decodeResult_logic = queue_1_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_1_bits_loadStore = queue_1_deq_bits_loadStore;
  wire         laneRequestSinkWire_1_bits_issueInst = queue_1_deq_bits_issueInst;
  wire         laneRequestSinkWire_1_bits_store = queue_1_deq_bits_store;
  wire         laneRequestSinkWire_1_bits_special = queue_1_deq_bits_special;
  wire         laneRequestSinkWire_1_bits_lsWholeReg = queue_1_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_1_bits_vs1 = queue_1_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_1_bits_vs2 = queue_1_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_1_bits_vd = queue_1_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_1_bits_loadStoreEEW = queue_1_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_1_bits_mask = queue_1_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_1_bits_segment = queue_1_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_1_bits_readFromScalar = queue_1_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_1_bits_csrInterface_vl = queue_1_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_1_bits_csrInterface_vStart = queue_1_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_1_bits_csrInterface_vlmul = queue_1_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_1_bits_csrInterface_vSew = queue_1_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_1_bits_csrInterface_vxrm = queue_1_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_1_bits_csrInterface_vta = queue_1_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_1_bits_csrInterface_vma = queue_1_deq_bits_csrInterface_vma;
  wire [1:0]   queue_1_enq_bits_csrInterface_vxrm;
  wire         queue_1_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_3 = {queue_1_enq_bits_csrInterface_vxrm, queue_1_enq_bits_csrInterface_vta};
  wire         queue_1_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_3 = {queue_dataIn_lo_hi_3, queue_1_enq_bits_csrInterface_vma};
  wire [2:0]   queue_1_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_1_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_3 = {queue_1_enq_bits_csrInterface_vlmul, queue_1_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_1_enq_bits_csrInterface_vl;
  wire [11:0]  queue_1_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_3 = {queue_1_enq_bits_csrInterface_vl, queue_1_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_3 = {queue_dataIn_hi_hi_3, queue_dataIn_hi_lo_3};
  wire         queue_1_enq_bits_decodeResult_shift;
  wire         queue_1_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_1 = {queue_1_enq_bits_decodeResult_shift, queue_1_enq_bits_decodeResult_adder};
  wire         queue_1_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_1 = {queue_dataIn_lo_lo_lo_lo_hi_1, queue_1_enq_bits_decodeResult_logic};
  wire         queue_1_enq_bits_decodeResult_multiCycle;
  wire         queue_1_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_multiCycle, queue_1_enq_bits_decodeResult_divider};
  wire         queue_1_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_1 = {queue_dataIn_lo_lo_lo_hi_hi_1, queue_1_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_1 = {queue_dataIn_lo_lo_lo_hi_1, queue_dataIn_lo_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_unsigned1;
  wire         queue_1_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_unsigned1, queue_1_enq_bits_decodeResult_unsigned0};
  wire         queue_1_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_1 = {queue_dataIn_lo_lo_hi_lo_hi_1, queue_1_enq_bits_decodeResult_other};
  wire         queue_1_enq_bits_decodeResult_red;
  wire         queue_1_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_red, queue_1_enq_bits_decodeResult_nr};
  wire         queue_1_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_1 = {queue_dataIn_lo_lo_hi_hi_hi_1, queue_1_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_2 = {queue_dataIn_lo_lo_hi_hi_1, queue_dataIn_lo_lo_hi_lo_1};
  wire [11:0]  queue_dataIn_lo_lo_2 = {queue_dataIn_lo_lo_hi_2, queue_dataIn_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_slid;
  wire         queue_1_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_1 = {queue_1_enq_bits_decodeResult_slid, queue_1_enq_bits_decodeResult_targetRd};
  wire         queue_1_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_1 = {queue_dataIn_lo_hi_lo_lo_hi_1, queue_1_enq_bits_decodeResult_widenReduce};
  wire         queue_1_enq_bits_decodeResult_compress;
  wire         queue_1_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_compress, queue_1_enq_bits_decodeResult_gather16};
  wire         queue_1_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_1 = {queue_dataIn_lo_hi_lo_hi_hi_1, queue_1_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_2 = {queue_dataIn_lo_hi_lo_hi_1, queue_dataIn_lo_hi_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_mv;
  wire         queue_1_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_mv, queue_1_enq_bits_decodeResult_extend};
  wire         queue_1_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_1 = {queue_dataIn_lo_hi_hi_lo_hi_1, queue_1_enq_bits_decodeResult_unOrderWrite};
  wire         queue_1_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_1_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_maskLogic, queue_1_enq_bits_decodeResult_uop};
  wire         queue_1_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_1 = {queue_dataIn_lo_hi_hi_hi_hi_1, queue_1_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_2 = {queue_dataIn_lo_hi_hi_hi_1, queue_dataIn_lo_hi_hi_lo_1};
  wire [14:0]  queue_dataIn_lo_hi_4 = {queue_dataIn_lo_hi_hi_2, queue_dataIn_lo_hi_lo_2};
  wire [26:0]  queue_dataIn_lo_4 = {queue_dataIn_lo_hi_4, queue_dataIn_lo_lo_2};
  wire         queue_1_enq_bits_decodeResult_readOnly;
  wire         queue_1_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_1 = {queue_1_enq_bits_decodeResult_readOnly, queue_1_enq_bits_decodeResult_maskSource};
  wire         queue_1_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_1 = {queue_dataIn_hi_lo_lo_lo_hi_1, queue_1_enq_bits_decodeResult_maskDestination};
  wire         queue_1_enq_bits_decodeResult_special;
  wire         queue_1_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_special, queue_1_enq_bits_decodeResult_saturate};
  wire         queue_1_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_1 = {queue_dataIn_hi_lo_lo_hi_hi_1, queue_1_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_2 = {queue_dataIn_hi_lo_lo_hi_1, queue_dataIn_hi_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_crossRead;
  wire         queue_1_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_crossRead, queue_1_enq_bits_decodeResult_crossWrite};
  wire         queue_1_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_1 = {queue_dataIn_hi_lo_hi_lo_hi_1, queue_1_enq_bits_decodeResult_maskUnit};
  wire         queue_1_enq_bits_decodeResult_sReadVD;
  wire         queue_1_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_sReadVD, queue_1_enq_bits_decodeResult_vtype};
  wire         queue_1_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_1 = {queue_dataIn_hi_lo_hi_hi_hi_1, queue_1_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_2 = {queue_dataIn_hi_lo_hi_hi_1, queue_dataIn_hi_lo_hi_lo_1};
  wire [11:0]  queue_dataIn_hi_lo_4 = {queue_dataIn_hi_lo_hi_2, queue_dataIn_hi_lo_lo_2};
  wire         queue_1_enq_bits_decodeResult_reverse;
  wire         queue_1_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_1 = {queue_1_enq_bits_decodeResult_reverse, queue_1_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_1_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_1 = {queue_dataIn_hi_hi_lo_lo_hi_1, queue_1_enq_bits_decodeResult_scheduler};
  wire         queue_1_enq_bits_decodeResult_popCount;
  wire         queue_1_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_popCount, queue_1_enq_bits_decodeResult_ffo};
  wire         queue_1_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_1 = {queue_dataIn_hi_hi_lo_hi_hi_1, queue_1_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_2 = {queue_dataIn_hi_hi_lo_hi_1, queue_dataIn_hi_hi_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_float;
  wire         queue_1_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_float, queue_1_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_1_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_1 = {queue_dataIn_hi_hi_hi_lo_hi_1, queue_1_enq_bits_decodeResult_topUop};
  wire         queue_1_enq_bits_decodeResult_orderReduce;
  wire         queue_1_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_orderReduce, queue_1_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_1_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_1 = {queue_dataIn_hi_hi_hi_hi_hi_1, queue_1_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_2 = {queue_dataIn_hi_hi_hi_hi_1, queue_dataIn_hi_hi_hi_lo_1};
  wire [16:0]  queue_dataIn_hi_hi_4 = {queue_dataIn_hi_hi_hi_2, queue_dataIn_hi_hi_lo_2};
  wire [28:0]  queue_dataIn_hi_4 = {queue_dataIn_hi_hi_4, queue_dataIn_hi_lo_4};
  wire [2:0]   queue_1_enq_bits_segment;
  wire [31:0]  queue_1_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_3 = {queue_1_enq_bits_segment, queue_1_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_3 = {queue_dataIn_lo_lo_hi_3, queue_dataIn_hi_3, queue_dataIn_lo_3};
  wire [1:0]   queue_1_enq_bits_loadStoreEEW;
  wire         queue_1_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_3 = {queue_1_enq_bits_loadStoreEEW, queue_1_enq_bits_mask};
  wire [4:0]   queue_1_enq_bits_vs2;
  wire [4:0]   queue_1_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_3 = {queue_1_enq_bits_vs2, queue_1_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_5 = {queue_dataIn_lo_hi_hi_3, queue_dataIn_lo_hi_lo_3};
  wire [80:0]  queue_dataIn_lo_5 = {queue_dataIn_lo_hi_5, queue_dataIn_lo_lo_3};
  wire         queue_1_enq_bits_lsWholeReg;
  wire [4:0]   queue_1_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_3 = {queue_1_enq_bits_lsWholeReg, queue_1_enq_bits_vs1};
  wire         queue_1_enq_bits_store;
  wire         queue_1_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_3 = {queue_1_enq_bits_store, queue_1_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_5 = {queue_dataIn_hi_lo_hi_3, queue_dataIn_hi_lo_lo_3};
  wire         queue_1_enq_bits_loadStore;
  wire         queue_1_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_3 = {queue_1_enq_bits_loadStore, queue_1_enq_bits_issueInst};
  wire [2:0]   queue_1_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_3 = {queue_1_enq_bits_instructionIndex, queue_dataIn_hi_4, queue_dataIn_lo_4};
  wire [60:0]  queue_dataIn_hi_hi_5 = {queue_dataIn_hi_hi_hi_3, queue_dataIn_hi_hi_lo_3};
  wire [68:0]  queue_dataIn_hi_5 = {queue_dataIn_hi_hi_5, queue_dataIn_hi_lo_5};
  wire [149:0] queue_dataIn_1 = {queue_dataIn_hi_5, queue_dataIn_lo_5};
  wire         queue_dataOut_1_csrInterface_vma = _queue_fifo_1_data_out[0];
  wire         queue_dataOut_1_csrInterface_vta = _queue_fifo_1_data_out[1];
  wire [1:0]   queue_dataOut_1_csrInterface_vxrm = _queue_fifo_1_data_out[3:2];
  wire [1:0]   queue_dataOut_1_csrInterface_vSew = _queue_fifo_1_data_out[5:4];
  wire [2:0]   queue_dataOut_1_csrInterface_vlmul = _queue_fifo_1_data_out[8:6];
  wire [11:0]  queue_dataOut_1_csrInterface_vStart = _queue_fifo_1_data_out[20:9];
  wire [11:0]  queue_dataOut_1_csrInterface_vl = _queue_fifo_1_data_out[32:21];
  wire [31:0]  queue_dataOut_1_readFromScalar = _queue_fifo_1_data_out[64:33];
  wire [2:0]   queue_dataOut_1_segment = _queue_fifo_1_data_out[67:65];
  wire         queue_dataOut_1_mask = _queue_fifo_1_data_out[68];
  wire [1:0]   queue_dataOut_1_loadStoreEEW = _queue_fifo_1_data_out[70:69];
  wire [4:0]   queue_dataOut_1_vd = _queue_fifo_1_data_out[75:71];
  wire [4:0]   queue_dataOut_1_vs2 = _queue_fifo_1_data_out[80:76];
  wire [4:0]   queue_dataOut_1_vs1 = _queue_fifo_1_data_out[85:81];
  wire         queue_dataOut_1_lsWholeReg = _queue_fifo_1_data_out[86];
  wire         queue_dataOut_1_special = _queue_fifo_1_data_out[87];
  wire         queue_dataOut_1_store = _queue_fifo_1_data_out[88];
  wire         queue_dataOut_1_issueInst = _queue_fifo_1_data_out[89];
  wire         queue_dataOut_1_loadStore = _queue_fifo_1_data_out[90];
  wire         queue_dataOut_1_decodeResult_logic = _queue_fifo_1_data_out[91];
  wire         queue_dataOut_1_decodeResult_adder = _queue_fifo_1_data_out[92];
  wire         queue_dataOut_1_decodeResult_shift = _queue_fifo_1_data_out[93];
  wire         queue_dataOut_1_decodeResult_multiplier = _queue_fifo_1_data_out[94];
  wire         queue_dataOut_1_decodeResult_divider = _queue_fifo_1_data_out[95];
  wire         queue_dataOut_1_decodeResult_multiCycle = _queue_fifo_1_data_out[96];
  wire         queue_dataOut_1_decodeResult_other = _queue_fifo_1_data_out[97];
  wire         queue_dataOut_1_decodeResult_unsigned0 = _queue_fifo_1_data_out[98];
  wire         queue_dataOut_1_decodeResult_unsigned1 = _queue_fifo_1_data_out[99];
  wire         queue_dataOut_1_decodeResult_itype = _queue_fifo_1_data_out[100];
  wire         queue_dataOut_1_decodeResult_nr = _queue_fifo_1_data_out[101];
  wire         queue_dataOut_1_decodeResult_red = _queue_fifo_1_data_out[102];
  wire         queue_dataOut_1_decodeResult_widenReduce = _queue_fifo_1_data_out[103];
  wire         queue_dataOut_1_decodeResult_targetRd = _queue_fifo_1_data_out[104];
  wire         queue_dataOut_1_decodeResult_slid = _queue_fifo_1_data_out[105];
  wire         queue_dataOut_1_decodeResult_gather = _queue_fifo_1_data_out[106];
  wire         queue_dataOut_1_decodeResult_gather16 = _queue_fifo_1_data_out[107];
  wire         queue_dataOut_1_decodeResult_compress = _queue_fifo_1_data_out[108];
  wire         queue_dataOut_1_decodeResult_unOrderWrite = _queue_fifo_1_data_out[109];
  wire         queue_dataOut_1_decodeResult_extend = _queue_fifo_1_data_out[110];
  wire         queue_dataOut_1_decodeResult_mv = _queue_fifo_1_data_out[111];
  wire         queue_dataOut_1_decodeResult_iota = _queue_fifo_1_data_out[112];
  wire [3:0]   queue_dataOut_1_decodeResult_uop = _queue_fifo_1_data_out[116:113];
  wire         queue_dataOut_1_decodeResult_maskLogic = _queue_fifo_1_data_out[117];
  wire         queue_dataOut_1_decodeResult_maskDestination = _queue_fifo_1_data_out[118];
  wire         queue_dataOut_1_decodeResult_maskSource = _queue_fifo_1_data_out[119];
  wire         queue_dataOut_1_decodeResult_readOnly = _queue_fifo_1_data_out[120];
  wire         queue_dataOut_1_decodeResult_vwmacc = _queue_fifo_1_data_out[121];
  wire         queue_dataOut_1_decodeResult_saturate = _queue_fifo_1_data_out[122];
  wire         queue_dataOut_1_decodeResult_special = _queue_fifo_1_data_out[123];
  wire         queue_dataOut_1_decodeResult_maskUnit = _queue_fifo_1_data_out[124];
  wire         queue_dataOut_1_decodeResult_crossWrite = _queue_fifo_1_data_out[125];
  wire         queue_dataOut_1_decodeResult_crossRead = _queue_fifo_1_data_out[126];
  wire         queue_dataOut_1_decodeResult_sWrite = _queue_fifo_1_data_out[127];
  wire         queue_dataOut_1_decodeResult_vtype = _queue_fifo_1_data_out[128];
  wire         queue_dataOut_1_decodeResult_sReadVD = _queue_fifo_1_data_out[129];
  wire         queue_dataOut_1_decodeResult_scheduler = _queue_fifo_1_data_out[130];
  wire         queue_dataOut_1_decodeResult_dontNeedExecuteInLane = _queue_fifo_1_data_out[131];
  wire         queue_dataOut_1_decodeResult_reverse = _queue_fifo_1_data_out[132];
  wire         queue_dataOut_1_decodeResult_average = _queue_fifo_1_data_out[133];
  wire         queue_dataOut_1_decodeResult_ffo = _queue_fifo_1_data_out[134];
  wire         queue_dataOut_1_decodeResult_popCount = _queue_fifo_1_data_out[135];
  wire [4:0]   queue_dataOut_1_decodeResult_topUop = _queue_fifo_1_data_out[140:136];
  wire         queue_dataOut_1_decodeResult_specialSlot = _queue_fifo_1_data_out[141];
  wire         queue_dataOut_1_decodeResult_float = _queue_fifo_1_data_out[142];
  wire [1:0]   queue_dataOut_1_decodeResult_fpExecutionType = _queue_fifo_1_data_out[144:143];
  wire         queue_dataOut_1_decodeResult_floatMul = _queue_fifo_1_data_out[145];
  wire         queue_dataOut_1_decodeResult_orderReduce = _queue_fifo_1_data_out[146];
  wire [2:0]   queue_dataOut_1_instructionIndex = _queue_fifo_1_data_out[149:147];
  wire         queue_1_enq_ready = ~_queue_fifo_1_full;
  wire         queue_1_enq_valid;
  assign queue_1_deq_valid = ~_queue_fifo_1_empty | queue_1_enq_valid;
  assign queue_1_deq_bits_instructionIndex = _queue_fifo_1_empty ? queue_1_enq_bits_instructionIndex : queue_dataOut_1_instructionIndex;
  assign queue_1_deq_bits_decodeResult_orderReduce = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_orderReduce : queue_dataOut_1_decodeResult_orderReduce;
  assign queue_1_deq_bits_decodeResult_floatMul = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_floatMul : queue_dataOut_1_decodeResult_floatMul;
  assign queue_1_deq_bits_decodeResult_fpExecutionType = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_fpExecutionType : queue_dataOut_1_decodeResult_fpExecutionType;
  assign queue_1_deq_bits_decodeResult_float = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_float : queue_dataOut_1_decodeResult_float;
  assign queue_1_deq_bits_decodeResult_specialSlot = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_specialSlot : queue_dataOut_1_decodeResult_specialSlot;
  assign queue_1_deq_bits_decodeResult_topUop = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_topUop : queue_dataOut_1_decodeResult_topUop;
  assign queue_1_deq_bits_decodeResult_popCount = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_popCount : queue_dataOut_1_decodeResult_popCount;
  assign queue_1_deq_bits_decodeResult_ffo = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_ffo : queue_dataOut_1_decodeResult_ffo;
  assign queue_1_deq_bits_decodeResult_average = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_average : queue_dataOut_1_decodeResult_average;
  assign queue_1_deq_bits_decodeResult_reverse = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_reverse : queue_dataOut_1_decodeResult_reverse;
  assign queue_1_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_1_decodeResult_dontNeedExecuteInLane;
  assign queue_1_deq_bits_decodeResult_scheduler = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_scheduler : queue_dataOut_1_decodeResult_scheduler;
  assign queue_1_deq_bits_decodeResult_sReadVD = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_sReadVD : queue_dataOut_1_decodeResult_sReadVD;
  assign queue_1_deq_bits_decodeResult_vtype = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_vtype : queue_dataOut_1_decodeResult_vtype;
  assign queue_1_deq_bits_decodeResult_sWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_sWrite : queue_dataOut_1_decodeResult_sWrite;
  assign queue_1_deq_bits_decodeResult_crossRead = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_crossRead : queue_dataOut_1_decodeResult_crossRead;
  assign queue_1_deq_bits_decodeResult_crossWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_crossWrite : queue_dataOut_1_decodeResult_crossWrite;
  assign queue_1_deq_bits_decodeResult_maskUnit = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskUnit : queue_dataOut_1_decodeResult_maskUnit;
  assign queue_1_deq_bits_decodeResult_special = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_special : queue_dataOut_1_decodeResult_special;
  assign queue_1_deq_bits_decodeResult_saturate = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_saturate : queue_dataOut_1_decodeResult_saturate;
  assign queue_1_deq_bits_decodeResult_vwmacc = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_vwmacc : queue_dataOut_1_decodeResult_vwmacc;
  assign queue_1_deq_bits_decodeResult_readOnly = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_readOnly : queue_dataOut_1_decodeResult_readOnly;
  assign queue_1_deq_bits_decodeResult_maskSource = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskSource : queue_dataOut_1_decodeResult_maskSource;
  assign queue_1_deq_bits_decodeResult_maskDestination = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskDestination : queue_dataOut_1_decodeResult_maskDestination;
  assign queue_1_deq_bits_decodeResult_maskLogic = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskLogic : queue_dataOut_1_decodeResult_maskLogic;
  assign queue_1_deq_bits_decodeResult_uop = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_uop : queue_dataOut_1_decodeResult_uop;
  assign queue_1_deq_bits_decodeResult_iota = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_iota : queue_dataOut_1_decodeResult_iota;
  assign queue_1_deq_bits_decodeResult_mv = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_mv : queue_dataOut_1_decodeResult_mv;
  assign queue_1_deq_bits_decodeResult_extend = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_extend : queue_dataOut_1_decodeResult_extend;
  assign queue_1_deq_bits_decodeResult_unOrderWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unOrderWrite : queue_dataOut_1_decodeResult_unOrderWrite;
  assign queue_1_deq_bits_decodeResult_compress = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_compress : queue_dataOut_1_decodeResult_compress;
  assign queue_1_deq_bits_decodeResult_gather16 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_gather16 : queue_dataOut_1_decodeResult_gather16;
  assign queue_1_deq_bits_decodeResult_gather = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_gather : queue_dataOut_1_decodeResult_gather;
  assign queue_1_deq_bits_decodeResult_slid = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_slid : queue_dataOut_1_decodeResult_slid;
  assign queue_1_deq_bits_decodeResult_targetRd = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_targetRd : queue_dataOut_1_decodeResult_targetRd;
  assign queue_1_deq_bits_decodeResult_widenReduce = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_widenReduce : queue_dataOut_1_decodeResult_widenReduce;
  assign queue_1_deq_bits_decodeResult_red = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_red : queue_dataOut_1_decodeResult_red;
  assign queue_1_deq_bits_decodeResult_nr = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_nr : queue_dataOut_1_decodeResult_nr;
  assign queue_1_deq_bits_decodeResult_itype = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_itype : queue_dataOut_1_decodeResult_itype;
  assign queue_1_deq_bits_decodeResult_unsigned1 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unsigned1 : queue_dataOut_1_decodeResult_unsigned1;
  assign queue_1_deq_bits_decodeResult_unsigned0 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unsigned0 : queue_dataOut_1_decodeResult_unsigned0;
  assign queue_1_deq_bits_decodeResult_other = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_other : queue_dataOut_1_decodeResult_other;
  assign queue_1_deq_bits_decodeResult_multiCycle = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_multiCycle : queue_dataOut_1_decodeResult_multiCycle;
  assign queue_1_deq_bits_decodeResult_divider = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_divider : queue_dataOut_1_decodeResult_divider;
  assign queue_1_deq_bits_decodeResult_multiplier = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_multiplier : queue_dataOut_1_decodeResult_multiplier;
  assign queue_1_deq_bits_decodeResult_shift = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_shift : queue_dataOut_1_decodeResult_shift;
  assign queue_1_deq_bits_decodeResult_adder = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_adder : queue_dataOut_1_decodeResult_adder;
  assign queue_1_deq_bits_decodeResult_logic = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_logic : queue_dataOut_1_decodeResult_logic;
  assign queue_1_deq_bits_loadStore = _queue_fifo_1_empty ? queue_1_enq_bits_loadStore : queue_dataOut_1_loadStore;
  assign queue_1_deq_bits_issueInst = _queue_fifo_1_empty ? queue_1_enq_bits_issueInst : queue_dataOut_1_issueInst;
  assign queue_1_deq_bits_store = _queue_fifo_1_empty ? queue_1_enq_bits_store : queue_dataOut_1_store;
  assign queue_1_deq_bits_special = _queue_fifo_1_empty ? queue_1_enq_bits_special : queue_dataOut_1_special;
  assign queue_1_deq_bits_lsWholeReg = _queue_fifo_1_empty ? queue_1_enq_bits_lsWholeReg : queue_dataOut_1_lsWholeReg;
  assign queue_1_deq_bits_vs1 = _queue_fifo_1_empty ? queue_1_enq_bits_vs1 : queue_dataOut_1_vs1;
  assign queue_1_deq_bits_vs2 = _queue_fifo_1_empty ? queue_1_enq_bits_vs2 : queue_dataOut_1_vs2;
  assign queue_1_deq_bits_vd = _queue_fifo_1_empty ? queue_1_enq_bits_vd : queue_dataOut_1_vd;
  assign queue_1_deq_bits_loadStoreEEW = _queue_fifo_1_empty ? queue_1_enq_bits_loadStoreEEW : queue_dataOut_1_loadStoreEEW;
  assign queue_1_deq_bits_mask = _queue_fifo_1_empty ? queue_1_enq_bits_mask : queue_dataOut_1_mask;
  assign queue_1_deq_bits_segment = _queue_fifo_1_empty ? queue_1_enq_bits_segment : queue_dataOut_1_segment;
  assign queue_1_deq_bits_readFromScalar = _queue_fifo_1_empty ? queue_1_enq_bits_readFromScalar : queue_dataOut_1_readFromScalar;
  assign queue_1_deq_bits_csrInterface_vl = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vl : queue_dataOut_1_csrInterface_vl;
  assign queue_1_deq_bits_csrInterface_vStart = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vStart : queue_dataOut_1_csrInterface_vStart;
  assign queue_1_deq_bits_csrInterface_vlmul = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vlmul : queue_dataOut_1_csrInterface_vlmul;
  assign queue_1_deq_bits_csrInterface_vSew = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vSew : queue_dataOut_1_csrInterface_vSew;
  assign queue_1_deq_bits_csrInterface_vxrm = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vxrm : queue_dataOut_1_csrInterface_vxrm;
  assign queue_1_deq_bits_csrInterface_vta = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vta : queue_dataOut_1_csrInterface_vta;
  assign queue_1_deq_bits_csrInterface_vma = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vma : queue_dataOut_1_csrInterface_vma;
  wire         laneVec_1_laneRequest_bits_issueInst = laneRequestSinkWire_1_ready & laneRequestSinkWire_1_valid;
  reg          releasePipe_pipe_v_1;
  wire         releasePipe_pipe_out_1_valid = releasePipe_pipe_v_1;
  wire         laneRequestSourceWire_1_ready;
  wire         validSource_1_valid = laneRequestSourceWire_1_ready & laneRequestSourceWire_1_valid;
  reg  [2:0]   tokenCheck_counter_1;
  wire [2:0]   tokenCheck_counterChange_1 = validSource_1_valid ? 3'h1 : 3'h7;
  assign tokenCheck_1 = ~(tokenCheck_counter_1[2]);
  assign laneRequestSourceWire_1_ready = tokenCheck_1;
  assign queue_1_enq_valid = validSink_1_valid;
  assign queue_1_enq_bits_instructionIndex = validSink_1_bits_instructionIndex;
  assign queue_1_enq_bits_decodeResult_orderReduce = validSink_1_bits_decodeResult_orderReduce;
  assign queue_1_enq_bits_decodeResult_floatMul = validSink_1_bits_decodeResult_floatMul;
  assign queue_1_enq_bits_decodeResult_fpExecutionType = validSink_1_bits_decodeResult_fpExecutionType;
  assign queue_1_enq_bits_decodeResult_float = validSink_1_bits_decodeResult_float;
  assign queue_1_enq_bits_decodeResult_specialSlot = validSink_1_bits_decodeResult_specialSlot;
  assign queue_1_enq_bits_decodeResult_topUop = validSink_1_bits_decodeResult_topUop;
  assign queue_1_enq_bits_decodeResult_popCount = validSink_1_bits_decodeResult_popCount;
  assign queue_1_enq_bits_decodeResult_ffo = validSink_1_bits_decodeResult_ffo;
  assign queue_1_enq_bits_decodeResult_average = validSink_1_bits_decodeResult_average;
  assign queue_1_enq_bits_decodeResult_reverse = validSink_1_bits_decodeResult_reverse;
  assign queue_1_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_1_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_1_enq_bits_decodeResult_scheduler = validSink_1_bits_decodeResult_scheduler;
  assign queue_1_enq_bits_decodeResult_sReadVD = validSink_1_bits_decodeResult_sReadVD;
  assign queue_1_enq_bits_decodeResult_vtype = validSink_1_bits_decodeResult_vtype;
  assign queue_1_enq_bits_decodeResult_sWrite = validSink_1_bits_decodeResult_sWrite;
  assign queue_1_enq_bits_decodeResult_crossRead = validSink_1_bits_decodeResult_crossRead;
  assign queue_1_enq_bits_decodeResult_crossWrite = validSink_1_bits_decodeResult_crossWrite;
  assign queue_1_enq_bits_decodeResult_maskUnit = validSink_1_bits_decodeResult_maskUnit;
  assign queue_1_enq_bits_decodeResult_special = validSink_1_bits_decodeResult_special;
  assign queue_1_enq_bits_decodeResult_saturate = validSink_1_bits_decodeResult_saturate;
  assign queue_1_enq_bits_decodeResult_vwmacc = validSink_1_bits_decodeResult_vwmacc;
  assign queue_1_enq_bits_decodeResult_readOnly = validSink_1_bits_decodeResult_readOnly;
  assign queue_1_enq_bits_decodeResult_maskSource = validSink_1_bits_decodeResult_maskSource;
  assign queue_1_enq_bits_decodeResult_maskDestination = validSink_1_bits_decodeResult_maskDestination;
  assign queue_1_enq_bits_decodeResult_maskLogic = validSink_1_bits_decodeResult_maskLogic;
  assign queue_1_enq_bits_decodeResult_uop = validSink_1_bits_decodeResult_uop;
  assign queue_1_enq_bits_decodeResult_iota = validSink_1_bits_decodeResult_iota;
  assign queue_1_enq_bits_decodeResult_mv = validSink_1_bits_decodeResult_mv;
  assign queue_1_enq_bits_decodeResult_extend = validSink_1_bits_decodeResult_extend;
  assign queue_1_enq_bits_decodeResult_unOrderWrite = validSink_1_bits_decodeResult_unOrderWrite;
  assign queue_1_enq_bits_decodeResult_compress = validSink_1_bits_decodeResult_compress;
  assign queue_1_enq_bits_decodeResult_gather16 = validSink_1_bits_decodeResult_gather16;
  assign queue_1_enq_bits_decodeResult_gather = validSink_1_bits_decodeResult_gather;
  assign queue_1_enq_bits_decodeResult_slid = validSink_1_bits_decodeResult_slid;
  assign queue_1_enq_bits_decodeResult_targetRd = validSink_1_bits_decodeResult_targetRd;
  assign queue_1_enq_bits_decodeResult_widenReduce = validSink_1_bits_decodeResult_widenReduce;
  assign queue_1_enq_bits_decodeResult_red = validSink_1_bits_decodeResult_red;
  assign queue_1_enq_bits_decodeResult_nr = validSink_1_bits_decodeResult_nr;
  assign queue_1_enq_bits_decodeResult_itype = validSink_1_bits_decodeResult_itype;
  assign queue_1_enq_bits_decodeResult_unsigned1 = validSink_1_bits_decodeResult_unsigned1;
  assign queue_1_enq_bits_decodeResult_unsigned0 = validSink_1_bits_decodeResult_unsigned0;
  assign queue_1_enq_bits_decodeResult_other = validSink_1_bits_decodeResult_other;
  assign queue_1_enq_bits_decodeResult_multiCycle = validSink_1_bits_decodeResult_multiCycle;
  assign queue_1_enq_bits_decodeResult_divider = validSink_1_bits_decodeResult_divider;
  assign queue_1_enq_bits_decodeResult_multiplier = validSink_1_bits_decodeResult_multiplier;
  assign queue_1_enq_bits_decodeResult_shift = validSink_1_bits_decodeResult_shift;
  assign queue_1_enq_bits_decodeResult_adder = validSink_1_bits_decodeResult_adder;
  assign queue_1_enq_bits_decodeResult_logic = validSink_1_bits_decodeResult_logic;
  assign queue_1_enq_bits_loadStore = validSink_1_bits_loadStore;
  assign queue_1_enq_bits_issueInst = validSink_1_bits_issueInst;
  assign queue_1_enq_bits_store = validSink_1_bits_store;
  assign queue_1_enq_bits_special = validSink_1_bits_special;
  assign queue_1_enq_bits_lsWholeReg = validSink_1_bits_lsWholeReg;
  assign queue_1_enq_bits_vs1 = validSink_1_bits_vs1;
  assign queue_1_enq_bits_vs2 = validSink_1_bits_vs2;
  assign queue_1_enq_bits_vd = validSink_1_bits_vd;
  assign queue_1_enq_bits_loadStoreEEW = validSink_1_bits_loadStoreEEW;
  assign queue_1_enq_bits_mask = validSink_1_bits_mask;
  assign queue_1_enq_bits_segment = validSink_1_bits_segment;
  assign queue_1_enq_bits_readFromScalar = validSink_1_bits_readFromScalar;
  assign queue_1_enq_bits_csrInterface_vl = validSink_1_bits_csrInterface_vl;
  assign queue_1_enq_bits_csrInterface_vStart = validSink_1_bits_csrInterface_vStart;
  assign queue_1_enq_bits_csrInterface_vlmul = validSink_1_bits_csrInterface_vlmul;
  assign queue_1_enq_bits_csrInterface_vSew = validSink_1_bits_csrInterface_vSew;
  assign queue_1_enq_bits_csrInterface_vxrm = validSink_1_bits_csrInterface_vxrm;
  assign queue_1_enq_bits_csrInterface_vta = validSink_1_bits_csrInterface_vta;
  assign queue_1_enq_bits_csrInterface_vma = validSink_1_bits_csrInterface_vma;
  reg          shifterReg_1_0_valid;
  assign validSink_1_valid = shifterReg_1_0_valid;
  reg  [2:0]   shifterReg_1_0_bits_instructionIndex;
  assign validSink_1_bits_instructionIndex = shifterReg_1_0_bits_instructionIndex;
  reg          shifterReg_1_0_bits_decodeResult_orderReduce;
  assign validSink_1_bits_decodeResult_orderReduce = shifterReg_1_0_bits_decodeResult_orderReduce;
  reg          shifterReg_1_0_bits_decodeResult_floatMul;
  assign validSink_1_bits_decodeResult_floatMul = shifterReg_1_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_1_0_bits_decodeResult_fpExecutionType;
  assign validSink_1_bits_decodeResult_fpExecutionType = shifterReg_1_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_1_0_bits_decodeResult_float;
  assign validSink_1_bits_decodeResult_float = shifterReg_1_0_bits_decodeResult_float;
  reg          shifterReg_1_0_bits_decodeResult_specialSlot;
  assign validSink_1_bits_decodeResult_specialSlot = shifterReg_1_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_1_0_bits_decodeResult_topUop;
  assign validSink_1_bits_decodeResult_topUop = shifterReg_1_0_bits_decodeResult_topUop;
  reg          shifterReg_1_0_bits_decodeResult_popCount;
  assign validSink_1_bits_decodeResult_popCount = shifterReg_1_0_bits_decodeResult_popCount;
  reg          shifterReg_1_0_bits_decodeResult_ffo;
  assign validSink_1_bits_decodeResult_ffo = shifterReg_1_0_bits_decodeResult_ffo;
  reg          shifterReg_1_0_bits_decodeResult_average;
  assign validSink_1_bits_decodeResult_average = shifterReg_1_0_bits_decodeResult_average;
  reg          shifterReg_1_0_bits_decodeResult_reverse;
  assign validSink_1_bits_decodeResult_reverse = shifterReg_1_0_bits_decodeResult_reverse;
  reg          shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_1_bits_decodeResult_dontNeedExecuteInLane = shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_1_0_bits_decodeResult_scheduler;
  assign validSink_1_bits_decodeResult_scheduler = shifterReg_1_0_bits_decodeResult_scheduler;
  reg          shifterReg_1_0_bits_decodeResult_sReadVD;
  assign validSink_1_bits_decodeResult_sReadVD = shifterReg_1_0_bits_decodeResult_sReadVD;
  reg          shifterReg_1_0_bits_decodeResult_vtype;
  assign validSink_1_bits_decodeResult_vtype = shifterReg_1_0_bits_decodeResult_vtype;
  reg          shifterReg_1_0_bits_decodeResult_sWrite;
  assign validSink_1_bits_decodeResult_sWrite = shifterReg_1_0_bits_decodeResult_sWrite;
  reg          shifterReg_1_0_bits_decodeResult_crossRead;
  assign validSink_1_bits_decodeResult_crossRead = shifterReg_1_0_bits_decodeResult_crossRead;
  reg          shifterReg_1_0_bits_decodeResult_crossWrite;
  assign validSink_1_bits_decodeResult_crossWrite = shifterReg_1_0_bits_decodeResult_crossWrite;
  reg          shifterReg_1_0_bits_decodeResult_maskUnit;
  assign validSink_1_bits_decodeResult_maskUnit = shifterReg_1_0_bits_decodeResult_maskUnit;
  reg          shifterReg_1_0_bits_decodeResult_special;
  assign validSink_1_bits_decodeResult_special = shifterReg_1_0_bits_decodeResult_special;
  reg          shifterReg_1_0_bits_decodeResult_saturate;
  assign validSink_1_bits_decodeResult_saturate = shifterReg_1_0_bits_decodeResult_saturate;
  reg          shifterReg_1_0_bits_decodeResult_vwmacc;
  assign validSink_1_bits_decodeResult_vwmacc = shifterReg_1_0_bits_decodeResult_vwmacc;
  reg          shifterReg_1_0_bits_decodeResult_readOnly;
  assign validSink_1_bits_decodeResult_readOnly = shifterReg_1_0_bits_decodeResult_readOnly;
  reg          shifterReg_1_0_bits_decodeResult_maskSource;
  assign validSink_1_bits_decodeResult_maskSource = shifterReg_1_0_bits_decodeResult_maskSource;
  reg          shifterReg_1_0_bits_decodeResult_maskDestination;
  assign validSink_1_bits_decodeResult_maskDestination = shifterReg_1_0_bits_decodeResult_maskDestination;
  reg          shifterReg_1_0_bits_decodeResult_maskLogic;
  assign validSink_1_bits_decodeResult_maskLogic = shifterReg_1_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_1_0_bits_decodeResult_uop;
  assign validSink_1_bits_decodeResult_uop = shifterReg_1_0_bits_decodeResult_uop;
  reg          shifterReg_1_0_bits_decodeResult_iota;
  assign validSink_1_bits_decodeResult_iota = shifterReg_1_0_bits_decodeResult_iota;
  reg          shifterReg_1_0_bits_decodeResult_mv;
  assign validSink_1_bits_decodeResult_mv = shifterReg_1_0_bits_decodeResult_mv;
  reg          shifterReg_1_0_bits_decodeResult_extend;
  assign validSink_1_bits_decodeResult_extend = shifterReg_1_0_bits_decodeResult_extend;
  reg          shifterReg_1_0_bits_decodeResult_unOrderWrite;
  assign validSink_1_bits_decodeResult_unOrderWrite = shifterReg_1_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_1_0_bits_decodeResult_compress;
  assign validSink_1_bits_decodeResult_compress = shifterReg_1_0_bits_decodeResult_compress;
  reg          shifterReg_1_0_bits_decodeResult_gather16;
  assign validSink_1_bits_decodeResult_gather16 = shifterReg_1_0_bits_decodeResult_gather16;
  reg          shifterReg_1_0_bits_decodeResult_gather;
  assign validSink_1_bits_decodeResult_gather = shifterReg_1_0_bits_decodeResult_gather;
  reg          shifterReg_1_0_bits_decodeResult_slid;
  assign validSink_1_bits_decodeResult_slid = shifterReg_1_0_bits_decodeResult_slid;
  reg          shifterReg_1_0_bits_decodeResult_targetRd;
  assign validSink_1_bits_decodeResult_targetRd = shifterReg_1_0_bits_decodeResult_targetRd;
  reg          shifterReg_1_0_bits_decodeResult_widenReduce;
  assign validSink_1_bits_decodeResult_widenReduce = shifterReg_1_0_bits_decodeResult_widenReduce;
  reg          shifterReg_1_0_bits_decodeResult_red;
  assign validSink_1_bits_decodeResult_red = shifterReg_1_0_bits_decodeResult_red;
  reg          shifterReg_1_0_bits_decodeResult_nr;
  assign validSink_1_bits_decodeResult_nr = shifterReg_1_0_bits_decodeResult_nr;
  reg          shifterReg_1_0_bits_decodeResult_itype;
  assign validSink_1_bits_decodeResult_itype = shifterReg_1_0_bits_decodeResult_itype;
  reg          shifterReg_1_0_bits_decodeResult_unsigned1;
  assign validSink_1_bits_decodeResult_unsigned1 = shifterReg_1_0_bits_decodeResult_unsigned1;
  reg          shifterReg_1_0_bits_decodeResult_unsigned0;
  assign validSink_1_bits_decodeResult_unsigned0 = shifterReg_1_0_bits_decodeResult_unsigned0;
  reg          shifterReg_1_0_bits_decodeResult_other;
  assign validSink_1_bits_decodeResult_other = shifterReg_1_0_bits_decodeResult_other;
  reg          shifterReg_1_0_bits_decodeResult_multiCycle;
  assign validSink_1_bits_decodeResult_multiCycle = shifterReg_1_0_bits_decodeResult_multiCycle;
  reg          shifterReg_1_0_bits_decodeResult_divider;
  assign validSink_1_bits_decodeResult_divider = shifterReg_1_0_bits_decodeResult_divider;
  reg          shifterReg_1_0_bits_decodeResult_multiplier;
  assign validSink_1_bits_decodeResult_multiplier = shifterReg_1_0_bits_decodeResult_multiplier;
  reg          shifterReg_1_0_bits_decodeResult_shift;
  assign validSink_1_bits_decodeResult_shift = shifterReg_1_0_bits_decodeResult_shift;
  reg          shifterReg_1_0_bits_decodeResult_adder;
  assign validSink_1_bits_decodeResult_adder = shifterReg_1_0_bits_decodeResult_adder;
  reg          shifterReg_1_0_bits_decodeResult_logic;
  assign validSink_1_bits_decodeResult_logic = shifterReg_1_0_bits_decodeResult_logic;
  reg          shifterReg_1_0_bits_loadStore;
  assign validSink_1_bits_loadStore = shifterReg_1_0_bits_loadStore;
  reg          shifterReg_1_0_bits_issueInst;
  assign validSink_1_bits_issueInst = shifterReg_1_0_bits_issueInst;
  reg          shifterReg_1_0_bits_store;
  assign validSink_1_bits_store = shifterReg_1_0_bits_store;
  reg          shifterReg_1_0_bits_special;
  assign validSink_1_bits_special = shifterReg_1_0_bits_special;
  reg          shifterReg_1_0_bits_lsWholeReg;
  assign validSink_1_bits_lsWholeReg = shifterReg_1_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_1_0_bits_vs1;
  assign validSink_1_bits_vs1 = shifterReg_1_0_bits_vs1;
  reg  [4:0]   shifterReg_1_0_bits_vs2;
  assign validSink_1_bits_vs2 = shifterReg_1_0_bits_vs2;
  reg  [4:0]   shifterReg_1_0_bits_vd;
  assign validSink_1_bits_vd = shifterReg_1_0_bits_vd;
  reg  [1:0]   shifterReg_1_0_bits_loadStoreEEW;
  assign validSink_1_bits_loadStoreEEW = shifterReg_1_0_bits_loadStoreEEW;
  reg          shifterReg_1_0_bits_mask;
  assign validSink_1_bits_mask = shifterReg_1_0_bits_mask;
  reg  [2:0]   shifterReg_1_0_bits_segment;
  assign validSink_1_bits_segment = shifterReg_1_0_bits_segment;
  reg  [31:0]  shifterReg_1_0_bits_readFromScalar;
  assign validSink_1_bits_readFromScalar = shifterReg_1_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_1_0_bits_csrInterface_vl;
  assign validSink_1_bits_csrInterface_vl = shifterReg_1_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_1_0_bits_csrInterface_vStart;
  assign validSink_1_bits_csrInterface_vStart = shifterReg_1_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_1_0_bits_csrInterface_vlmul;
  assign validSink_1_bits_csrInterface_vlmul = shifterReg_1_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_1_0_bits_csrInterface_vSew;
  assign validSink_1_bits_csrInterface_vSew = shifterReg_1_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_1_0_bits_csrInterface_vxrm;
  assign validSink_1_bits_csrInterface_vxrm = shifterReg_1_0_bits_csrInterface_vxrm;
  reg          shifterReg_1_0_bits_csrInterface_vta;
  assign validSink_1_bits_csrInterface_vta = shifterReg_1_0_bits_csrInterface_vta;
  reg          shifterReg_1_0_bits_csrInterface_vma;
  assign validSink_1_bits_csrInterface_vma = shifterReg_1_0_bits_csrInterface_vma;
  wire         shifterValid_1 = shifterReg_1_0_valid | validSource_1_valid;
  wire         validSink_2_valid;
  wire [2:0]   validSink_2_bits_instructionIndex;
  wire         validSink_2_bits_decodeResult_orderReduce;
  wire         validSink_2_bits_decodeResult_floatMul;
  wire [1:0]   validSink_2_bits_decodeResult_fpExecutionType;
  wire         validSink_2_bits_decodeResult_float;
  wire         validSink_2_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_2_bits_decodeResult_topUop;
  wire         validSink_2_bits_decodeResult_popCount;
  wire         validSink_2_bits_decodeResult_ffo;
  wire         validSink_2_bits_decodeResult_average;
  wire         validSink_2_bits_decodeResult_reverse;
  wire         validSink_2_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_2_bits_decodeResult_scheduler;
  wire         validSink_2_bits_decodeResult_sReadVD;
  wire         validSink_2_bits_decodeResult_vtype;
  wire         validSink_2_bits_decodeResult_sWrite;
  wire         validSink_2_bits_decodeResult_crossRead;
  wire         validSink_2_bits_decodeResult_crossWrite;
  wire         validSink_2_bits_decodeResult_maskUnit;
  wire         validSink_2_bits_decodeResult_special;
  wire         validSink_2_bits_decodeResult_saturate;
  wire         validSink_2_bits_decodeResult_vwmacc;
  wire         validSink_2_bits_decodeResult_readOnly;
  wire         validSink_2_bits_decodeResult_maskSource;
  wire         validSink_2_bits_decodeResult_maskDestination;
  wire         validSink_2_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_2_bits_decodeResult_uop;
  wire         validSink_2_bits_decodeResult_iota;
  wire         validSink_2_bits_decodeResult_mv;
  wire         validSink_2_bits_decodeResult_extend;
  wire         validSink_2_bits_decodeResult_unOrderWrite;
  wire         validSink_2_bits_decodeResult_compress;
  wire         validSink_2_bits_decodeResult_gather16;
  wire         validSink_2_bits_decodeResult_gather;
  wire         validSink_2_bits_decodeResult_slid;
  wire         validSink_2_bits_decodeResult_targetRd;
  wire         validSink_2_bits_decodeResult_widenReduce;
  wire         validSink_2_bits_decodeResult_red;
  wire         validSink_2_bits_decodeResult_nr;
  wire         validSink_2_bits_decodeResult_itype;
  wire         validSink_2_bits_decodeResult_unsigned1;
  wire         validSink_2_bits_decodeResult_unsigned0;
  wire         validSink_2_bits_decodeResult_other;
  wire         validSink_2_bits_decodeResult_multiCycle;
  wire         validSink_2_bits_decodeResult_divider;
  wire         validSink_2_bits_decodeResult_multiplier;
  wire         validSink_2_bits_decodeResult_shift;
  wire         validSink_2_bits_decodeResult_adder;
  wire         validSink_2_bits_decodeResult_logic;
  wire         validSink_2_bits_loadStore;
  wire         validSink_2_bits_issueInst;
  wire         validSink_2_bits_store;
  wire         validSink_2_bits_special;
  wire         validSink_2_bits_lsWholeReg;
  wire [4:0]   validSink_2_bits_vs1;
  wire [4:0]   validSink_2_bits_vs2;
  wire [4:0]   validSink_2_bits_vd;
  wire [1:0]   validSink_2_bits_loadStoreEEW;
  wire         validSink_2_bits_mask;
  wire [2:0]   validSink_2_bits_segment;
  wire [31:0]  validSink_2_bits_readFromScalar;
  wire [11:0]  validSink_2_bits_csrInterface_vl;
  wire [11:0]  validSink_2_bits_csrInterface_vStart;
  wire [2:0]   validSink_2_bits_csrInterface_vlmul;
  wire [1:0]   validSink_2_bits_csrInterface_vSew;
  wire [1:0]   validSink_2_bits_csrInterface_vxrm;
  wire         validSink_2_bits_csrInterface_vta;
  wire         validSink_2_bits_csrInterface_vma;
  wire         laneRequestSinkWire_2_valid = queue_2_deq_valid;
  wire [2:0]   laneRequestSinkWire_2_bits_instructionIndex = queue_2_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_2_bits_decodeResult_orderReduce = queue_2_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_2_bits_decodeResult_floatMul = queue_2_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_2_bits_decodeResult_fpExecutionType = queue_2_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_2_bits_decodeResult_float = queue_2_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_2_bits_decodeResult_specialSlot = queue_2_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_2_bits_decodeResult_topUop = queue_2_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_2_bits_decodeResult_popCount = queue_2_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_2_bits_decodeResult_ffo = queue_2_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_2_bits_decodeResult_average = queue_2_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_2_bits_decodeResult_reverse = queue_2_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_2_bits_decodeResult_dontNeedExecuteInLane = queue_2_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_2_bits_decodeResult_scheduler = queue_2_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_2_bits_decodeResult_sReadVD = queue_2_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_2_bits_decodeResult_vtype = queue_2_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_2_bits_decodeResult_sWrite = queue_2_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_crossRead = queue_2_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_2_bits_decodeResult_crossWrite = queue_2_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskUnit = queue_2_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_2_bits_decodeResult_special = queue_2_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_2_bits_decodeResult_saturate = queue_2_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_2_bits_decodeResult_vwmacc = queue_2_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_2_bits_decodeResult_readOnly = queue_2_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskSource = queue_2_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskDestination = queue_2_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskLogic = queue_2_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_2_bits_decodeResult_uop = queue_2_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_2_bits_decodeResult_iota = queue_2_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_2_bits_decodeResult_mv = queue_2_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_2_bits_decodeResult_extend = queue_2_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_2_bits_decodeResult_unOrderWrite = queue_2_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_compress = queue_2_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_2_bits_decodeResult_gather16 = queue_2_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_2_bits_decodeResult_gather = queue_2_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_2_bits_decodeResult_slid = queue_2_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_2_bits_decodeResult_targetRd = queue_2_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_2_bits_decodeResult_widenReduce = queue_2_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_2_bits_decodeResult_red = queue_2_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_2_bits_decodeResult_nr = queue_2_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_2_bits_decodeResult_itype = queue_2_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_2_bits_decodeResult_unsigned1 = queue_2_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_2_bits_decodeResult_unsigned0 = queue_2_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_2_bits_decodeResult_other = queue_2_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_2_bits_decodeResult_multiCycle = queue_2_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_2_bits_decodeResult_divider = queue_2_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_2_bits_decodeResult_multiplier = queue_2_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_2_bits_decodeResult_shift = queue_2_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_2_bits_decodeResult_adder = queue_2_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_2_bits_decodeResult_logic = queue_2_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_2_bits_loadStore = queue_2_deq_bits_loadStore;
  wire         laneRequestSinkWire_2_bits_issueInst = queue_2_deq_bits_issueInst;
  wire         laneRequestSinkWire_2_bits_store = queue_2_deq_bits_store;
  wire         laneRequestSinkWire_2_bits_special = queue_2_deq_bits_special;
  wire         laneRequestSinkWire_2_bits_lsWholeReg = queue_2_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_2_bits_vs1 = queue_2_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_2_bits_vs2 = queue_2_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_2_bits_vd = queue_2_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_2_bits_loadStoreEEW = queue_2_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_2_bits_mask = queue_2_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_2_bits_segment = queue_2_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_2_bits_readFromScalar = queue_2_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_2_bits_csrInterface_vl = queue_2_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_2_bits_csrInterface_vStart = queue_2_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_2_bits_csrInterface_vlmul = queue_2_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_2_bits_csrInterface_vSew = queue_2_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_2_bits_csrInterface_vxrm = queue_2_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_2_bits_csrInterface_vta = queue_2_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_2_bits_csrInterface_vma = queue_2_deq_bits_csrInterface_vma;
  wire [1:0]   queue_2_enq_bits_csrInterface_vxrm;
  wire         queue_2_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_6 = {queue_2_enq_bits_csrInterface_vxrm, queue_2_enq_bits_csrInterface_vta};
  wire         queue_2_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_6 = {queue_dataIn_lo_hi_6, queue_2_enq_bits_csrInterface_vma};
  wire [2:0]   queue_2_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_2_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_6 = {queue_2_enq_bits_csrInterface_vlmul, queue_2_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_2_enq_bits_csrInterface_vl;
  wire [11:0]  queue_2_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_6 = {queue_2_enq_bits_csrInterface_vl, queue_2_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_6 = {queue_dataIn_hi_hi_6, queue_dataIn_hi_lo_6};
  wire         queue_2_enq_bits_decodeResult_shift;
  wire         queue_2_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_2 = {queue_2_enq_bits_decodeResult_shift, queue_2_enq_bits_decodeResult_adder};
  wire         queue_2_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_2 = {queue_dataIn_lo_lo_lo_lo_hi_2, queue_2_enq_bits_decodeResult_logic};
  wire         queue_2_enq_bits_decodeResult_multiCycle;
  wire         queue_2_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_multiCycle, queue_2_enq_bits_decodeResult_divider};
  wire         queue_2_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_2 = {queue_dataIn_lo_lo_lo_hi_hi_2, queue_2_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_2 = {queue_dataIn_lo_lo_lo_hi_2, queue_dataIn_lo_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_unsigned1;
  wire         queue_2_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_unsigned1, queue_2_enq_bits_decodeResult_unsigned0};
  wire         queue_2_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_2 = {queue_dataIn_lo_lo_hi_lo_hi_2, queue_2_enq_bits_decodeResult_other};
  wire         queue_2_enq_bits_decodeResult_red;
  wire         queue_2_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_red, queue_2_enq_bits_decodeResult_nr};
  wire         queue_2_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_2 = {queue_dataIn_lo_lo_hi_hi_hi_2, queue_2_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_4 = {queue_dataIn_lo_lo_hi_hi_2, queue_dataIn_lo_lo_hi_lo_2};
  wire [11:0]  queue_dataIn_lo_lo_4 = {queue_dataIn_lo_lo_hi_4, queue_dataIn_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_slid;
  wire         queue_2_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_2 = {queue_2_enq_bits_decodeResult_slid, queue_2_enq_bits_decodeResult_targetRd};
  wire         queue_2_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_2 = {queue_dataIn_lo_hi_lo_lo_hi_2, queue_2_enq_bits_decodeResult_widenReduce};
  wire         queue_2_enq_bits_decodeResult_compress;
  wire         queue_2_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_compress, queue_2_enq_bits_decodeResult_gather16};
  wire         queue_2_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_2 = {queue_dataIn_lo_hi_lo_hi_hi_2, queue_2_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_4 = {queue_dataIn_lo_hi_lo_hi_2, queue_dataIn_lo_hi_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_mv;
  wire         queue_2_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_mv, queue_2_enq_bits_decodeResult_extend};
  wire         queue_2_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_2 = {queue_dataIn_lo_hi_hi_lo_hi_2, queue_2_enq_bits_decodeResult_unOrderWrite};
  wire         queue_2_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_2_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_maskLogic, queue_2_enq_bits_decodeResult_uop};
  wire         queue_2_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_2 = {queue_dataIn_lo_hi_hi_hi_hi_2, queue_2_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_4 = {queue_dataIn_lo_hi_hi_hi_2, queue_dataIn_lo_hi_hi_lo_2};
  wire [14:0]  queue_dataIn_lo_hi_7 = {queue_dataIn_lo_hi_hi_4, queue_dataIn_lo_hi_lo_4};
  wire [26:0]  queue_dataIn_lo_7 = {queue_dataIn_lo_hi_7, queue_dataIn_lo_lo_4};
  wire         queue_2_enq_bits_decodeResult_readOnly;
  wire         queue_2_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_2 = {queue_2_enq_bits_decodeResult_readOnly, queue_2_enq_bits_decodeResult_maskSource};
  wire         queue_2_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_2 = {queue_dataIn_hi_lo_lo_lo_hi_2, queue_2_enq_bits_decodeResult_maskDestination};
  wire         queue_2_enq_bits_decodeResult_special;
  wire         queue_2_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_special, queue_2_enq_bits_decodeResult_saturate};
  wire         queue_2_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_2 = {queue_dataIn_hi_lo_lo_hi_hi_2, queue_2_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_4 = {queue_dataIn_hi_lo_lo_hi_2, queue_dataIn_hi_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_crossRead;
  wire         queue_2_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_crossRead, queue_2_enq_bits_decodeResult_crossWrite};
  wire         queue_2_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_2 = {queue_dataIn_hi_lo_hi_lo_hi_2, queue_2_enq_bits_decodeResult_maskUnit};
  wire         queue_2_enq_bits_decodeResult_sReadVD;
  wire         queue_2_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_sReadVD, queue_2_enq_bits_decodeResult_vtype};
  wire         queue_2_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_2 = {queue_dataIn_hi_lo_hi_hi_hi_2, queue_2_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_4 = {queue_dataIn_hi_lo_hi_hi_2, queue_dataIn_hi_lo_hi_lo_2};
  wire [11:0]  queue_dataIn_hi_lo_7 = {queue_dataIn_hi_lo_hi_4, queue_dataIn_hi_lo_lo_4};
  wire         queue_2_enq_bits_decodeResult_reverse;
  wire         queue_2_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_2 = {queue_2_enq_bits_decodeResult_reverse, queue_2_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_2_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_2 = {queue_dataIn_hi_hi_lo_lo_hi_2, queue_2_enq_bits_decodeResult_scheduler};
  wire         queue_2_enq_bits_decodeResult_popCount;
  wire         queue_2_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_popCount, queue_2_enq_bits_decodeResult_ffo};
  wire         queue_2_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_2 = {queue_dataIn_hi_hi_lo_hi_hi_2, queue_2_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_4 = {queue_dataIn_hi_hi_lo_hi_2, queue_dataIn_hi_hi_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_float;
  wire         queue_2_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_float, queue_2_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_2_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_2 = {queue_dataIn_hi_hi_hi_lo_hi_2, queue_2_enq_bits_decodeResult_topUop};
  wire         queue_2_enq_bits_decodeResult_orderReduce;
  wire         queue_2_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_orderReduce, queue_2_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_2_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_2 = {queue_dataIn_hi_hi_hi_hi_hi_2, queue_2_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_4 = {queue_dataIn_hi_hi_hi_hi_2, queue_dataIn_hi_hi_hi_lo_2};
  wire [16:0]  queue_dataIn_hi_hi_7 = {queue_dataIn_hi_hi_hi_4, queue_dataIn_hi_hi_lo_4};
  wire [28:0]  queue_dataIn_hi_7 = {queue_dataIn_hi_hi_7, queue_dataIn_hi_lo_7};
  wire [2:0]   queue_2_enq_bits_segment;
  wire [31:0]  queue_2_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_5 = {queue_2_enq_bits_segment, queue_2_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_5 = {queue_dataIn_lo_lo_hi_5, queue_dataIn_hi_6, queue_dataIn_lo_6};
  wire [1:0]   queue_2_enq_bits_loadStoreEEW;
  wire         queue_2_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_5 = {queue_2_enq_bits_loadStoreEEW, queue_2_enq_bits_mask};
  wire [4:0]   queue_2_enq_bits_vs2;
  wire [4:0]   queue_2_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_5 = {queue_2_enq_bits_vs2, queue_2_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_8 = {queue_dataIn_lo_hi_hi_5, queue_dataIn_lo_hi_lo_5};
  wire [80:0]  queue_dataIn_lo_8 = {queue_dataIn_lo_hi_8, queue_dataIn_lo_lo_5};
  wire         queue_2_enq_bits_lsWholeReg;
  wire [4:0]   queue_2_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_5 = {queue_2_enq_bits_lsWholeReg, queue_2_enq_bits_vs1};
  wire         queue_2_enq_bits_store;
  wire         queue_2_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_5 = {queue_2_enq_bits_store, queue_2_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_8 = {queue_dataIn_hi_lo_hi_5, queue_dataIn_hi_lo_lo_5};
  wire         queue_2_enq_bits_loadStore;
  wire         queue_2_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_5 = {queue_2_enq_bits_loadStore, queue_2_enq_bits_issueInst};
  wire [2:0]   queue_2_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_5 = {queue_2_enq_bits_instructionIndex, queue_dataIn_hi_7, queue_dataIn_lo_7};
  wire [60:0]  queue_dataIn_hi_hi_8 = {queue_dataIn_hi_hi_hi_5, queue_dataIn_hi_hi_lo_5};
  wire [68:0]  queue_dataIn_hi_8 = {queue_dataIn_hi_hi_8, queue_dataIn_hi_lo_8};
  wire [149:0] queue_dataIn_2 = {queue_dataIn_hi_8, queue_dataIn_lo_8};
  wire         queue_dataOut_2_csrInterface_vma = _queue_fifo_2_data_out[0];
  wire         queue_dataOut_2_csrInterface_vta = _queue_fifo_2_data_out[1];
  wire [1:0]   queue_dataOut_2_csrInterface_vxrm = _queue_fifo_2_data_out[3:2];
  wire [1:0]   queue_dataOut_2_csrInterface_vSew = _queue_fifo_2_data_out[5:4];
  wire [2:0]   queue_dataOut_2_csrInterface_vlmul = _queue_fifo_2_data_out[8:6];
  wire [11:0]  queue_dataOut_2_csrInterface_vStart = _queue_fifo_2_data_out[20:9];
  wire [11:0]  queue_dataOut_2_csrInterface_vl = _queue_fifo_2_data_out[32:21];
  wire [31:0]  queue_dataOut_2_readFromScalar = _queue_fifo_2_data_out[64:33];
  wire [2:0]   queue_dataOut_2_segment = _queue_fifo_2_data_out[67:65];
  wire         queue_dataOut_2_mask = _queue_fifo_2_data_out[68];
  wire [1:0]   queue_dataOut_2_loadStoreEEW = _queue_fifo_2_data_out[70:69];
  wire [4:0]   queue_dataOut_2_vd = _queue_fifo_2_data_out[75:71];
  wire [4:0]   queue_dataOut_2_vs2 = _queue_fifo_2_data_out[80:76];
  wire [4:0]   queue_dataOut_2_vs1 = _queue_fifo_2_data_out[85:81];
  wire         queue_dataOut_2_lsWholeReg = _queue_fifo_2_data_out[86];
  wire         queue_dataOut_2_special = _queue_fifo_2_data_out[87];
  wire         queue_dataOut_2_store = _queue_fifo_2_data_out[88];
  wire         queue_dataOut_2_issueInst = _queue_fifo_2_data_out[89];
  wire         queue_dataOut_2_loadStore = _queue_fifo_2_data_out[90];
  wire         queue_dataOut_2_decodeResult_logic = _queue_fifo_2_data_out[91];
  wire         queue_dataOut_2_decodeResult_adder = _queue_fifo_2_data_out[92];
  wire         queue_dataOut_2_decodeResult_shift = _queue_fifo_2_data_out[93];
  wire         queue_dataOut_2_decodeResult_multiplier = _queue_fifo_2_data_out[94];
  wire         queue_dataOut_2_decodeResult_divider = _queue_fifo_2_data_out[95];
  wire         queue_dataOut_2_decodeResult_multiCycle = _queue_fifo_2_data_out[96];
  wire         queue_dataOut_2_decodeResult_other = _queue_fifo_2_data_out[97];
  wire         queue_dataOut_2_decodeResult_unsigned0 = _queue_fifo_2_data_out[98];
  wire         queue_dataOut_2_decodeResult_unsigned1 = _queue_fifo_2_data_out[99];
  wire         queue_dataOut_2_decodeResult_itype = _queue_fifo_2_data_out[100];
  wire         queue_dataOut_2_decodeResult_nr = _queue_fifo_2_data_out[101];
  wire         queue_dataOut_2_decodeResult_red = _queue_fifo_2_data_out[102];
  wire         queue_dataOut_2_decodeResult_widenReduce = _queue_fifo_2_data_out[103];
  wire         queue_dataOut_2_decodeResult_targetRd = _queue_fifo_2_data_out[104];
  wire         queue_dataOut_2_decodeResult_slid = _queue_fifo_2_data_out[105];
  wire         queue_dataOut_2_decodeResult_gather = _queue_fifo_2_data_out[106];
  wire         queue_dataOut_2_decodeResult_gather16 = _queue_fifo_2_data_out[107];
  wire         queue_dataOut_2_decodeResult_compress = _queue_fifo_2_data_out[108];
  wire         queue_dataOut_2_decodeResult_unOrderWrite = _queue_fifo_2_data_out[109];
  wire         queue_dataOut_2_decodeResult_extend = _queue_fifo_2_data_out[110];
  wire         queue_dataOut_2_decodeResult_mv = _queue_fifo_2_data_out[111];
  wire         queue_dataOut_2_decodeResult_iota = _queue_fifo_2_data_out[112];
  wire [3:0]   queue_dataOut_2_decodeResult_uop = _queue_fifo_2_data_out[116:113];
  wire         queue_dataOut_2_decodeResult_maskLogic = _queue_fifo_2_data_out[117];
  wire         queue_dataOut_2_decodeResult_maskDestination = _queue_fifo_2_data_out[118];
  wire         queue_dataOut_2_decodeResult_maskSource = _queue_fifo_2_data_out[119];
  wire         queue_dataOut_2_decodeResult_readOnly = _queue_fifo_2_data_out[120];
  wire         queue_dataOut_2_decodeResult_vwmacc = _queue_fifo_2_data_out[121];
  wire         queue_dataOut_2_decodeResult_saturate = _queue_fifo_2_data_out[122];
  wire         queue_dataOut_2_decodeResult_special = _queue_fifo_2_data_out[123];
  wire         queue_dataOut_2_decodeResult_maskUnit = _queue_fifo_2_data_out[124];
  wire         queue_dataOut_2_decodeResult_crossWrite = _queue_fifo_2_data_out[125];
  wire         queue_dataOut_2_decodeResult_crossRead = _queue_fifo_2_data_out[126];
  wire         queue_dataOut_2_decodeResult_sWrite = _queue_fifo_2_data_out[127];
  wire         queue_dataOut_2_decodeResult_vtype = _queue_fifo_2_data_out[128];
  wire         queue_dataOut_2_decodeResult_sReadVD = _queue_fifo_2_data_out[129];
  wire         queue_dataOut_2_decodeResult_scheduler = _queue_fifo_2_data_out[130];
  wire         queue_dataOut_2_decodeResult_dontNeedExecuteInLane = _queue_fifo_2_data_out[131];
  wire         queue_dataOut_2_decodeResult_reverse = _queue_fifo_2_data_out[132];
  wire         queue_dataOut_2_decodeResult_average = _queue_fifo_2_data_out[133];
  wire         queue_dataOut_2_decodeResult_ffo = _queue_fifo_2_data_out[134];
  wire         queue_dataOut_2_decodeResult_popCount = _queue_fifo_2_data_out[135];
  wire [4:0]   queue_dataOut_2_decodeResult_topUop = _queue_fifo_2_data_out[140:136];
  wire         queue_dataOut_2_decodeResult_specialSlot = _queue_fifo_2_data_out[141];
  wire         queue_dataOut_2_decodeResult_float = _queue_fifo_2_data_out[142];
  wire [1:0]   queue_dataOut_2_decodeResult_fpExecutionType = _queue_fifo_2_data_out[144:143];
  wire         queue_dataOut_2_decodeResult_floatMul = _queue_fifo_2_data_out[145];
  wire         queue_dataOut_2_decodeResult_orderReduce = _queue_fifo_2_data_out[146];
  wire [2:0]   queue_dataOut_2_instructionIndex = _queue_fifo_2_data_out[149:147];
  wire         queue_2_enq_ready = ~_queue_fifo_2_full;
  wire         queue_2_enq_valid;
  assign queue_2_deq_valid = ~_queue_fifo_2_empty | queue_2_enq_valid;
  assign queue_2_deq_bits_instructionIndex = _queue_fifo_2_empty ? queue_2_enq_bits_instructionIndex : queue_dataOut_2_instructionIndex;
  assign queue_2_deq_bits_decodeResult_orderReduce = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_orderReduce : queue_dataOut_2_decodeResult_orderReduce;
  assign queue_2_deq_bits_decodeResult_floatMul = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_floatMul : queue_dataOut_2_decodeResult_floatMul;
  assign queue_2_deq_bits_decodeResult_fpExecutionType = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_fpExecutionType : queue_dataOut_2_decodeResult_fpExecutionType;
  assign queue_2_deq_bits_decodeResult_float = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_float : queue_dataOut_2_decodeResult_float;
  assign queue_2_deq_bits_decodeResult_specialSlot = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_specialSlot : queue_dataOut_2_decodeResult_specialSlot;
  assign queue_2_deq_bits_decodeResult_topUop = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_topUop : queue_dataOut_2_decodeResult_topUop;
  assign queue_2_deq_bits_decodeResult_popCount = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_popCount : queue_dataOut_2_decodeResult_popCount;
  assign queue_2_deq_bits_decodeResult_ffo = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_ffo : queue_dataOut_2_decodeResult_ffo;
  assign queue_2_deq_bits_decodeResult_average = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_average : queue_dataOut_2_decodeResult_average;
  assign queue_2_deq_bits_decodeResult_reverse = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_reverse : queue_dataOut_2_decodeResult_reverse;
  assign queue_2_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_2_decodeResult_dontNeedExecuteInLane;
  assign queue_2_deq_bits_decodeResult_scheduler = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_scheduler : queue_dataOut_2_decodeResult_scheduler;
  assign queue_2_deq_bits_decodeResult_sReadVD = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_sReadVD : queue_dataOut_2_decodeResult_sReadVD;
  assign queue_2_deq_bits_decodeResult_vtype = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_vtype : queue_dataOut_2_decodeResult_vtype;
  assign queue_2_deq_bits_decodeResult_sWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_sWrite : queue_dataOut_2_decodeResult_sWrite;
  assign queue_2_deq_bits_decodeResult_crossRead = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_crossRead : queue_dataOut_2_decodeResult_crossRead;
  assign queue_2_deq_bits_decodeResult_crossWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_crossWrite : queue_dataOut_2_decodeResult_crossWrite;
  assign queue_2_deq_bits_decodeResult_maskUnit = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskUnit : queue_dataOut_2_decodeResult_maskUnit;
  assign queue_2_deq_bits_decodeResult_special = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_special : queue_dataOut_2_decodeResult_special;
  assign queue_2_deq_bits_decodeResult_saturate = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_saturate : queue_dataOut_2_decodeResult_saturate;
  assign queue_2_deq_bits_decodeResult_vwmacc = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_vwmacc : queue_dataOut_2_decodeResult_vwmacc;
  assign queue_2_deq_bits_decodeResult_readOnly = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_readOnly : queue_dataOut_2_decodeResult_readOnly;
  assign queue_2_deq_bits_decodeResult_maskSource = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskSource : queue_dataOut_2_decodeResult_maskSource;
  assign queue_2_deq_bits_decodeResult_maskDestination = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskDestination : queue_dataOut_2_decodeResult_maskDestination;
  assign queue_2_deq_bits_decodeResult_maskLogic = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskLogic : queue_dataOut_2_decodeResult_maskLogic;
  assign queue_2_deq_bits_decodeResult_uop = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_uop : queue_dataOut_2_decodeResult_uop;
  assign queue_2_deq_bits_decodeResult_iota = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_iota : queue_dataOut_2_decodeResult_iota;
  assign queue_2_deq_bits_decodeResult_mv = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_mv : queue_dataOut_2_decodeResult_mv;
  assign queue_2_deq_bits_decodeResult_extend = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_extend : queue_dataOut_2_decodeResult_extend;
  assign queue_2_deq_bits_decodeResult_unOrderWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unOrderWrite : queue_dataOut_2_decodeResult_unOrderWrite;
  assign queue_2_deq_bits_decodeResult_compress = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_compress : queue_dataOut_2_decodeResult_compress;
  assign queue_2_deq_bits_decodeResult_gather16 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_gather16 : queue_dataOut_2_decodeResult_gather16;
  assign queue_2_deq_bits_decodeResult_gather = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_gather : queue_dataOut_2_decodeResult_gather;
  assign queue_2_deq_bits_decodeResult_slid = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_slid : queue_dataOut_2_decodeResult_slid;
  assign queue_2_deq_bits_decodeResult_targetRd = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_targetRd : queue_dataOut_2_decodeResult_targetRd;
  assign queue_2_deq_bits_decodeResult_widenReduce = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_widenReduce : queue_dataOut_2_decodeResult_widenReduce;
  assign queue_2_deq_bits_decodeResult_red = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_red : queue_dataOut_2_decodeResult_red;
  assign queue_2_deq_bits_decodeResult_nr = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_nr : queue_dataOut_2_decodeResult_nr;
  assign queue_2_deq_bits_decodeResult_itype = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_itype : queue_dataOut_2_decodeResult_itype;
  assign queue_2_deq_bits_decodeResult_unsigned1 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unsigned1 : queue_dataOut_2_decodeResult_unsigned1;
  assign queue_2_deq_bits_decodeResult_unsigned0 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unsigned0 : queue_dataOut_2_decodeResult_unsigned0;
  assign queue_2_deq_bits_decodeResult_other = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_other : queue_dataOut_2_decodeResult_other;
  assign queue_2_deq_bits_decodeResult_multiCycle = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_multiCycle : queue_dataOut_2_decodeResult_multiCycle;
  assign queue_2_deq_bits_decodeResult_divider = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_divider : queue_dataOut_2_decodeResult_divider;
  assign queue_2_deq_bits_decodeResult_multiplier = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_multiplier : queue_dataOut_2_decodeResult_multiplier;
  assign queue_2_deq_bits_decodeResult_shift = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_shift : queue_dataOut_2_decodeResult_shift;
  assign queue_2_deq_bits_decodeResult_adder = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_adder : queue_dataOut_2_decodeResult_adder;
  assign queue_2_deq_bits_decodeResult_logic = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_logic : queue_dataOut_2_decodeResult_logic;
  assign queue_2_deq_bits_loadStore = _queue_fifo_2_empty ? queue_2_enq_bits_loadStore : queue_dataOut_2_loadStore;
  assign queue_2_deq_bits_issueInst = _queue_fifo_2_empty ? queue_2_enq_bits_issueInst : queue_dataOut_2_issueInst;
  assign queue_2_deq_bits_store = _queue_fifo_2_empty ? queue_2_enq_bits_store : queue_dataOut_2_store;
  assign queue_2_deq_bits_special = _queue_fifo_2_empty ? queue_2_enq_bits_special : queue_dataOut_2_special;
  assign queue_2_deq_bits_lsWholeReg = _queue_fifo_2_empty ? queue_2_enq_bits_lsWholeReg : queue_dataOut_2_lsWholeReg;
  assign queue_2_deq_bits_vs1 = _queue_fifo_2_empty ? queue_2_enq_bits_vs1 : queue_dataOut_2_vs1;
  assign queue_2_deq_bits_vs2 = _queue_fifo_2_empty ? queue_2_enq_bits_vs2 : queue_dataOut_2_vs2;
  assign queue_2_deq_bits_vd = _queue_fifo_2_empty ? queue_2_enq_bits_vd : queue_dataOut_2_vd;
  assign queue_2_deq_bits_loadStoreEEW = _queue_fifo_2_empty ? queue_2_enq_bits_loadStoreEEW : queue_dataOut_2_loadStoreEEW;
  assign queue_2_deq_bits_mask = _queue_fifo_2_empty ? queue_2_enq_bits_mask : queue_dataOut_2_mask;
  assign queue_2_deq_bits_segment = _queue_fifo_2_empty ? queue_2_enq_bits_segment : queue_dataOut_2_segment;
  assign queue_2_deq_bits_readFromScalar = _queue_fifo_2_empty ? queue_2_enq_bits_readFromScalar : queue_dataOut_2_readFromScalar;
  assign queue_2_deq_bits_csrInterface_vl = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vl : queue_dataOut_2_csrInterface_vl;
  assign queue_2_deq_bits_csrInterface_vStart = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vStart : queue_dataOut_2_csrInterface_vStart;
  assign queue_2_deq_bits_csrInterface_vlmul = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vlmul : queue_dataOut_2_csrInterface_vlmul;
  assign queue_2_deq_bits_csrInterface_vSew = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vSew : queue_dataOut_2_csrInterface_vSew;
  assign queue_2_deq_bits_csrInterface_vxrm = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vxrm : queue_dataOut_2_csrInterface_vxrm;
  assign queue_2_deq_bits_csrInterface_vta = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vta : queue_dataOut_2_csrInterface_vta;
  assign queue_2_deq_bits_csrInterface_vma = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vma : queue_dataOut_2_csrInterface_vma;
  wire         laneVec_2_laneRequest_bits_issueInst = laneRequestSinkWire_2_ready & laneRequestSinkWire_2_valid;
  reg          releasePipe_pipe_v_2;
  wire         releasePipe_pipe_out_2_valid = releasePipe_pipe_v_2;
  wire         laneRequestSourceWire_2_ready;
  wire         validSource_2_valid = laneRequestSourceWire_2_ready & laneRequestSourceWire_2_valid;
  reg  [2:0]   tokenCheck_counter_2;
  wire [2:0]   tokenCheck_counterChange_2 = validSource_2_valid ? 3'h1 : 3'h7;
  assign tokenCheck_2 = ~(tokenCheck_counter_2[2]);
  assign laneRequestSourceWire_2_ready = tokenCheck_2;
  assign queue_2_enq_valid = validSink_2_valid;
  assign queue_2_enq_bits_instructionIndex = validSink_2_bits_instructionIndex;
  assign queue_2_enq_bits_decodeResult_orderReduce = validSink_2_bits_decodeResult_orderReduce;
  assign queue_2_enq_bits_decodeResult_floatMul = validSink_2_bits_decodeResult_floatMul;
  assign queue_2_enq_bits_decodeResult_fpExecutionType = validSink_2_bits_decodeResult_fpExecutionType;
  assign queue_2_enq_bits_decodeResult_float = validSink_2_bits_decodeResult_float;
  assign queue_2_enq_bits_decodeResult_specialSlot = validSink_2_bits_decodeResult_specialSlot;
  assign queue_2_enq_bits_decodeResult_topUop = validSink_2_bits_decodeResult_topUop;
  assign queue_2_enq_bits_decodeResult_popCount = validSink_2_bits_decodeResult_popCount;
  assign queue_2_enq_bits_decodeResult_ffo = validSink_2_bits_decodeResult_ffo;
  assign queue_2_enq_bits_decodeResult_average = validSink_2_bits_decodeResult_average;
  assign queue_2_enq_bits_decodeResult_reverse = validSink_2_bits_decodeResult_reverse;
  assign queue_2_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_2_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_2_enq_bits_decodeResult_scheduler = validSink_2_bits_decodeResult_scheduler;
  assign queue_2_enq_bits_decodeResult_sReadVD = validSink_2_bits_decodeResult_sReadVD;
  assign queue_2_enq_bits_decodeResult_vtype = validSink_2_bits_decodeResult_vtype;
  assign queue_2_enq_bits_decodeResult_sWrite = validSink_2_bits_decodeResult_sWrite;
  assign queue_2_enq_bits_decodeResult_crossRead = validSink_2_bits_decodeResult_crossRead;
  assign queue_2_enq_bits_decodeResult_crossWrite = validSink_2_bits_decodeResult_crossWrite;
  assign queue_2_enq_bits_decodeResult_maskUnit = validSink_2_bits_decodeResult_maskUnit;
  assign queue_2_enq_bits_decodeResult_special = validSink_2_bits_decodeResult_special;
  assign queue_2_enq_bits_decodeResult_saturate = validSink_2_bits_decodeResult_saturate;
  assign queue_2_enq_bits_decodeResult_vwmacc = validSink_2_bits_decodeResult_vwmacc;
  assign queue_2_enq_bits_decodeResult_readOnly = validSink_2_bits_decodeResult_readOnly;
  assign queue_2_enq_bits_decodeResult_maskSource = validSink_2_bits_decodeResult_maskSource;
  assign queue_2_enq_bits_decodeResult_maskDestination = validSink_2_bits_decodeResult_maskDestination;
  assign queue_2_enq_bits_decodeResult_maskLogic = validSink_2_bits_decodeResult_maskLogic;
  assign queue_2_enq_bits_decodeResult_uop = validSink_2_bits_decodeResult_uop;
  assign queue_2_enq_bits_decodeResult_iota = validSink_2_bits_decodeResult_iota;
  assign queue_2_enq_bits_decodeResult_mv = validSink_2_bits_decodeResult_mv;
  assign queue_2_enq_bits_decodeResult_extend = validSink_2_bits_decodeResult_extend;
  assign queue_2_enq_bits_decodeResult_unOrderWrite = validSink_2_bits_decodeResult_unOrderWrite;
  assign queue_2_enq_bits_decodeResult_compress = validSink_2_bits_decodeResult_compress;
  assign queue_2_enq_bits_decodeResult_gather16 = validSink_2_bits_decodeResult_gather16;
  assign queue_2_enq_bits_decodeResult_gather = validSink_2_bits_decodeResult_gather;
  assign queue_2_enq_bits_decodeResult_slid = validSink_2_bits_decodeResult_slid;
  assign queue_2_enq_bits_decodeResult_targetRd = validSink_2_bits_decodeResult_targetRd;
  assign queue_2_enq_bits_decodeResult_widenReduce = validSink_2_bits_decodeResult_widenReduce;
  assign queue_2_enq_bits_decodeResult_red = validSink_2_bits_decodeResult_red;
  assign queue_2_enq_bits_decodeResult_nr = validSink_2_bits_decodeResult_nr;
  assign queue_2_enq_bits_decodeResult_itype = validSink_2_bits_decodeResult_itype;
  assign queue_2_enq_bits_decodeResult_unsigned1 = validSink_2_bits_decodeResult_unsigned1;
  assign queue_2_enq_bits_decodeResult_unsigned0 = validSink_2_bits_decodeResult_unsigned0;
  assign queue_2_enq_bits_decodeResult_other = validSink_2_bits_decodeResult_other;
  assign queue_2_enq_bits_decodeResult_multiCycle = validSink_2_bits_decodeResult_multiCycle;
  assign queue_2_enq_bits_decodeResult_divider = validSink_2_bits_decodeResult_divider;
  assign queue_2_enq_bits_decodeResult_multiplier = validSink_2_bits_decodeResult_multiplier;
  assign queue_2_enq_bits_decodeResult_shift = validSink_2_bits_decodeResult_shift;
  assign queue_2_enq_bits_decodeResult_adder = validSink_2_bits_decodeResult_adder;
  assign queue_2_enq_bits_decodeResult_logic = validSink_2_bits_decodeResult_logic;
  assign queue_2_enq_bits_loadStore = validSink_2_bits_loadStore;
  assign queue_2_enq_bits_issueInst = validSink_2_bits_issueInst;
  assign queue_2_enq_bits_store = validSink_2_bits_store;
  assign queue_2_enq_bits_special = validSink_2_bits_special;
  assign queue_2_enq_bits_lsWholeReg = validSink_2_bits_lsWholeReg;
  assign queue_2_enq_bits_vs1 = validSink_2_bits_vs1;
  assign queue_2_enq_bits_vs2 = validSink_2_bits_vs2;
  assign queue_2_enq_bits_vd = validSink_2_bits_vd;
  assign queue_2_enq_bits_loadStoreEEW = validSink_2_bits_loadStoreEEW;
  assign queue_2_enq_bits_mask = validSink_2_bits_mask;
  assign queue_2_enq_bits_segment = validSink_2_bits_segment;
  assign queue_2_enq_bits_readFromScalar = validSink_2_bits_readFromScalar;
  assign queue_2_enq_bits_csrInterface_vl = validSink_2_bits_csrInterface_vl;
  assign queue_2_enq_bits_csrInterface_vStart = validSink_2_bits_csrInterface_vStart;
  assign queue_2_enq_bits_csrInterface_vlmul = validSink_2_bits_csrInterface_vlmul;
  assign queue_2_enq_bits_csrInterface_vSew = validSink_2_bits_csrInterface_vSew;
  assign queue_2_enq_bits_csrInterface_vxrm = validSink_2_bits_csrInterface_vxrm;
  assign queue_2_enq_bits_csrInterface_vta = validSink_2_bits_csrInterface_vta;
  assign queue_2_enq_bits_csrInterface_vma = validSink_2_bits_csrInterface_vma;
  reg          shifterReg_2_0_valid;
  assign validSink_2_valid = shifterReg_2_0_valid;
  reg  [2:0]   shifterReg_2_0_bits_instructionIndex;
  assign validSink_2_bits_instructionIndex = shifterReg_2_0_bits_instructionIndex;
  reg          shifterReg_2_0_bits_decodeResult_orderReduce;
  assign validSink_2_bits_decodeResult_orderReduce = shifterReg_2_0_bits_decodeResult_orderReduce;
  reg          shifterReg_2_0_bits_decodeResult_floatMul;
  assign validSink_2_bits_decodeResult_floatMul = shifterReg_2_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_2_0_bits_decodeResult_fpExecutionType;
  assign validSink_2_bits_decodeResult_fpExecutionType = shifterReg_2_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_2_0_bits_decodeResult_float;
  assign validSink_2_bits_decodeResult_float = shifterReg_2_0_bits_decodeResult_float;
  reg          shifterReg_2_0_bits_decodeResult_specialSlot;
  assign validSink_2_bits_decodeResult_specialSlot = shifterReg_2_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_2_0_bits_decodeResult_topUop;
  assign validSink_2_bits_decodeResult_topUop = shifterReg_2_0_bits_decodeResult_topUop;
  reg          shifterReg_2_0_bits_decodeResult_popCount;
  assign validSink_2_bits_decodeResult_popCount = shifterReg_2_0_bits_decodeResult_popCount;
  reg          shifterReg_2_0_bits_decodeResult_ffo;
  assign validSink_2_bits_decodeResult_ffo = shifterReg_2_0_bits_decodeResult_ffo;
  reg          shifterReg_2_0_bits_decodeResult_average;
  assign validSink_2_bits_decodeResult_average = shifterReg_2_0_bits_decodeResult_average;
  reg          shifterReg_2_0_bits_decodeResult_reverse;
  assign validSink_2_bits_decodeResult_reverse = shifterReg_2_0_bits_decodeResult_reverse;
  reg          shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_2_bits_decodeResult_dontNeedExecuteInLane = shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_2_0_bits_decodeResult_scheduler;
  assign validSink_2_bits_decodeResult_scheduler = shifterReg_2_0_bits_decodeResult_scheduler;
  reg          shifterReg_2_0_bits_decodeResult_sReadVD;
  assign validSink_2_bits_decodeResult_sReadVD = shifterReg_2_0_bits_decodeResult_sReadVD;
  reg          shifterReg_2_0_bits_decodeResult_vtype;
  assign validSink_2_bits_decodeResult_vtype = shifterReg_2_0_bits_decodeResult_vtype;
  reg          shifterReg_2_0_bits_decodeResult_sWrite;
  assign validSink_2_bits_decodeResult_sWrite = shifterReg_2_0_bits_decodeResult_sWrite;
  reg          shifterReg_2_0_bits_decodeResult_crossRead;
  assign validSink_2_bits_decodeResult_crossRead = shifterReg_2_0_bits_decodeResult_crossRead;
  reg          shifterReg_2_0_bits_decodeResult_crossWrite;
  assign validSink_2_bits_decodeResult_crossWrite = shifterReg_2_0_bits_decodeResult_crossWrite;
  reg          shifterReg_2_0_bits_decodeResult_maskUnit;
  assign validSink_2_bits_decodeResult_maskUnit = shifterReg_2_0_bits_decodeResult_maskUnit;
  reg          shifterReg_2_0_bits_decodeResult_special;
  assign validSink_2_bits_decodeResult_special = shifterReg_2_0_bits_decodeResult_special;
  reg          shifterReg_2_0_bits_decodeResult_saturate;
  assign validSink_2_bits_decodeResult_saturate = shifterReg_2_0_bits_decodeResult_saturate;
  reg          shifterReg_2_0_bits_decodeResult_vwmacc;
  assign validSink_2_bits_decodeResult_vwmacc = shifterReg_2_0_bits_decodeResult_vwmacc;
  reg          shifterReg_2_0_bits_decodeResult_readOnly;
  assign validSink_2_bits_decodeResult_readOnly = shifterReg_2_0_bits_decodeResult_readOnly;
  reg          shifterReg_2_0_bits_decodeResult_maskSource;
  assign validSink_2_bits_decodeResult_maskSource = shifterReg_2_0_bits_decodeResult_maskSource;
  reg          shifterReg_2_0_bits_decodeResult_maskDestination;
  assign validSink_2_bits_decodeResult_maskDestination = shifterReg_2_0_bits_decodeResult_maskDestination;
  reg          shifterReg_2_0_bits_decodeResult_maskLogic;
  assign validSink_2_bits_decodeResult_maskLogic = shifterReg_2_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_2_0_bits_decodeResult_uop;
  assign validSink_2_bits_decodeResult_uop = shifterReg_2_0_bits_decodeResult_uop;
  reg          shifterReg_2_0_bits_decodeResult_iota;
  assign validSink_2_bits_decodeResult_iota = shifterReg_2_0_bits_decodeResult_iota;
  reg          shifterReg_2_0_bits_decodeResult_mv;
  assign validSink_2_bits_decodeResult_mv = shifterReg_2_0_bits_decodeResult_mv;
  reg          shifterReg_2_0_bits_decodeResult_extend;
  assign validSink_2_bits_decodeResult_extend = shifterReg_2_0_bits_decodeResult_extend;
  reg          shifterReg_2_0_bits_decodeResult_unOrderWrite;
  assign validSink_2_bits_decodeResult_unOrderWrite = shifterReg_2_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_2_0_bits_decodeResult_compress;
  assign validSink_2_bits_decodeResult_compress = shifterReg_2_0_bits_decodeResult_compress;
  reg          shifterReg_2_0_bits_decodeResult_gather16;
  assign validSink_2_bits_decodeResult_gather16 = shifterReg_2_0_bits_decodeResult_gather16;
  reg          shifterReg_2_0_bits_decodeResult_gather;
  assign validSink_2_bits_decodeResult_gather = shifterReg_2_0_bits_decodeResult_gather;
  reg          shifterReg_2_0_bits_decodeResult_slid;
  assign validSink_2_bits_decodeResult_slid = shifterReg_2_0_bits_decodeResult_slid;
  reg          shifterReg_2_0_bits_decodeResult_targetRd;
  assign validSink_2_bits_decodeResult_targetRd = shifterReg_2_0_bits_decodeResult_targetRd;
  reg          shifterReg_2_0_bits_decodeResult_widenReduce;
  assign validSink_2_bits_decodeResult_widenReduce = shifterReg_2_0_bits_decodeResult_widenReduce;
  reg          shifterReg_2_0_bits_decodeResult_red;
  assign validSink_2_bits_decodeResult_red = shifterReg_2_0_bits_decodeResult_red;
  reg          shifterReg_2_0_bits_decodeResult_nr;
  assign validSink_2_bits_decodeResult_nr = shifterReg_2_0_bits_decodeResult_nr;
  reg          shifterReg_2_0_bits_decodeResult_itype;
  assign validSink_2_bits_decodeResult_itype = shifterReg_2_0_bits_decodeResult_itype;
  reg          shifterReg_2_0_bits_decodeResult_unsigned1;
  assign validSink_2_bits_decodeResult_unsigned1 = shifterReg_2_0_bits_decodeResult_unsigned1;
  reg          shifterReg_2_0_bits_decodeResult_unsigned0;
  assign validSink_2_bits_decodeResult_unsigned0 = shifterReg_2_0_bits_decodeResult_unsigned0;
  reg          shifterReg_2_0_bits_decodeResult_other;
  assign validSink_2_bits_decodeResult_other = shifterReg_2_0_bits_decodeResult_other;
  reg          shifterReg_2_0_bits_decodeResult_multiCycle;
  assign validSink_2_bits_decodeResult_multiCycle = shifterReg_2_0_bits_decodeResult_multiCycle;
  reg          shifterReg_2_0_bits_decodeResult_divider;
  assign validSink_2_bits_decodeResult_divider = shifterReg_2_0_bits_decodeResult_divider;
  reg          shifterReg_2_0_bits_decodeResult_multiplier;
  assign validSink_2_bits_decodeResult_multiplier = shifterReg_2_0_bits_decodeResult_multiplier;
  reg          shifterReg_2_0_bits_decodeResult_shift;
  assign validSink_2_bits_decodeResult_shift = shifterReg_2_0_bits_decodeResult_shift;
  reg          shifterReg_2_0_bits_decodeResult_adder;
  assign validSink_2_bits_decodeResult_adder = shifterReg_2_0_bits_decodeResult_adder;
  reg          shifterReg_2_0_bits_decodeResult_logic;
  assign validSink_2_bits_decodeResult_logic = shifterReg_2_0_bits_decodeResult_logic;
  reg          shifterReg_2_0_bits_loadStore;
  assign validSink_2_bits_loadStore = shifterReg_2_0_bits_loadStore;
  reg          shifterReg_2_0_bits_issueInst;
  assign validSink_2_bits_issueInst = shifterReg_2_0_bits_issueInst;
  reg          shifterReg_2_0_bits_store;
  assign validSink_2_bits_store = shifterReg_2_0_bits_store;
  reg          shifterReg_2_0_bits_special;
  assign validSink_2_bits_special = shifterReg_2_0_bits_special;
  reg          shifterReg_2_0_bits_lsWholeReg;
  assign validSink_2_bits_lsWholeReg = shifterReg_2_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_2_0_bits_vs1;
  assign validSink_2_bits_vs1 = shifterReg_2_0_bits_vs1;
  reg  [4:0]   shifterReg_2_0_bits_vs2;
  assign validSink_2_bits_vs2 = shifterReg_2_0_bits_vs2;
  reg  [4:0]   shifterReg_2_0_bits_vd;
  assign validSink_2_bits_vd = shifterReg_2_0_bits_vd;
  reg  [1:0]   shifterReg_2_0_bits_loadStoreEEW;
  assign validSink_2_bits_loadStoreEEW = shifterReg_2_0_bits_loadStoreEEW;
  reg          shifterReg_2_0_bits_mask;
  assign validSink_2_bits_mask = shifterReg_2_0_bits_mask;
  reg  [2:0]   shifterReg_2_0_bits_segment;
  assign validSink_2_bits_segment = shifterReg_2_0_bits_segment;
  reg  [31:0]  shifterReg_2_0_bits_readFromScalar;
  assign validSink_2_bits_readFromScalar = shifterReg_2_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_2_0_bits_csrInterface_vl;
  assign validSink_2_bits_csrInterface_vl = shifterReg_2_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_2_0_bits_csrInterface_vStart;
  assign validSink_2_bits_csrInterface_vStart = shifterReg_2_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_2_0_bits_csrInterface_vlmul;
  assign validSink_2_bits_csrInterface_vlmul = shifterReg_2_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_2_0_bits_csrInterface_vSew;
  assign validSink_2_bits_csrInterface_vSew = shifterReg_2_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_2_0_bits_csrInterface_vxrm;
  assign validSink_2_bits_csrInterface_vxrm = shifterReg_2_0_bits_csrInterface_vxrm;
  reg          shifterReg_2_0_bits_csrInterface_vta;
  assign validSink_2_bits_csrInterface_vta = shifterReg_2_0_bits_csrInterface_vta;
  reg          shifterReg_2_0_bits_csrInterface_vma;
  assign validSink_2_bits_csrInterface_vma = shifterReg_2_0_bits_csrInterface_vma;
  wire         shifterValid_2 = shifterReg_2_0_valid | validSource_2_valid;
  wire         validSink_3_valid;
  wire [2:0]   validSink_3_bits_instructionIndex;
  wire         validSink_3_bits_decodeResult_orderReduce;
  wire         validSink_3_bits_decodeResult_floatMul;
  wire [1:0]   validSink_3_bits_decodeResult_fpExecutionType;
  wire         validSink_3_bits_decodeResult_float;
  wire         validSink_3_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_3_bits_decodeResult_topUop;
  wire         validSink_3_bits_decodeResult_popCount;
  wire         validSink_3_bits_decodeResult_ffo;
  wire         validSink_3_bits_decodeResult_average;
  wire         validSink_3_bits_decodeResult_reverse;
  wire         validSink_3_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_3_bits_decodeResult_scheduler;
  wire         validSink_3_bits_decodeResult_sReadVD;
  wire         validSink_3_bits_decodeResult_vtype;
  wire         validSink_3_bits_decodeResult_sWrite;
  wire         validSink_3_bits_decodeResult_crossRead;
  wire         validSink_3_bits_decodeResult_crossWrite;
  wire         validSink_3_bits_decodeResult_maskUnit;
  wire         validSink_3_bits_decodeResult_special;
  wire         validSink_3_bits_decodeResult_saturate;
  wire         validSink_3_bits_decodeResult_vwmacc;
  wire         validSink_3_bits_decodeResult_readOnly;
  wire         validSink_3_bits_decodeResult_maskSource;
  wire         validSink_3_bits_decodeResult_maskDestination;
  wire         validSink_3_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_3_bits_decodeResult_uop;
  wire         validSink_3_bits_decodeResult_iota;
  wire         validSink_3_bits_decodeResult_mv;
  wire         validSink_3_bits_decodeResult_extend;
  wire         validSink_3_bits_decodeResult_unOrderWrite;
  wire         validSink_3_bits_decodeResult_compress;
  wire         validSink_3_bits_decodeResult_gather16;
  wire         validSink_3_bits_decodeResult_gather;
  wire         validSink_3_bits_decodeResult_slid;
  wire         validSink_3_bits_decodeResult_targetRd;
  wire         validSink_3_bits_decodeResult_widenReduce;
  wire         validSink_3_bits_decodeResult_red;
  wire         validSink_3_bits_decodeResult_nr;
  wire         validSink_3_bits_decodeResult_itype;
  wire         validSink_3_bits_decodeResult_unsigned1;
  wire         validSink_3_bits_decodeResult_unsigned0;
  wire         validSink_3_bits_decodeResult_other;
  wire         validSink_3_bits_decodeResult_multiCycle;
  wire         validSink_3_bits_decodeResult_divider;
  wire         validSink_3_bits_decodeResult_multiplier;
  wire         validSink_3_bits_decodeResult_shift;
  wire         validSink_3_bits_decodeResult_adder;
  wire         validSink_3_bits_decodeResult_logic;
  wire         validSink_3_bits_loadStore;
  wire         validSink_3_bits_issueInst;
  wire         validSink_3_bits_store;
  wire         validSink_3_bits_special;
  wire         validSink_3_bits_lsWholeReg;
  wire [4:0]   validSink_3_bits_vs1;
  wire [4:0]   validSink_3_bits_vs2;
  wire [4:0]   validSink_3_bits_vd;
  wire [1:0]   validSink_3_bits_loadStoreEEW;
  wire         validSink_3_bits_mask;
  wire [2:0]   validSink_3_bits_segment;
  wire [31:0]  validSink_3_bits_readFromScalar;
  wire [11:0]  validSink_3_bits_csrInterface_vl;
  wire [11:0]  validSink_3_bits_csrInterface_vStart;
  wire [2:0]   validSink_3_bits_csrInterface_vlmul;
  wire [1:0]   validSink_3_bits_csrInterface_vSew;
  wire [1:0]   validSink_3_bits_csrInterface_vxrm;
  wire         validSink_3_bits_csrInterface_vta;
  wire         validSink_3_bits_csrInterface_vma;
  wire         laneRequestSinkWire_3_valid = queue_3_deq_valid;
  wire [2:0]   laneRequestSinkWire_3_bits_instructionIndex = queue_3_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_3_bits_decodeResult_orderReduce = queue_3_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_3_bits_decodeResult_floatMul = queue_3_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_3_bits_decodeResult_fpExecutionType = queue_3_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_3_bits_decodeResult_float = queue_3_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_3_bits_decodeResult_specialSlot = queue_3_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_3_bits_decodeResult_topUop = queue_3_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_3_bits_decodeResult_popCount = queue_3_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_3_bits_decodeResult_ffo = queue_3_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_3_bits_decodeResult_average = queue_3_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_3_bits_decodeResult_reverse = queue_3_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_3_bits_decodeResult_dontNeedExecuteInLane = queue_3_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_3_bits_decodeResult_scheduler = queue_3_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_3_bits_decodeResult_sReadVD = queue_3_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_3_bits_decodeResult_vtype = queue_3_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_3_bits_decodeResult_sWrite = queue_3_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_crossRead = queue_3_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_3_bits_decodeResult_crossWrite = queue_3_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskUnit = queue_3_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_3_bits_decodeResult_special = queue_3_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_3_bits_decodeResult_saturate = queue_3_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_3_bits_decodeResult_vwmacc = queue_3_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_3_bits_decodeResult_readOnly = queue_3_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskSource = queue_3_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskDestination = queue_3_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskLogic = queue_3_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_3_bits_decodeResult_uop = queue_3_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_3_bits_decodeResult_iota = queue_3_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_3_bits_decodeResult_mv = queue_3_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_3_bits_decodeResult_extend = queue_3_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_3_bits_decodeResult_unOrderWrite = queue_3_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_compress = queue_3_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_3_bits_decodeResult_gather16 = queue_3_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_3_bits_decodeResult_gather = queue_3_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_3_bits_decodeResult_slid = queue_3_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_3_bits_decodeResult_targetRd = queue_3_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_3_bits_decodeResult_widenReduce = queue_3_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_3_bits_decodeResult_red = queue_3_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_3_bits_decodeResult_nr = queue_3_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_3_bits_decodeResult_itype = queue_3_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_3_bits_decodeResult_unsigned1 = queue_3_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_3_bits_decodeResult_unsigned0 = queue_3_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_3_bits_decodeResult_other = queue_3_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_3_bits_decodeResult_multiCycle = queue_3_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_3_bits_decodeResult_divider = queue_3_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_3_bits_decodeResult_multiplier = queue_3_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_3_bits_decodeResult_shift = queue_3_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_3_bits_decodeResult_adder = queue_3_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_3_bits_decodeResult_logic = queue_3_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_3_bits_loadStore = queue_3_deq_bits_loadStore;
  wire         laneRequestSinkWire_3_bits_issueInst = queue_3_deq_bits_issueInst;
  wire         laneRequestSinkWire_3_bits_store = queue_3_deq_bits_store;
  wire         laneRequestSinkWire_3_bits_special = queue_3_deq_bits_special;
  wire         laneRequestSinkWire_3_bits_lsWholeReg = queue_3_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_3_bits_vs1 = queue_3_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_3_bits_vs2 = queue_3_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_3_bits_vd = queue_3_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_3_bits_loadStoreEEW = queue_3_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_3_bits_mask = queue_3_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_3_bits_segment = queue_3_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_3_bits_readFromScalar = queue_3_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_3_bits_csrInterface_vl = queue_3_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_3_bits_csrInterface_vStart = queue_3_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_3_bits_csrInterface_vlmul = queue_3_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_3_bits_csrInterface_vSew = queue_3_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_3_bits_csrInterface_vxrm = queue_3_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_3_bits_csrInterface_vta = queue_3_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_3_bits_csrInterface_vma = queue_3_deq_bits_csrInterface_vma;
  wire [1:0]   queue_3_enq_bits_csrInterface_vxrm;
  wire         queue_3_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_9 = {queue_3_enq_bits_csrInterface_vxrm, queue_3_enq_bits_csrInterface_vta};
  wire         queue_3_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_9 = {queue_dataIn_lo_hi_9, queue_3_enq_bits_csrInterface_vma};
  wire [2:0]   queue_3_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_3_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_9 = {queue_3_enq_bits_csrInterface_vlmul, queue_3_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_3_enq_bits_csrInterface_vl;
  wire [11:0]  queue_3_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_9 = {queue_3_enq_bits_csrInterface_vl, queue_3_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_9 = {queue_dataIn_hi_hi_9, queue_dataIn_hi_lo_9};
  wire         queue_3_enq_bits_decodeResult_shift;
  wire         queue_3_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_3 = {queue_3_enq_bits_decodeResult_shift, queue_3_enq_bits_decodeResult_adder};
  wire         queue_3_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_3 = {queue_dataIn_lo_lo_lo_lo_hi_3, queue_3_enq_bits_decodeResult_logic};
  wire         queue_3_enq_bits_decodeResult_multiCycle;
  wire         queue_3_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_multiCycle, queue_3_enq_bits_decodeResult_divider};
  wire         queue_3_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_3 = {queue_dataIn_lo_lo_lo_hi_hi_3, queue_3_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_3 = {queue_dataIn_lo_lo_lo_hi_3, queue_dataIn_lo_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_unsigned1;
  wire         queue_3_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_unsigned1, queue_3_enq_bits_decodeResult_unsigned0};
  wire         queue_3_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_3 = {queue_dataIn_lo_lo_hi_lo_hi_3, queue_3_enq_bits_decodeResult_other};
  wire         queue_3_enq_bits_decodeResult_red;
  wire         queue_3_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_red, queue_3_enq_bits_decodeResult_nr};
  wire         queue_3_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_3 = {queue_dataIn_lo_lo_hi_hi_hi_3, queue_3_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_6 = {queue_dataIn_lo_lo_hi_hi_3, queue_dataIn_lo_lo_hi_lo_3};
  wire [11:0]  queue_dataIn_lo_lo_6 = {queue_dataIn_lo_lo_hi_6, queue_dataIn_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_slid;
  wire         queue_3_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_3 = {queue_3_enq_bits_decodeResult_slid, queue_3_enq_bits_decodeResult_targetRd};
  wire         queue_3_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_3 = {queue_dataIn_lo_hi_lo_lo_hi_3, queue_3_enq_bits_decodeResult_widenReduce};
  wire         queue_3_enq_bits_decodeResult_compress;
  wire         queue_3_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_compress, queue_3_enq_bits_decodeResult_gather16};
  wire         queue_3_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_3 = {queue_dataIn_lo_hi_lo_hi_hi_3, queue_3_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_6 = {queue_dataIn_lo_hi_lo_hi_3, queue_dataIn_lo_hi_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_mv;
  wire         queue_3_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_mv, queue_3_enq_bits_decodeResult_extend};
  wire         queue_3_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_3 = {queue_dataIn_lo_hi_hi_lo_hi_3, queue_3_enq_bits_decodeResult_unOrderWrite};
  wire         queue_3_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_3_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_maskLogic, queue_3_enq_bits_decodeResult_uop};
  wire         queue_3_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_3 = {queue_dataIn_lo_hi_hi_hi_hi_3, queue_3_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_6 = {queue_dataIn_lo_hi_hi_hi_3, queue_dataIn_lo_hi_hi_lo_3};
  wire [14:0]  queue_dataIn_lo_hi_10 = {queue_dataIn_lo_hi_hi_6, queue_dataIn_lo_hi_lo_6};
  wire [26:0]  queue_dataIn_lo_10 = {queue_dataIn_lo_hi_10, queue_dataIn_lo_lo_6};
  wire         queue_3_enq_bits_decodeResult_readOnly;
  wire         queue_3_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_3 = {queue_3_enq_bits_decodeResult_readOnly, queue_3_enq_bits_decodeResult_maskSource};
  wire         queue_3_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_3 = {queue_dataIn_hi_lo_lo_lo_hi_3, queue_3_enq_bits_decodeResult_maskDestination};
  wire         queue_3_enq_bits_decodeResult_special;
  wire         queue_3_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_special, queue_3_enq_bits_decodeResult_saturate};
  wire         queue_3_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_3 = {queue_dataIn_hi_lo_lo_hi_hi_3, queue_3_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_6 = {queue_dataIn_hi_lo_lo_hi_3, queue_dataIn_hi_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_crossRead;
  wire         queue_3_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_crossRead, queue_3_enq_bits_decodeResult_crossWrite};
  wire         queue_3_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_3 = {queue_dataIn_hi_lo_hi_lo_hi_3, queue_3_enq_bits_decodeResult_maskUnit};
  wire         queue_3_enq_bits_decodeResult_sReadVD;
  wire         queue_3_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_sReadVD, queue_3_enq_bits_decodeResult_vtype};
  wire         queue_3_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_3 = {queue_dataIn_hi_lo_hi_hi_hi_3, queue_3_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_6 = {queue_dataIn_hi_lo_hi_hi_3, queue_dataIn_hi_lo_hi_lo_3};
  wire [11:0]  queue_dataIn_hi_lo_10 = {queue_dataIn_hi_lo_hi_6, queue_dataIn_hi_lo_lo_6};
  wire         queue_3_enq_bits_decodeResult_reverse;
  wire         queue_3_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_3 = {queue_3_enq_bits_decodeResult_reverse, queue_3_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_3_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_3 = {queue_dataIn_hi_hi_lo_lo_hi_3, queue_3_enq_bits_decodeResult_scheduler};
  wire         queue_3_enq_bits_decodeResult_popCount;
  wire         queue_3_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_popCount, queue_3_enq_bits_decodeResult_ffo};
  wire         queue_3_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_3 = {queue_dataIn_hi_hi_lo_hi_hi_3, queue_3_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_6 = {queue_dataIn_hi_hi_lo_hi_3, queue_dataIn_hi_hi_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_float;
  wire         queue_3_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_float, queue_3_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_3_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_3 = {queue_dataIn_hi_hi_hi_lo_hi_3, queue_3_enq_bits_decodeResult_topUop};
  wire         queue_3_enq_bits_decodeResult_orderReduce;
  wire         queue_3_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_orderReduce, queue_3_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_3_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_3 = {queue_dataIn_hi_hi_hi_hi_hi_3, queue_3_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_6 = {queue_dataIn_hi_hi_hi_hi_3, queue_dataIn_hi_hi_hi_lo_3};
  wire [16:0]  queue_dataIn_hi_hi_10 = {queue_dataIn_hi_hi_hi_6, queue_dataIn_hi_hi_lo_6};
  wire [28:0]  queue_dataIn_hi_10 = {queue_dataIn_hi_hi_10, queue_dataIn_hi_lo_10};
  wire [2:0]   queue_3_enq_bits_segment;
  wire [31:0]  queue_3_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_7 = {queue_3_enq_bits_segment, queue_3_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_7 = {queue_dataIn_lo_lo_hi_7, queue_dataIn_hi_9, queue_dataIn_lo_9};
  wire [1:0]   queue_3_enq_bits_loadStoreEEW;
  wire         queue_3_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_7 = {queue_3_enq_bits_loadStoreEEW, queue_3_enq_bits_mask};
  wire [4:0]   queue_3_enq_bits_vs2;
  wire [4:0]   queue_3_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_7 = {queue_3_enq_bits_vs2, queue_3_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_11 = {queue_dataIn_lo_hi_hi_7, queue_dataIn_lo_hi_lo_7};
  wire [80:0]  queue_dataIn_lo_11 = {queue_dataIn_lo_hi_11, queue_dataIn_lo_lo_7};
  wire         queue_3_enq_bits_lsWholeReg;
  wire [4:0]   queue_3_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_7 = {queue_3_enq_bits_lsWholeReg, queue_3_enq_bits_vs1};
  wire         queue_3_enq_bits_store;
  wire         queue_3_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_7 = {queue_3_enq_bits_store, queue_3_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_11 = {queue_dataIn_hi_lo_hi_7, queue_dataIn_hi_lo_lo_7};
  wire         queue_3_enq_bits_loadStore;
  wire         queue_3_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_7 = {queue_3_enq_bits_loadStore, queue_3_enq_bits_issueInst};
  wire [2:0]   queue_3_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_7 = {queue_3_enq_bits_instructionIndex, queue_dataIn_hi_10, queue_dataIn_lo_10};
  wire [60:0]  queue_dataIn_hi_hi_11 = {queue_dataIn_hi_hi_hi_7, queue_dataIn_hi_hi_lo_7};
  wire [68:0]  queue_dataIn_hi_11 = {queue_dataIn_hi_hi_11, queue_dataIn_hi_lo_11};
  wire [149:0] queue_dataIn_3 = {queue_dataIn_hi_11, queue_dataIn_lo_11};
  wire         queue_dataOut_3_csrInterface_vma = _queue_fifo_3_data_out[0];
  wire         queue_dataOut_3_csrInterface_vta = _queue_fifo_3_data_out[1];
  wire [1:0]   queue_dataOut_3_csrInterface_vxrm = _queue_fifo_3_data_out[3:2];
  wire [1:0]   queue_dataOut_3_csrInterface_vSew = _queue_fifo_3_data_out[5:4];
  wire [2:0]   queue_dataOut_3_csrInterface_vlmul = _queue_fifo_3_data_out[8:6];
  wire [11:0]  queue_dataOut_3_csrInterface_vStart = _queue_fifo_3_data_out[20:9];
  wire [11:0]  queue_dataOut_3_csrInterface_vl = _queue_fifo_3_data_out[32:21];
  wire [31:0]  queue_dataOut_3_readFromScalar = _queue_fifo_3_data_out[64:33];
  wire [2:0]   queue_dataOut_3_segment = _queue_fifo_3_data_out[67:65];
  wire         queue_dataOut_3_mask = _queue_fifo_3_data_out[68];
  wire [1:0]   queue_dataOut_3_loadStoreEEW = _queue_fifo_3_data_out[70:69];
  wire [4:0]   queue_dataOut_3_vd = _queue_fifo_3_data_out[75:71];
  wire [4:0]   queue_dataOut_3_vs2 = _queue_fifo_3_data_out[80:76];
  wire [4:0]   queue_dataOut_3_vs1 = _queue_fifo_3_data_out[85:81];
  wire         queue_dataOut_3_lsWholeReg = _queue_fifo_3_data_out[86];
  wire         queue_dataOut_3_special = _queue_fifo_3_data_out[87];
  wire         queue_dataOut_3_store = _queue_fifo_3_data_out[88];
  wire         queue_dataOut_3_issueInst = _queue_fifo_3_data_out[89];
  wire         queue_dataOut_3_loadStore = _queue_fifo_3_data_out[90];
  wire         queue_dataOut_3_decodeResult_logic = _queue_fifo_3_data_out[91];
  wire         queue_dataOut_3_decodeResult_adder = _queue_fifo_3_data_out[92];
  wire         queue_dataOut_3_decodeResult_shift = _queue_fifo_3_data_out[93];
  wire         queue_dataOut_3_decodeResult_multiplier = _queue_fifo_3_data_out[94];
  wire         queue_dataOut_3_decodeResult_divider = _queue_fifo_3_data_out[95];
  wire         queue_dataOut_3_decodeResult_multiCycle = _queue_fifo_3_data_out[96];
  wire         queue_dataOut_3_decodeResult_other = _queue_fifo_3_data_out[97];
  wire         queue_dataOut_3_decodeResult_unsigned0 = _queue_fifo_3_data_out[98];
  wire         queue_dataOut_3_decodeResult_unsigned1 = _queue_fifo_3_data_out[99];
  wire         queue_dataOut_3_decodeResult_itype = _queue_fifo_3_data_out[100];
  wire         queue_dataOut_3_decodeResult_nr = _queue_fifo_3_data_out[101];
  wire         queue_dataOut_3_decodeResult_red = _queue_fifo_3_data_out[102];
  wire         queue_dataOut_3_decodeResult_widenReduce = _queue_fifo_3_data_out[103];
  wire         queue_dataOut_3_decodeResult_targetRd = _queue_fifo_3_data_out[104];
  wire         queue_dataOut_3_decodeResult_slid = _queue_fifo_3_data_out[105];
  wire         queue_dataOut_3_decodeResult_gather = _queue_fifo_3_data_out[106];
  wire         queue_dataOut_3_decodeResult_gather16 = _queue_fifo_3_data_out[107];
  wire         queue_dataOut_3_decodeResult_compress = _queue_fifo_3_data_out[108];
  wire         queue_dataOut_3_decodeResult_unOrderWrite = _queue_fifo_3_data_out[109];
  wire         queue_dataOut_3_decodeResult_extend = _queue_fifo_3_data_out[110];
  wire         queue_dataOut_3_decodeResult_mv = _queue_fifo_3_data_out[111];
  wire         queue_dataOut_3_decodeResult_iota = _queue_fifo_3_data_out[112];
  wire [3:0]   queue_dataOut_3_decodeResult_uop = _queue_fifo_3_data_out[116:113];
  wire         queue_dataOut_3_decodeResult_maskLogic = _queue_fifo_3_data_out[117];
  wire         queue_dataOut_3_decodeResult_maskDestination = _queue_fifo_3_data_out[118];
  wire         queue_dataOut_3_decodeResult_maskSource = _queue_fifo_3_data_out[119];
  wire         queue_dataOut_3_decodeResult_readOnly = _queue_fifo_3_data_out[120];
  wire         queue_dataOut_3_decodeResult_vwmacc = _queue_fifo_3_data_out[121];
  wire         queue_dataOut_3_decodeResult_saturate = _queue_fifo_3_data_out[122];
  wire         queue_dataOut_3_decodeResult_special = _queue_fifo_3_data_out[123];
  wire         queue_dataOut_3_decodeResult_maskUnit = _queue_fifo_3_data_out[124];
  wire         queue_dataOut_3_decodeResult_crossWrite = _queue_fifo_3_data_out[125];
  wire         queue_dataOut_3_decodeResult_crossRead = _queue_fifo_3_data_out[126];
  wire         queue_dataOut_3_decodeResult_sWrite = _queue_fifo_3_data_out[127];
  wire         queue_dataOut_3_decodeResult_vtype = _queue_fifo_3_data_out[128];
  wire         queue_dataOut_3_decodeResult_sReadVD = _queue_fifo_3_data_out[129];
  wire         queue_dataOut_3_decodeResult_scheduler = _queue_fifo_3_data_out[130];
  wire         queue_dataOut_3_decodeResult_dontNeedExecuteInLane = _queue_fifo_3_data_out[131];
  wire         queue_dataOut_3_decodeResult_reverse = _queue_fifo_3_data_out[132];
  wire         queue_dataOut_3_decodeResult_average = _queue_fifo_3_data_out[133];
  wire         queue_dataOut_3_decodeResult_ffo = _queue_fifo_3_data_out[134];
  wire         queue_dataOut_3_decodeResult_popCount = _queue_fifo_3_data_out[135];
  wire [4:0]   queue_dataOut_3_decodeResult_topUop = _queue_fifo_3_data_out[140:136];
  wire         queue_dataOut_3_decodeResult_specialSlot = _queue_fifo_3_data_out[141];
  wire         queue_dataOut_3_decodeResult_float = _queue_fifo_3_data_out[142];
  wire [1:0]   queue_dataOut_3_decodeResult_fpExecutionType = _queue_fifo_3_data_out[144:143];
  wire         queue_dataOut_3_decodeResult_floatMul = _queue_fifo_3_data_out[145];
  wire         queue_dataOut_3_decodeResult_orderReduce = _queue_fifo_3_data_out[146];
  wire [2:0]   queue_dataOut_3_instructionIndex = _queue_fifo_3_data_out[149:147];
  wire         queue_3_enq_ready = ~_queue_fifo_3_full;
  wire         queue_3_enq_valid;
  assign queue_3_deq_valid = ~_queue_fifo_3_empty | queue_3_enq_valid;
  assign queue_3_deq_bits_instructionIndex = _queue_fifo_3_empty ? queue_3_enq_bits_instructionIndex : queue_dataOut_3_instructionIndex;
  assign queue_3_deq_bits_decodeResult_orderReduce = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_orderReduce : queue_dataOut_3_decodeResult_orderReduce;
  assign queue_3_deq_bits_decodeResult_floatMul = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_floatMul : queue_dataOut_3_decodeResult_floatMul;
  assign queue_3_deq_bits_decodeResult_fpExecutionType = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_fpExecutionType : queue_dataOut_3_decodeResult_fpExecutionType;
  assign queue_3_deq_bits_decodeResult_float = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_float : queue_dataOut_3_decodeResult_float;
  assign queue_3_deq_bits_decodeResult_specialSlot = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_specialSlot : queue_dataOut_3_decodeResult_specialSlot;
  assign queue_3_deq_bits_decodeResult_topUop = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_topUop : queue_dataOut_3_decodeResult_topUop;
  assign queue_3_deq_bits_decodeResult_popCount = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_popCount : queue_dataOut_3_decodeResult_popCount;
  assign queue_3_deq_bits_decodeResult_ffo = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_ffo : queue_dataOut_3_decodeResult_ffo;
  assign queue_3_deq_bits_decodeResult_average = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_average : queue_dataOut_3_decodeResult_average;
  assign queue_3_deq_bits_decodeResult_reverse = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_reverse : queue_dataOut_3_decodeResult_reverse;
  assign queue_3_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_3_decodeResult_dontNeedExecuteInLane;
  assign queue_3_deq_bits_decodeResult_scheduler = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_scheduler : queue_dataOut_3_decodeResult_scheduler;
  assign queue_3_deq_bits_decodeResult_sReadVD = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_sReadVD : queue_dataOut_3_decodeResult_sReadVD;
  assign queue_3_deq_bits_decodeResult_vtype = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_vtype : queue_dataOut_3_decodeResult_vtype;
  assign queue_3_deq_bits_decodeResult_sWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_sWrite : queue_dataOut_3_decodeResult_sWrite;
  assign queue_3_deq_bits_decodeResult_crossRead = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_crossRead : queue_dataOut_3_decodeResult_crossRead;
  assign queue_3_deq_bits_decodeResult_crossWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_crossWrite : queue_dataOut_3_decodeResult_crossWrite;
  assign queue_3_deq_bits_decodeResult_maskUnit = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskUnit : queue_dataOut_3_decodeResult_maskUnit;
  assign queue_3_deq_bits_decodeResult_special = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_special : queue_dataOut_3_decodeResult_special;
  assign queue_3_deq_bits_decodeResult_saturate = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_saturate : queue_dataOut_3_decodeResult_saturate;
  assign queue_3_deq_bits_decodeResult_vwmacc = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_vwmacc : queue_dataOut_3_decodeResult_vwmacc;
  assign queue_3_deq_bits_decodeResult_readOnly = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_readOnly : queue_dataOut_3_decodeResult_readOnly;
  assign queue_3_deq_bits_decodeResult_maskSource = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskSource : queue_dataOut_3_decodeResult_maskSource;
  assign queue_3_deq_bits_decodeResult_maskDestination = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskDestination : queue_dataOut_3_decodeResult_maskDestination;
  assign queue_3_deq_bits_decodeResult_maskLogic = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskLogic : queue_dataOut_3_decodeResult_maskLogic;
  assign queue_3_deq_bits_decodeResult_uop = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_uop : queue_dataOut_3_decodeResult_uop;
  assign queue_3_deq_bits_decodeResult_iota = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_iota : queue_dataOut_3_decodeResult_iota;
  assign queue_3_deq_bits_decodeResult_mv = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_mv : queue_dataOut_3_decodeResult_mv;
  assign queue_3_deq_bits_decodeResult_extend = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_extend : queue_dataOut_3_decodeResult_extend;
  assign queue_3_deq_bits_decodeResult_unOrderWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unOrderWrite : queue_dataOut_3_decodeResult_unOrderWrite;
  assign queue_3_deq_bits_decodeResult_compress = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_compress : queue_dataOut_3_decodeResult_compress;
  assign queue_3_deq_bits_decodeResult_gather16 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_gather16 : queue_dataOut_3_decodeResult_gather16;
  assign queue_3_deq_bits_decodeResult_gather = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_gather : queue_dataOut_3_decodeResult_gather;
  assign queue_3_deq_bits_decodeResult_slid = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_slid : queue_dataOut_3_decodeResult_slid;
  assign queue_3_deq_bits_decodeResult_targetRd = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_targetRd : queue_dataOut_3_decodeResult_targetRd;
  assign queue_3_deq_bits_decodeResult_widenReduce = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_widenReduce : queue_dataOut_3_decodeResult_widenReduce;
  assign queue_3_deq_bits_decodeResult_red = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_red : queue_dataOut_3_decodeResult_red;
  assign queue_3_deq_bits_decodeResult_nr = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_nr : queue_dataOut_3_decodeResult_nr;
  assign queue_3_deq_bits_decodeResult_itype = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_itype : queue_dataOut_3_decodeResult_itype;
  assign queue_3_deq_bits_decodeResult_unsigned1 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unsigned1 : queue_dataOut_3_decodeResult_unsigned1;
  assign queue_3_deq_bits_decodeResult_unsigned0 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unsigned0 : queue_dataOut_3_decodeResult_unsigned0;
  assign queue_3_deq_bits_decodeResult_other = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_other : queue_dataOut_3_decodeResult_other;
  assign queue_3_deq_bits_decodeResult_multiCycle = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_multiCycle : queue_dataOut_3_decodeResult_multiCycle;
  assign queue_3_deq_bits_decodeResult_divider = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_divider : queue_dataOut_3_decodeResult_divider;
  assign queue_3_deq_bits_decodeResult_multiplier = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_multiplier : queue_dataOut_3_decodeResult_multiplier;
  assign queue_3_deq_bits_decodeResult_shift = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_shift : queue_dataOut_3_decodeResult_shift;
  assign queue_3_deq_bits_decodeResult_adder = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_adder : queue_dataOut_3_decodeResult_adder;
  assign queue_3_deq_bits_decodeResult_logic = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_logic : queue_dataOut_3_decodeResult_logic;
  assign queue_3_deq_bits_loadStore = _queue_fifo_3_empty ? queue_3_enq_bits_loadStore : queue_dataOut_3_loadStore;
  assign queue_3_deq_bits_issueInst = _queue_fifo_3_empty ? queue_3_enq_bits_issueInst : queue_dataOut_3_issueInst;
  assign queue_3_deq_bits_store = _queue_fifo_3_empty ? queue_3_enq_bits_store : queue_dataOut_3_store;
  assign queue_3_deq_bits_special = _queue_fifo_3_empty ? queue_3_enq_bits_special : queue_dataOut_3_special;
  assign queue_3_deq_bits_lsWholeReg = _queue_fifo_3_empty ? queue_3_enq_bits_lsWholeReg : queue_dataOut_3_lsWholeReg;
  assign queue_3_deq_bits_vs1 = _queue_fifo_3_empty ? queue_3_enq_bits_vs1 : queue_dataOut_3_vs1;
  assign queue_3_deq_bits_vs2 = _queue_fifo_3_empty ? queue_3_enq_bits_vs2 : queue_dataOut_3_vs2;
  assign queue_3_deq_bits_vd = _queue_fifo_3_empty ? queue_3_enq_bits_vd : queue_dataOut_3_vd;
  assign queue_3_deq_bits_loadStoreEEW = _queue_fifo_3_empty ? queue_3_enq_bits_loadStoreEEW : queue_dataOut_3_loadStoreEEW;
  assign queue_3_deq_bits_mask = _queue_fifo_3_empty ? queue_3_enq_bits_mask : queue_dataOut_3_mask;
  assign queue_3_deq_bits_segment = _queue_fifo_3_empty ? queue_3_enq_bits_segment : queue_dataOut_3_segment;
  assign queue_3_deq_bits_readFromScalar = _queue_fifo_3_empty ? queue_3_enq_bits_readFromScalar : queue_dataOut_3_readFromScalar;
  assign queue_3_deq_bits_csrInterface_vl = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vl : queue_dataOut_3_csrInterface_vl;
  assign queue_3_deq_bits_csrInterface_vStart = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vStart : queue_dataOut_3_csrInterface_vStart;
  assign queue_3_deq_bits_csrInterface_vlmul = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vlmul : queue_dataOut_3_csrInterface_vlmul;
  assign queue_3_deq_bits_csrInterface_vSew = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vSew : queue_dataOut_3_csrInterface_vSew;
  assign queue_3_deq_bits_csrInterface_vxrm = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vxrm : queue_dataOut_3_csrInterface_vxrm;
  assign queue_3_deq_bits_csrInterface_vta = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vta : queue_dataOut_3_csrInterface_vta;
  assign queue_3_deq_bits_csrInterface_vma = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vma : queue_dataOut_3_csrInterface_vma;
  wire         laneVec_3_laneRequest_bits_issueInst = laneRequestSinkWire_3_ready & laneRequestSinkWire_3_valid;
  reg          releasePipe_pipe_v_3;
  wire         releasePipe_pipe_out_3_valid = releasePipe_pipe_v_3;
  wire         laneRequestSourceWire_3_ready;
  wire         validSource_3_valid = laneRequestSourceWire_3_ready & laneRequestSourceWire_3_valid;
  reg  [2:0]   tokenCheck_counter_3;
  wire [2:0]   tokenCheck_counterChange_3 = validSource_3_valid ? 3'h1 : 3'h7;
  assign tokenCheck_3 = ~(tokenCheck_counter_3[2]);
  assign laneRequestSourceWire_3_ready = tokenCheck_3;
  assign queue_3_enq_valid = validSink_3_valid;
  assign queue_3_enq_bits_instructionIndex = validSink_3_bits_instructionIndex;
  assign queue_3_enq_bits_decodeResult_orderReduce = validSink_3_bits_decodeResult_orderReduce;
  assign queue_3_enq_bits_decodeResult_floatMul = validSink_3_bits_decodeResult_floatMul;
  assign queue_3_enq_bits_decodeResult_fpExecutionType = validSink_3_bits_decodeResult_fpExecutionType;
  assign queue_3_enq_bits_decodeResult_float = validSink_3_bits_decodeResult_float;
  assign queue_3_enq_bits_decodeResult_specialSlot = validSink_3_bits_decodeResult_specialSlot;
  assign queue_3_enq_bits_decodeResult_topUop = validSink_3_bits_decodeResult_topUop;
  assign queue_3_enq_bits_decodeResult_popCount = validSink_3_bits_decodeResult_popCount;
  assign queue_3_enq_bits_decodeResult_ffo = validSink_3_bits_decodeResult_ffo;
  assign queue_3_enq_bits_decodeResult_average = validSink_3_bits_decodeResult_average;
  assign queue_3_enq_bits_decodeResult_reverse = validSink_3_bits_decodeResult_reverse;
  assign queue_3_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_3_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_3_enq_bits_decodeResult_scheduler = validSink_3_bits_decodeResult_scheduler;
  assign queue_3_enq_bits_decodeResult_sReadVD = validSink_3_bits_decodeResult_sReadVD;
  assign queue_3_enq_bits_decodeResult_vtype = validSink_3_bits_decodeResult_vtype;
  assign queue_3_enq_bits_decodeResult_sWrite = validSink_3_bits_decodeResult_sWrite;
  assign queue_3_enq_bits_decodeResult_crossRead = validSink_3_bits_decodeResult_crossRead;
  assign queue_3_enq_bits_decodeResult_crossWrite = validSink_3_bits_decodeResult_crossWrite;
  assign queue_3_enq_bits_decodeResult_maskUnit = validSink_3_bits_decodeResult_maskUnit;
  assign queue_3_enq_bits_decodeResult_special = validSink_3_bits_decodeResult_special;
  assign queue_3_enq_bits_decodeResult_saturate = validSink_3_bits_decodeResult_saturate;
  assign queue_3_enq_bits_decodeResult_vwmacc = validSink_3_bits_decodeResult_vwmacc;
  assign queue_3_enq_bits_decodeResult_readOnly = validSink_3_bits_decodeResult_readOnly;
  assign queue_3_enq_bits_decodeResult_maskSource = validSink_3_bits_decodeResult_maskSource;
  assign queue_3_enq_bits_decodeResult_maskDestination = validSink_3_bits_decodeResult_maskDestination;
  assign queue_3_enq_bits_decodeResult_maskLogic = validSink_3_bits_decodeResult_maskLogic;
  assign queue_3_enq_bits_decodeResult_uop = validSink_3_bits_decodeResult_uop;
  assign queue_3_enq_bits_decodeResult_iota = validSink_3_bits_decodeResult_iota;
  assign queue_3_enq_bits_decodeResult_mv = validSink_3_bits_decodeResult_mv;
  assign queue_3_enq_bits_decodeResult_extend = validSink_3_bits_decodeResult_extend;
  assign queue_3_enq_bits_decodeResult_unOrderWrite = validSink_3_bits_decodeResult_unOrderWrite;
  assign queue_3_enq_bits_decodeResult_compress = validSink_3_bits_decodeResult_compress;
  assign queue_3_enq_bits_decodeResult_gather16 = validSink_3_bits_decodeResult_gather16;
  assign queue_3_enq_bits_decodeResult_gather = validSink_3_bits_decodeResult_gather;
  assign queue_3_enq_bits_decodeResult_slid = validSink_3_bits_decodeResult_slid;
  assign queue_3_enq_bits_decodeResult_targetRd = validSink_3_bits_decodeResult_targetRd;
  assign queue_3_enq_bits_decodeResult_widenReduce = validSink_3_bits_decodeResult_widenReduce;
  assign queue_3_enq_bits_decodeResult_red = validSink_3_bits_decodeResult_red;
  assign queue_3_enq_bits_decodeResult_nr = validSink_3_bits_decodeResult_nr;
  assign queue_3_enq_bits_decodeResult_itype = validSink_3_bits_decodeResult_itype;
  assign queue_3_enq_bits_decodeResult_unsigned1 = validSink_3_bits_decodeResult_unsigned1;
  assign queue_3_enq_bits_decodeResult_unsigned0 = validSink_3_bits_decodeResult_unsigned0;
  assign queue_3_enq_bits_decodeResult_other = validSink_3_bits_decodeResult_other;
  assign queue_3_enq_bits_decodeResult_multiCycle = validSink_3_bits_decodeResult_multiCycle;
  assign queue_3_enq_bits_decodeResult_divider = validSink_3_bits_decodeResult_divider;
  assign queue_3_enq_bits_decodeResult_multiplier = validSink_3_bits_decodeResult_multiplier;
  assign queue_3_enq_bits_decodeResult_shift = validSink_3_bits_decodeResult_shift;
  assign queue_3_enq_bits_decodeResult_adder = validSink_3_bits_decodeResult_adder;
  assign queue_3_enq_bits_decodeResult_logic = validSink_3_bits_decodeResult_logic;
  assign queue_3_enq_bits_loadStore = validSink_3_bits_loadStore;
  assign queue_3_enq_bits_issueInst = validSink_3_bits_issueInst;
  assign queue_3_enq_bits_store = validSink_3_bits_store;
  assign queue_3_enq_bits_special = validSink_3_bits_special;
  assign queue_3_enq_bits_lsWholeReg = validSink_3_bits_lsWholeReg;
  assign queue_3_enq_bits_vs1 = validSink_3_bits_vs1;
  assign queue_3_enq_bits_vs2 = validSink_3_bits_vs2;
  assign queue_3_enq_bits_vd = validSink_3_bits_vd;
  assign queue_3_enq_bits_loadStoreEEW = validSink_3_bits_loadStoreEEW;
  assign queue_3_enq_bits_mask = validSink_3_bits_mask;
  assign queue_3_enq_bits_segment = validSink_3_bits_segment;
  assign queue_3_enq_bits_readFromScalar = validSink_3_bits_readFromScalar;
  assign queue_3_enq_bits_csrInterface_vl = validSink_3_bits_csrInterface_vl;
  assign queue_3_enq_bits_csrInterface_vStart = validSink_3_bits_csrInterface_vStart;
  assign queue_3_enq_bits_csrInterface_vlmul = validSink_3_bits_csrInterface_vlmul;
  assign queue_3_enq_bits_csrInterface_vSew = validSink_3_bits_csrInterface_vSew;
  assign queue_3_enq_bits_csrInterface_vxrm = validSink_3_bits_csrInterface_vxrm;
  assign queue_3_enq_bits_csrInterface_vta = validSink_3_bits_csrInterface_vta;
  assign queue_3_enq_bits_csrInterface_vma = validSink_3_bits_csrInterface_vma;
  reg          shifterReg_3_0_valid;
  assign validSink_3_valid = shifterReg_3_0_valid;
  reg  [2:0]   shifterReg_3_0_bits_instructionIndex;
  assign validSink_3_bits_instructionIndex = shifterReg_3_0_bits_instructionIndex;
  reg          shifterReg_3_0_bits_decodeResult_orderReduce;
  assign validSink_3_bits_decodeResult_orderReduce = shifterReg_3_0_bits_decodeResult_orderReduce;
  reg          shifterReg_3_0_bits_decodeResult_floatMul;
  assign validSink_3_bits_decodeResult_floatMul = shifterReg_3_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_3_0_bits_decodeResult_fpExecutionType;
  assign validSink_3_bits_decodeResult_fpExecutionType = shifterReg_3_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_3_0_bits_decodeResult_float;
  assign validSink_3_bits_decodeResult_float = shifterReg_3_0_bits_decodeResult_float;
  reg          shifterReg_3_0_bits_decodeResult_specialSlot;
  assign validSink_3_bits_decodeResult_specialSlot = shifterReg_3_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_3_0_bits_decodeResult_topUop;
  assign validSink_3_bits_decodeResult_topUop = shifterReg_3_0_bits_decodeResult_topUop;
  reg          shifterReg_3_0_bits_decodeResult_popCount;
  assign validSink_3_bits_decodeResult_popCount = shifterReg_3_0_bits_decodeResult_popCount;
  reg          shifterReg_3_0_bits_decodeResult_ffo;
  assign validSink_3_bits_decodeResult_ffo = shifterReg_3_0_bits_decodeResult_ffo;
  reg          shifterReg_3_0_bits_decodeResult_average;
  assign validSink_3_bits_decodeResult_average = shifterReg_3_0_bits_decodeResult_average;
  reg          shifterReg_3_0_bits_decodeResult_reverse;
  assign validSink_3_bits_decodeResult_reverse = shifterReg_3_0_bits_decodeResult_reverse;
  reg          shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_3_bits_decodeResult_dontNeedExecuteInLane = shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_3_0_bits_decodeResult_scheduler;
  assign validSink_3_bits_decodeResult_scheduler = shifterReg_3_0_bits_decodeResult_scheduler;
  reg          shifterReg_3_0_bits_decodeResult_sReadVD;
  assign validSink_3_bits_decodeResult_sReadVD = shifterReg_3_0_bits_decodeResult_sReadVD;
  reg          shifterReg_3_0_bits_decodeResult_vtype;
  assign validSink_3_bits_decodeResult_vtype = shifterReg_3_0_bits_decodeResult_vtype;
  reg          shifterReg_3_0_bits_decodeResult_sWrite;
  assign validSink_3_bits_decodeResult_sWrite = shifterReg_3_0_bits_decodeResult_sWrite;
  reg          shifterReg_3_0_bits_decodeResult_crossRead;
  assign validSink_3_bits_decodeResult_crossRead = shifterReg_3_0_bits_decodeResult_crossRead;
  reg          shifterReg_3_0_bits_decodeResult_crossWrite;
  assign validSink_3_bits_decodeResult_crossWrite = shifterReg_3_0_bits_decodeResult_crossWrite;
  reg          shifterReg_3_0_bits_decodeResult_maskUnit;
  assign validSink_3_bits_decodeResult_maskUnit = shifterReg_3_0_bits_decodeResult_maskUnit;
  reg          shifterReg_3_0_bits_decodeResult_special;
  assign validSink_3_bits_decodeResult_special = shifterReg_3_0_bits_decodeResult_special;
  reg          shifterReg_3_0_bits_decodeResult_saturate;
  assign validSink_3_bits_decodeResult_saturate = shifterReg_3_0_bits_decodeResult_saturate;
  reg          shifterReg_3_0_bits_decodeResult_vwmacc;
  assign validSink_3_bits_decodeResult_vwmacc = shifterReg_3_0_bits_decodeResult_vwmacc;
  reg          shifterReg_3_0_bits_decodeResult_readOnly;
  assign validSink_3_bits_decodeResult_readOnly = shifterReg_3_0_bits_decodeResult_readOnly;
  reg          shifterReg_3_0_bits_decodeResult_maskSource;
  assign validSink_3_bits_decodeResult_maskSource = shifterReg_3_0_bits_decodeResult_maskSource;
  reg          shifterReg_3_0_bits_decodeResult_maskDestination;
  assign validSink_3_bits_decodeResult_maskDestination = shifterReg_3_0_bits_decodeResult_maskDestination;
  reg          shifterReg_3_0_bits_decodeResult_maskLogic;
  assign validSink_3_bits_decodeResult_maskLogic = shifterReg_3_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_3_0_bits_decodeResult_uop;
  assign validSink_3_bits_decodeResult_uop = shifterReg_3_0_bits_decodeResult_uop;
  reg          shifterReg_3_0_bits_decodeResult_iota;
  assign validSink_3_bits_decodeResult_iota = shifterReg_3_0_bits_decodeResult_iota;
  reg          shifterReg_3_0_bits_decodeResult_mv;
  assign validSink_3_bits_decodeResult_mv = shifterReg_3_0_bits_decodeResult_mv;
  reg          shifterReg_3_0_bits_decodeResult_extend;
  assign validSink_3_bits_decodeResult_extend = shifterReg_3_0_bits_decodeResult_extend;
  reg          shifterReg_3_0_bits_decodeResult_unOrderWrite;
  assign validSink_3_bits_decodeResult_unOrderWrite = shifterReg_3_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_3_0_bits_decodeResult_compress;
  assign validSink_3_bits_decodeResult_compress = shifterReg_3_0_bits_decodeResult_compress;
  reg          shifterReg_3_0_bits_decodeResult_gather16;
  assign validSink_3_bits_decodeResult_gather16 = shifterReg_3_0_bits_decodeResult_gather16;
  reg          shifterReg_3_0_bits_decodeResult_gather;
  assign validSink_3_bits_decodeResult_gather = shifterReg_3_0_bits_decodeResult_gather;
  reg          shifterReg_3_0_bits_decodeResult_slid;
  assign validSink_3_bits_decodeResult_slid = shifterReg_3_0_bits_decodeResult_slid;
  reg          shifterReg_3_0_bits_decodeResult_targetRd;
  assign validSink_3_bits_decodeResult_targetRd = shifterReg_3_0_bits_decodeResult_targetRd;
  reg          shifterReg_3_0_bits_decodeResult_widenReduce;
  assign validSink_3_bits_decodeResult_widenReduce = shifterReg_3_0_bits_decodeResult_widenReduce;
  reg          shifterReg_3_0_bits_decodeResult_red;
  assign validSink_3_bits_decodeResult_red = shifterReg_3_0_bits_decodeResult_red;
  reg          shifterReg_3_0_bits_decodeResult_nr;
  assign validSink_3_bits_decodeResult_nr = shifterReg_3_0_bits_decodeResult_nr;
  reg          shifterReg_3_0_bits_decodeResult_itype;
  assign validSink_3_bits_decodeResult_itype = shifterReg_3_0_bits_decodeResult_itype;
  reg          shifterReg_3_0_bits_decodeResult_unsigned1;
  assign validSink_3_bits_decodeResult_unsigned1 = shifterReg_3_0_bits_decodeResult_unsigned1;
  reg          shifterReg_3_0_bits_decodeResult_unsigned0;
  assign validSink_3_bits_decodeResult_unsigned0 = shifterReg_3_0_bits_decodeResult_unsigned0;
  reg          shifterReg_3_0_bits_decodeResult_other;
  assign validSink_3_bits_decodeResult_other = shifterReg_3_0_bits_decodeResult_other;
  reg          shifterReg_3_0_bits_decodeResult_multiCycle;
  assign validSink_3_bits_decodeResult_multiCycle = shifterReg_3_0_bits_decodeResult_multiCycle;
  reg          shifterReg_3_0_bits_decodeResult_divider;
  assign validSink_3_bits_decodeResult_divider = shifterReg_3_0_bits_decodeResult_divider;
  reg          shifterReg_3_0_bits_decodeResult_multiplier;
  assign validSink_3_bits_decodeResult_multiplier = shifterReg_3_0_bits_decodeResult_multiplier;
  reg          shifterReg_3_0_bits_decodeResult_shift;
  assign validSink_3_bits_decodeResult_shift = shifterReg_3_0_bits_decodeResult_shift;
  reg          shifterReg_3_0_bits_decodeResult_adder;
  assign validSink_3_bits_decodeResult_adder = shifterReg_3_0_bits_decodeResult_adder;
  reg          shifterReg_3_0_bits_decodeResult_logic;
  assign validSink_3_bits_decodeResult_logic = shifterReg_3_0_bits_decodeResult_logic;
  reg          shifterReg_3_0_bits_loadStore;
  assign validSink_3_bits_loadStore = shifterReg_3_0_bits_loadStore;
  reg          shifterReg_3_0_bits_issueInst;
  assign validSink_3_bits_issueInst = shifterReg_3_0_bits_issueInst;
  reg          shifterReg_3_0_bits_store;
  assign validSink_3_bits_store = shifterReg_3_0_bits_store;
  reg          shifterReg_3_0_bits_special;
  assign validSink_3_bits_special = shifterReg_3_0_bits_special;
  reg          shifterReg_3_0_bits_lsWholeReg;
  assign validSink_3_bits_lsWholeReg = shifterReg_3_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_3_0_bits_vs1;
  assign validSink_3_bits_vs1 = shifterReg_3_0_bits_vs1;
  reg  [4:0]   shifterReg_3_0_bits_vs2;
  assign validSink_3_bits_vs2 = shifterReg_3_0_bits_vs2;
  reg  [4:0]   shifterReg_3_0_bits_vd;
  assign validSink_3_bits_vd = shifterReg_3_0_bits_vd;
  reg  [1:0]   shifterReg_3_0_bits_loadStoreEEW;
  assign validSink_3_bits_loadStoreEEW = shifterReg_3_0_bits_loadStoreEEW;
  reg          shifterReg_3_0_bits_mask;
  assign validSink_3_bits_mask = shifterReg_3_0_bits_mask;
  reg  [2:0]   shifterReg_3_0_bits_segment;
  assign validSink_3_bits_segment = shifterReg_3_0_bits_segment;
  reg  [31:0]  shifterReg_3_0_bits_readFromScalar;
  assign validSink_3_bits_readFromScalar = shifterReg_3_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_3_0_bits_csrInterface_vl;
  assign validSink_3_bits_csrInterface_vl = shifterReg_3_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_3_0_bits_csrInterface_vStart;
  assign validSink_3_bits_csrInterface_vStart = shifterReg_3_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_3_0_bits_csrInterface_vlmul;
  assign validSink_3_bits_csrInterface_vlmul = shifterReg_3_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_3_0_bits_csrInterface_vSew;
  assign validSink_3_bits_csrInterface_vSew = shifterReg_3_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_3_0_bits_csrInterface_vxrm;
  assign validSink_3_bits_csrInterface_vxrm = shifterReg_3_0_bits_csrInterface_vxrm;
  reg          shifterReg_3_0_bits_csrInterface_vta;
  assign validSink_3_bits_csrInterface_vta = shifterReg_3_0_bits_csrInterface_vta;
  reg          shifterReg_3_0_bits_csrInterface_vma;
  assign validSink_3_bits_csrInterface_vma = shifterReg_3_0_bits_csrInterface_vma;
  wire         shifterValid_3 = shifterReg_3_0_valid | validSource_3_valid;
  wire         validSink_4_valid;
  wire [2:0]   validSink_4_bits_instructionIndex;
  wire         validSink_4_bits_decodeResult_orderReduce;
  wire         validSink_4_bits_decodeResult_floatMul;
  wire [1:0]   validSink_4_bits_decodeResult_fpExecutionType;
  wire         validSink_4_bits_decodeResult_float;
  wire         validSink_4_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_4_bits_decodeResult_topUop;
  wire         validSink_4_bits_decodeResult_popCount;
  wire         validSink_4_bits_decodeResult_ffo;
  wire         validSink_4_bits_decodeResult_average;
  wire         validSink_4_bits_decodeResult_reverse;
  wire         validSink_4_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_4_bits_decodeResult_scheduler;
  wire         validSink_4_bits_decodeResult_sReadVD;
  wire         validSink_4_bits_decodeResult_vtype;
  wire         validSink_4_bits_decodeResult_sWrite;
  wire         validSink_4_bits_decodeResult_crossRead;
  wire         validSink_4_bits_decodeResult_crossWrite;
  wire         validSink_4_bits_decodeResult_maskUnit;
  wire         validSink_4_bits_decodeResult_special;
  wire         validSink_4_bits_decodeResult_saturate;
  wire         validSink_4_bits_decodeResult_vwmacc;
  wire         validSink_4_bits_decodeResult_readOnly;
  wire         validSink_4_bits_decodeResult_maskSource;
  wire         validSink_4_bits_decodeResult_maskDestination;
  wire         validSink_4_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_4_bits_decodeResult_uop;
  wire         validSink_4_bits_decodeResult_iota;
  wire         validSink_4_bits_decodeResult_mv;
  wire         validSink_4_bits_decodeResult_extend;
  wire         validSink_4_bits_decodeResult_unOrderWrite;
  wire         validSink_4_bits_decodeResult_compress;
  wire         validSink_4_bits_decodeResult_gather16;
  wire         validSink_4_bits_decodeResult_gather;
  wire         validSink_4_bits_decodeResult_slid;
  wire         validSink_4_bits_decodeResult_targetRd;
  wire         validSink_4_bits_decodeResult_widenReduce;
  wire         validSink_4_bits_decodeResult_red;
  wire         validSink_4_bits_decodeResult_nr;
  wire         validSink_4_bits_decodeResult_itype;
  wire         validSink_4_bits_decodeResult_unsigned1;
  wire         validSink_4_bits_decodeResult_unsigned0;
  wire         validSink_4_bits_decodeResult_other;
  wire         validSink_4_bits_decodeResult_multiCycle;
  wire         validSink_4_bits_decodeResult_divider;
  wire         validSink_4_bits_decodeResult_multiplier;
  wire         validSink_4_bits_decodeResult_shift;
  wire         validSink_4_bits_decodeResult_adder;
  wire         validSink_4_bits_decodeResult_logic;
  wire         validSink_4_bits_loadStore;
  wire         validSink_4_bits_issueInst;
  wire         validSink_4_bits_store;
  wire         validSink_4_bits_special;
  wire         validSink_4_bits_lsWholeReg;
  wire [4:0]   validSink_4_bits_vs1;
  wire [4:0]   validSink_4_bits_vs2;
  wire [4:0]   validSink_4_bits_vd;
  wire [1:0]   validSink_4_bits_loadStoreEEW;
  wire         validSink_4_bits_mask;
  wire [2:0]   validSink_4_bits_segment;
  wire [31:0]  validSink_4_bits_readFromScalar;
  wire [11:0]  validSink_4_bits_csrInterface_vl;
  wire [11:0]  validSink_4_bits_csrInterface_vStart;
  wire [2:0]   validSink_4_bits_csrInterface_vlmul;
  wire [1:0]   validSink_4_bits_csrInterface_vSew;
  wire [1:0]   validSink_4_bits_csrInterface_vxrm;
  wire         validSink_4_bits_csrInterface_vta;
  wire         validSink_4_bits_csrInterface_vma;
  wire         laneRequestSinkWire_4_valid = queue_4_deq_valid;
  wire [2:0]   laneRequestSinkWire_4_bits_instructionIndex = queue_4_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_4_bits_decodeResult_orderReduce = queue_4_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_4_bits_decodeResult_floatMul = queue_4_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_4_bits_decodeResult_fpExecutionType = queue_4_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_4_bits_decodeResult_float = queue_4_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_4_bits_decodeResult_specialSlot = queue_4_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_4_bits_decodeResult_topUop = queue_4_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_4_bits_decodeResult_popCount = queue_4_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_4_bits_decodeResult_ffo = queue_4_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_4_bits_decodeResult_average = queue_4_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_4_bits_decodeResult_reverse = queue_4_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_4_bits_decodeResult_dontNeedExecuteInLane = queue_4_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_4_bits_decodeResult_scheduler = queue_4_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_4_bits_decodeResult_sReadVD = queue_4_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_4_bits_decodeResult_vtype = queue_4_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_4_bits_decodeResult_sWrite = queue_4_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_crossRead = queue_4_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_4_bits_decodeResult_crossWrite = queue_4_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskUnit = queue_4_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_4_bits_decodeResult_special = queue_4_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_4_bits_decodeResult_saturate = queue_4_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_4_bits_decodeResult_vwmacc = queue_4_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_4_bits_decodeResult_readOnly = queue_4_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskSource = queue_4_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskDestination = queue_4_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskLogic = queue_4_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_4_bits_decodeResult_uop = queue_4_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_4_bits_decodeResult_iota = queue_4_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_4_bits_decodeResult_mv = queue_4_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_4_bits_decodeResult_extend = queue_4_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_4_bits_decodeResult_unOrderWrite = queue_4_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_compress = queue_4_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_4_bits_decodeResult_gather16 = queue_4_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_4_bits_decodeResult_gather = queue_4_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_4_bits_decodeResult_slid = queue_4_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_4_bits_decodeResult_targetRd = queue_4_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_4_bits_decodeResult_widenReduce = queue_4_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_4_bits_decodeResult_red = queue_4_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_4_bits_decodeResult_nr = queue_4_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_4_bits_decodeResult_itype = queue_4_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_4_bits_decodeResult_unsigned1 = queue_4_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_4_bits_decodeResult_unsigned0 = queue_4_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_4_bits_decodeResult_other = queue_4_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_4_bits_decodeResult_multiCycle = queue_4_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_4_bits_decodeResult_divider = queue_4_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_4_bits_decodeResult_multiplier = queue_4_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_4_bits_decodeResult_shift = queue_4_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_4_bits_decodeResult_adder = queue_4_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_4_bits_decodeResult_logic = queue_4_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_4_bits_loadStore = queue_4_deq_bits_loadStore;
  wire         laneRequestSinkWire_4_bits_issueInst = queue_4_deq_bits_issueInst;
  wire         laneRequestSinkWire_4_bits_store = queue_4_deq_bits_store;
  wire         laneRequestSinkWire_4_bits_special = queue_4_deq_bits_special;
  wire         laneRequestSinkWire_4_bits_lsWholeReg = queue_4_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_4_bits_vs1 = queue_4_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_4_bits_vs2 = queue_4_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_4_bits_vd = queue_4_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_4_bits_loadStoreEEW = queue_4_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_4_bits_mask = queue_4_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_4_bits_segment = queue_4_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_4_bits_readFromScalar = queue_4_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_4_bits_csrInterface_vl = queue_4_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_4_bits_csrInterface_vStart = queue_4_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_4_bits_csrInterface_vlmul = queue_4_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_4_bits_csrInterface_vSew = queue_4_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_4_bits_csrInterface_vxrm = queue_4_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_4_bits_csrInterface_vta = queue_4_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_4_bits_csrInterface_vma = queue_4_deq_bits_csrInterface_vma;
  wire [1:0]   queue_4_enq_bits_csrInterface_vxrm;
  wire         queue_4_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_12 = {queue_4_enq_bits_csrInterface_vxrm, queue_4_enq_bits_csrInterface_vta};
  wire         queue_4_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_12 = {queue_dataIn_lo_hi_12, queue_4_enq_bits_csrInterface_vma};
  wire [2:0]   queue_4_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_4_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_12 = {queue_4_enq_bits_csrInterface_vlmul, queue_4_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_4_enq_bits_csrInterface_vl;
  wire [11:0]  queue_4_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_12 = {queue_4_enq_bits_csrInterface_vl, queue_4_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_12 = {queue_dataIn_hi_hi_12, queue_dataIn_hi_lo_12};
  wire         queue_4_enq_bits_decodeResult_shift;
  wire         queue_4_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_4 = {queue_4_enq_bits_decodeResult_shift, queue_4_enq_bits_decodeResult_adder};
  wire         queue_4_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_4 = {queue_dataIn_lo_lo_lo_lo_hi_4, queue_4_enq_bits_decodeResult_logic};
  wire         queue_4_enq_bits_decodeResult_multiCycle;
  wire         queue_4_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_multiCycle, queue_4_enq_bits_decodeResult_divider};
  wire         queue_4_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_4 = {queue_dataIn_lo_lo_lo_hi_hi_4, queue_4_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_4 = {queue_dataIn_lo_lo_lo_hi_4, queue_dataIn_lo_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_unsigned1;
  wire         queue_4_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_unsigned1, queue_4_enq_bits_decodeResult_unsigned0};
  wire         queue_4_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_4 = {queue_dataIn_lo_lo_hi_lo_hi_4, queue_4_enq_bits_decodeResult_other};
  wire         queue_4_enq_bits_decodeResult_red;
  wire         queue_4_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_red, queue_4_enq_bits_decodeResult_nr};
  wire         queue_4_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_4 = {queue_dataIn_lo_lo_hi_hi_hi_4, queue_4_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_8 = {queue_dataIn_lo_lo_hi_hi_4, queue_dataIn_lo_lo_hi_lo_4};
  wire [11:0]  queue_dataIn_lo_lo_8 = {queue_dataIn_lo_lo_hi_8, queue_dataIn_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_slid;
  wire         queue_4_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_4 = {queue_4_enq_bits_decodeResult_slid, queue_4_enq_bits_decodeResult_targetRd};
  wire         queue_4_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_4 = {queue_dataIn_lo_hi_lo_lo_hi_4, queue_4_enq_bits_decodeResult_widenReduce};
  wire         queue_4_enq_bits_decodeResult_compress;
  wire         queue_4_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_compress, queue_4_enq_bits_decodeResult_gather16};
  wire         queue_4_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_4 = {queue_dataIn_lo_hi_lo_hi_hi_4, queue_4_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_8 = {queue_dataIn_lo_hi_lo_hi_4, queue_dataIn_lo_hi_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_mv;
  wire         queue_4_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_mv, queue_4_enq_bits_decodeResult_extend};
  wire         queue_4_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_4 = {queue_dataIn_lo_hi_hi_lo_hi_4, queue_4_enq_bits_decodeResult_unOrderWrite};
  wire         queue_4_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_4_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_maskLogic, queue_4_enq_bits_decodeResult_uop};
  wire         queue_4_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_4 = {queue_dataIn_lo_hi_hi_hi_hi_4, queue_4_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_8 = {queue_dataIn_lo_hi_hi_hi_4, queue_dataIn_lo_hi_hi_lo_4};
  wire [14:0]  queue_dataIn_lo_hi_13 = {queue_dataIn_lo_hi_hi_8, queue_dataIn_lo_hi_lo_8};
  wire [26:0]  queue_dataIn_lo_13 = {queue_dataIn_lo_hi_13, queue_dataIn_lo_lo_8};
  wire         queue_4_enq_bits_decodeResult_readOnly;
  wire         queue_4_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_4 = {queue_4_enq_bits_decodeResult_readOnly, queue_4_enq_bits_decodeResult_maskSource};
  wire         queue_4_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_4 = {queue_dataIn_hi_lo_lo_lo_hi_4, queue_4_enq_bits_decodeResult_maskDestination};
  wire         queue_4_enq_bits_decodeResult_special;
  wire         queue_4_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_special, queue_4_enq_bits_decodeResult_saturate};
  wire         queue_4_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_4 = {queue_dataIn_hi_lo_lo_hi_hi_4, queue_4_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_8 = {queue_dataIn_hi_lo_lo_hi_4, queue_dataIn_hi_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_crossRead;
  wire         queue_4_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_crossRead, queue_4_enq_bits_decodeResult_crossWrite};
  wire         queue_4_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_4 = {queue_dataIn_hi_lo_hi_lo_hi_4, queue_4_enq_bits_decodeResult_maskUnit};
  wire         queue_4_enq_bits_decodeResult_sReadVD;
  wire         queue_4_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_sReadVD, queue_4_enq_bits_decodeResult_vtype};
  wire         queue_4_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_4 = {queue_dataIn_hi_lo_hi_hi_hi_4, queue_4_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_8 = {queue_dataIn_hi_lo_hi_hi_4, queue_dataIn_hi_lo_hi_lo_4};
  wire [11:0]  queue_dataIn_hi_lo_13 = {queue_dataIn_hi_lo_hi_8, queue_dataIn_hi_lo_lo_8};
  wire         queue_4_enq_bits_decodeResult_reverse;
  wire         queue_4_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_4 = {queue_4_enq_bits_decodeResult_reverse, queue_4_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_4_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_4 = {queue_dataIn_hi_hi_lo_lo_hi_4, queue_4_enq_bits_decodeResult_scheduler};
  wire         queue_4_enq_bits_decodeResult_popCount;
  wire         queue_4_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_popCount, queue_4_enq_bits_decodeResult_ffo};
  wire         queue_4_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_4 = {queue_dataIn_hi_hi_lo_hi_hi_4, queue_4_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_8 = {queue_dataIn_hi_hi_lo_hi_4, queue_dataIn_hi_hi_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_float;
  wire         queue_4_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_float, queue_4_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_4_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_4 = {queue_dataIn_hi_hi_hi_lo_hi_4, queue_4_enq_bits_decodeResult_topUop};
  wire         queue_4_enq_bits_decodeResult_orderReduce;
  wire         queue_4_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_orderReduce, queue_4_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_4_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_4 = {queue_dataIn_hi_hi_hi_hi_hi_4, queue_4_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_8 = {queue_dataIn_hi_hi_hi_hi_4, queue_dataIn_hi_hi_hi_lo_4};
  wire [16:0]  queue_dataIn_hi_hi_13 = {queue_dataIn_hi_hi_hi_8, queue_dataIn_hi_hi_lo_8};
  wire [28:0]  queue_dataIn_hi_13 = {queue_dataIn_hi_hi_13, queue_dataIn_hi_lo_13};
  wire [2:0]   queue_4_enq_bits_segment;
  wire [31:0]  queue_4_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_9 = {queue_4_enq_bits_segment, queue_4_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_9 = {queue_dataIn_lo_lo_hi_9, queue_dataIn_hi_12, queue_dataIn_lo_12};
  wire [1:0]   queue_4_enq_bits_loadStoreEEW;
  wire         queue_4_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_9 = {queue_4_enq_bits_loadStoreEEW, queue_4_enq_bits_mask};
  wire [4:0]   queue_4_enq_bits_vs2;
  wire [4:0]   queue_4_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_9 = {queue_4_enq_bits_vs2, queue_4_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_14 = {queue_dataIn_lo_hi_hi_9, queue_dataIn_lo_hi_lo_9};
  wire [80:0]  queue_dataIn_lo_14 = {queue_dataIn_lo_hi_14, queue_dataIn_lo_lo_9};
  wire         queue_4_enq_bits_lsWholeReg;
  wire [4:0]   queue_4_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_9 = {queue_4_enq_bits_lsWholeReg, queue_4_enq_bits_vs1};
  wire         queue_4_enq_bits_store;
  wire         queue_4_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_9 = {queue_4_enq_bits_store, queue_4_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_14 = {queue_dataIn_hi_lo_hi_9, queue_dataIn_hi_lo_lo_9};
  wire         queue_4_enq_bits_loadStore;
  wire         queue_4_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_9 = {queue_4_enq_bits_loadStore, queue_4_enq_bits_issueInst};
  wire [2:0]   queue_4_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_9 = {queue_4_enq_bits_instructionIndex, queue_dataIn_hi_13, queue_dataIn_lo_13};
  wire [60:0]  queue_dataIn_hi_hi_14 = {queue_dataIn_hi_hi_hi_9, queue_dataIn_hi_hi_lo_9};
  wire [68:0]  queue_dataIn_hi_14 = {queue_dataIn_hi_hi_14, queue_dataIn_hi_lo_14};
  wire [149:0] queue_dataIn_4 = {queue_dataIn_hi_14, queue_dataIn_lo_14};
  wire         queue_dataOut_4_csrInterface_vma = _queue_fifo_4_data_out[0];
  wire         queue_dataOut_4_csrInterface_vta = _queue_fifo_4_data_out[1];
  wire [1:0]   queue_dataOut_4_csrInterface_vxrm = _queue_fifo_4_data_out[3:2];
  wire [1:0]   queue_dataOut_4_csrInterface_vSew = _queue_fifo_4_data_out[5:4];
  wire [2:0]   queue_dataOut_4_csrInterface_vlmul = _queue_fifo_4_data_out[8:6];
  wire [11:0]  queue_dataOut_4_csrInterface_vStart = _queue_fifo_4_data_out[20:9];
  wire [11:0]  queue_dataOut_4_csrInterface_vl = _queue_fifo_4_data_out[32:21];
  wire [31:0]  queue_dataOut_4_readFromScalar = _queue_fifo_4_data_out[64:33];
  wire [2:0]   queue_dataOut_4_segment = _queue_fifo_4_data_out[67:65];
  wire         queue_dataOut_4_mask = _queue_fifo_4_data_out[68];
  wire [1:0]   queue_dataOut_4_loadStoreEEW = _queue_fifo_4_data_out[70:69];
  wire [4:0]   queue_dataOut_4_vd = _queue_fifo_4_data_out[75:71];
  wire [4:0]   queue_dataOut_4_vs2 = _queue_fifo_4_data_out[80:76];
  wire [4:0]   queue_dataOut_4_vs1 = _queue_fifo_4_data_out[85:81];
  wire         queue_dataOut_4_lsWholeReg = _queue_fifo_4_data_out[86];
  wire         queue_dataOut_4_special = _queue_fifo_4_data_out[87];
  wire         queue_dataOut_4_store = _queue_fifo_4_data_out[88];
  wire         queue_dataOut_4_issueInst = _queue_fifo_4_data_out[89];
  wire         queue_dataOut_4_loadStore = _queue_fifo_4_data_out[90];
  wire         queue_dataOut_4_decodeResult_logic = _queue_fifo_4_data_out[91];
  wire         queue_dataOut_4_decodeResult_adder = _queue_fifo_4_data_out[92];
  wire         queue_dataOut_4_decodeResult_shift = _queue_fifo_4_data_out[93];
  wire         queue_dataOut_4_decodeResult_multiplier = _queue_fifo_4_data_out[94];
  wire         queue_dataOut_4_decodeResult_divider = _queue_fifo_4_data_out[95];
  wire         queue_dataOut_4_decodeResult_multiCycle = _queue_fifo_4_data_out[96];
  wire         queue_dataOut_4_decodeResult_other = _queue_fifo_4_data_out[97];
  wire         queue_dataOut_4_decodeResult_unsigned0 = _queue_fifo_4_data_out[98];
  wire         queue_dataOut_4_decodeResult_unsigned1 = _queue_fifo_4_data_out[99];
  wire         queue_dataOut_4_decodeResult_itype = _queue_fifo_4_data_out[100];
  wire         queue_dataOut_4_decodeResult_nr = _queue_fifo_4_data_out[101];
  wire         queue_dataOut_4_decodeResult_red = _queue_fifo_4_data_out[102];
  wire         queue_dataOut_4_decodeResult_widenReduce = _queue_fifo_4_data_out[103];
  wire         queue_dataOut_4_decodeResult_targetRd = _queue_fifo_4_data_out[104];
  wire         queue_dataOut_4_decodeResult_slid = _queue_fifo_4_data_out[105];
  wire         queue_dataOut_4_decodeResult_gather = _queue_fifo_4_data_out[106];
  wire         queue_dataOut_4_decodeResult_gather16 = _queue_fifo_4_data_out[107];
  wire         queue_dataOut_4_decodeResult_compress = _queue_fifo_4_data_out[108];
  wire         queue_dataOut_4_decodeResult_unOrderWrite = _queue_fifo_4_data_out[109];
  wire         queue_dataOut_4_decodeResult_extend = _queue_fifo_4_data_out[110];
  wire         queue_dataOut_4_decodeResult_mv = _queue_fifo_4_data_out[111];
  wire         queue_dataOut_4_decodeResult_iota = _queue_fifo_4_data_out[112];
  wire [3:0]   queue_dataOut_4_decodeResult_uop = _queue_fifo_4_data_out[116:113];
  wire         queue_dataOut_4_decodeResult_maskLogic = _queue_fifo_4_data_out[117];
  wire         queue_dataOut_4_decodeResult_maskDestination = _queue_fifo_4_data_out[118];
  wire         queue_dataOut_4_decodeResult_maskSource = _queue_fifo_4_data_out[119];
  wire         queue_dataOut_4_decodeResult_readOnly = _queue_fifo_4_data_out[120];
  wire         queue_dataOut_4_decodeResult_vwmacc = _queue_fifo_4_data_out[121];
  wire         queue_dataOut_4_decodeResult_saturate = _queue_fifo_4_data_out[122];
  wire         queue_dataOut_4_decodeResult_special = _queue_fifo_4_data_out[123];
  wire         queue_dataOut_4_decodeResult_maskUnit = _queue_fifo_4_data_out[124];
  wire         queue_dataOut_4_decodeResult_crossWrite = _queue_fifo_4_data_out[125];
  wire         queue_dataOut_4_decodeResult_crossRead = _queue_fifo_4_data_out[126];
  wire         queue_dataOut_4_decodeResult_sWrite = _queue_fifo_4_data_out[127];
  wire         queue_dataOut_4_decodeResult_vtype = _queue_fifo_4_data_out[128];
  wire         queue_dataOut_4_decodeResult_sReadVD = _queue_fifo_4_data_out[129];
  wire         queue_dataOut_4_decodeResult_scheduler = _queue_fifo_4_data_out[130];
  wire         queue_dataOut_4_decodeResult_dontNeedExecuteInLane = _queue_fifo_4_data_out[131];
  wire         queue_dataOut_4_decodeResult_reverse = _queue_fifo_4_data_out[132];
  wire         queue_dataOut_4_decodeResult_average = _queue_fifo_4_data_out[133];
  wire         queue_dataOut_4_decodeResult_ffo = _queue_fifo_4_data_out[134];
  wire         queue_dataOut_4_decodeResult_popCount = _queue_fifo_4_data_out[135];
  wire [4:0]   queue_dataOut_4_decodeResult_topUop = _queue_fifo_4_data_out[140:136];
  wire         queue_dataOut_4_decodeResult_specialSlot = _queue_fifo_4_data_out[141];
  wire         queue_dataOut_4_decodeResult_float = _queue_fifo_4_data_out[142];
  wire [1:0]   queue_dataOut_4_decodeResult_fpExecutionType = _queue_fifo_4_data_out[144:143];
  wire         queue_dataOut_4_decodeResult_floatMul = _queue_fifo_4_data_out[145];
  wire         queue_dataOut_4_decodeResult_orderReduce = _queue_fifo_4_data_out[146];
  wire [2:0]   queue_dataOut_4_instructionIndex = _queue_fifo_4_data_out[149:147];
  wire         queue_4_enq_ready = ~_queue_fifo_4_full;
  wire         queue_4_enq_valid;
  assign queue_4_deq_valid = ~_queue_fifo_4_empty | queue_4_enq_valid;
  assign queue_4_deq_bits_instructionIndex = _queue_fifo_4_empty ? queue_4_enq_bits_instructionIndex : queue_dataOut_4_instructionIndex;
  assign queue_4_deq_bits_decodeResult_orderReduce = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_orderReduce : queue_dataOut_4_decodeResult_orderReduce;
  assign queue_4_deq_bits_decodeResult_floatMul = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_floatMul : queue_dataOut_4_decodeResult_floatMul;
  assign queue_4_deq_bits_decodeResult_fpExecutionType = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_fpExecutionType : queue_dataOut_4_decodeResult_fpExecutionType;
  assign queue_4_deq_bits_decodeResult_float = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_float : queue_dataOut_4_decodeResult_float;
  assign queue_4_deq_bits_decodeResult_specialSlot = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_specialSlot : queue_dataOut_4_decodeResult_specialSlot;
  assign queue_4_deq_bits_decodeResult_topUop = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_topUop : queue_dataOut_4_decodeResult_topUop;
  assign queue_4_deq_bits_decodeResult_popCount = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_popCount : queue_dataOut_4_decodeResult_popCount;
  assign queue_4_deq_bits_decodeResult_ffo = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_ffo : queue_dataOut_4_decodeResult_ffo;
  assign queue_4_deq_bits_decodeResult_average = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_average : queue_dataOut_4_decodeResult_average;
  assign queue_4_deq_bits_decodeResult_reverse = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_reverse : queue_dataOut_4_decodeResult_reverse;
  assign queue_4_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_4_decodeResult_dontNeedExecuteInLane;
  assign queue_4_deq_bits_decodeResult_scheduler = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_scheduler : queue_dataOut_4_decodeResult_scheduler;
  assign queue_4_deq_bits_decodeResult_sReadVD = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_sReadVD : queue_dataOut_4_decodeResult_sReadVD;
  assign queue_4_deq_bits_decodeResult_vtype = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_vtype : queue_dataOut_4_decodeResult_vtype;
  assign queue_4_deq_bits_decodeResult_sWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_sWrite : queue_dataOut_4_decodeResult_sWrite;
  assign queue_4_deq_bits_decodeResult_crossRead = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_crossRead : queue_dataOut_4_decodeResult_crossRead;
  assign queue_4_deq_bits_decodeResult_crossWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_crossWrite : queue_dataOut_4_decodeResult_crossWrite;
  assign queue_4_deq_bits_decodeResult_maskUnit = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskUnit : queue_dataOut_4_decodeResult_maskUnit;
  assign queue_4_deq_bits_decodeResult_special = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_special : queue_dataOut_4_decodeResult_special;
  assign queue_4_deq_bits_decodeResult_saturate = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_saturate : queue_dataOut_4_decodeResult_saturate;
  assign queue_4_deq_bits_decodeResult_vwmacc = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_vwmacc : queue_dataOut_4_decodeResult_vwmacc;
  assign queue_4_deq_bits_decodeResult_readOnly = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_readOnly : queue_dataOut_4_decodeResult_readOnly;
  assign queue_4_deq_bits_decodeResult_maskSource = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskSource : queue_dataOut_4_decodeResult_maskSource;
  assign queue_4_deq_bits_decodeResult_maskDestination = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskDestination : queue_dataOut_4_decodeResult_maskDestination;
  assign queue_4_deq_bits_decodeResult_maskLogic = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskLogic : queue_dataOut_4_decodeResult_maskLogic;
  assign queue_4_deq_bits_decodeResult_uop = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_uop : queue_dataOut_4_decodeResult_uop;
  assign queue_4_deq_bits_decodeResult_iota = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_iota : queue_dataOut_4_decodeResult_iota;
  assign queue_4_deq_bits_decodeResult_mv = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_mv : queue_dataOut_4_decodeResult_mv;
  assign queue_4_deq_bits_decodeResult_extend = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_extend : queue_dataOut_4_decodeResult_extend;
  assign queue_4_deq_bits_decodeResult_unOrderWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unOrderWrite : queue_dataOut_4_decodeResult_unOrderWrite;
  assign queue_4_deq_bits_decodeResult_compress = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_compress : queue_dataOut_4_decodeResult_compress;
  assign queue_4_deq_bits_decodeResult_gather16 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_gather16 : queue_dataOut_4_decodeResult_gather16;
  assign queue_4_deq_bits_decodeResult_gather = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_gather : queue_dataOut_4_decodeResult_gather;
  assign queue_4_deq_bits_decodeResult_slid = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_slid : queue_dataOut_4_decodeResult_slid;
  assign queue_4_deq_bits_decodeResult_targetRd = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_targetRd : queue_dataOut_4_decodeResult_targetRd;
  assign queue_4_deq_bits_decodeResult_widenReduce = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_widenReduce : queue_dataOut_4_decodeResult_widenReduce;
  assign queue_4_deq_bits_decodeResult_red = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_red : queue_dataOut_4_decodeResult_red;
  assign queue_4_deq_bits_decodeResult_nr = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_nr : queue_dataOut_4_decodeResult_nr;
  assign queue_4_deq_bits_decodeResult_itype = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_itype : queue_dataOut_4_decodeResult_itype;
  assign queue_4_deq_bits_decodeResult_unsigned1 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unsigned1 : queue_dataOut_4_decodeResult_unsigned1;
  assign queue_4_deq_bits_decodeResult_unsigned0 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unsigned0 : queue_dataOut_4_decodeResult_unsigned0;
  assign queue_4_deq_bits_decodeResult_other = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_other : queue_dataOut_4_decodeResult_other;
  assign queue_4_deq_bits_decodeResult_multiCycle = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_multiCycle : queue_dataOut_4_decodeResult_multiCycle;
  assign queue_4_deq_bits_decodeResult_divider = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_divider : queue_dataOut_4_decodeResult_divider;
  assign queue_4_deq_bits_decodeResult_multiplier = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_multiplier : queue_dataOut_4_decodeResult_multiplier;
  assign queue_4_deq_bits_decodeResult_shift = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_shift : queue_dataOut_4_decodeResult_shift;
  assign queue_4_deq_bits_decodeResult_adder = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_adder : queue_dataOut_4_decodeResult_adder;
  assign queue_4_deq_bits_decodeResult_logic = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_logic : queue_dataOut_4_decodeResult_logic;
  assign queue_4_deq_bits_loadStore = _queue_fifo_4_empty ? queue_4_enq_bits_loadStore : queue_dataOut_4_loadStore;
  assign queue_4_deq_bits_issueInst = _queue_fifo_4_empty ? queue_4_enq_bits_issueInst : queue_dataOut_4_issueInst;
  assign queue_4_deq_bits_store = _queue_fifo_4_empty ? queue_4_enq_bits_store : queue_dataOut_4_store;
  assign queue_4_deq_bits_special = _queue_fifo_4_empty ? queue_4_enq_bits_special : queue_dataOut_4_special;
  assign queue_4_deq_bits_lsWholeReg = _queue_fifo_4_empty ? queue_4_enq_bits_lsWholeReg : queue_dataOut_4_lsWholeReg;
  assign queue_4_deq_bits_vs1 = _queue_fifo_4_empty ? queue_4_enq_bits_vs1 : queue_dataOut_4_vs1;
  assign queue_4_deq_bits_vs2 = _queue_fifo_4_empty ? queue_4_enq_bits_vs2 : queue_dataOut_4_vs2;
  assign queue_4_deq_bits_vd = _queue_fifo_4_empty ? queue_4_enq_bits_vd : queue_dataOut_4_vd;
  assign queue_4_deq_bits_loadStoreEEW = _queue_fifo_4_empty ? queue_4_enq_bits_loadStoreEEW : queue_dataOut_4_loadStoreEEW;
  assign queue_4_deq_bits_mask = _queue_fifo_4_empty ? queue_4_enq_bits_mask : queue_dataOut_4_mask;
  assign queue_4_deq_bits_segment = _queue_fifo_4_empty ? queue_4_enq_bits_segment : queue_dataOut_4_segment;
  assign queue_4_deq_bits_readFromScalar = _queue_fifo_4_empty ? queue_4_enq_bits_readFromScalar : queue_dataOut_4_readFromScalar;
  assign queue_4_deq_bits_csrInterface_vl = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vl : queue_dataOut_4_csrInterface_vl;
  assign queue_4_deq_bits_csrInterface_vStart = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vStart : queue_dataOut_4_csrInterface_vStart;
  assign queue_4_deq_bits_csrInterface_vlmul = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vlmul : queue_dataOut_4_csrInterface_vlmul;
  assign queue_4_deq_bits_csrInterface_vSew = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vSew : queue_dataOut_4_csrInterface_vSew;
  assign queue_4_deq_bits_csrInterface_vxrm = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vxrm : queue_dataOut_4_csrInterface_vxrm;
  assign queue_4_deq_bits_csrInterface_vta = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vta : queue_dataOut_4_csrInterface_vta;
  assign queue_4_deq_bits_csrInterface_vma = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vma : queue_dataOut_4_csrInterface_vma;
  wire         laneVec_4_laneRequest_bits_issueInst = laneRequestSinkWire_4_ready & laneRequestSinkWire_4_valid;
  reg          releasePipe_pipe_v_4;
  wire         releasePipe_pipe_out_4_valid = releasePipe_pipe_v_4;
  wire         laneRequestSourceWire_4_ready;
  wire         validSource_4_valid = laneRequestSourceWire_4_ready & laneRequestSourceWire_4_valid;
  reg  [2:0]   tokenCheck_counter_4;
  wire [2:0]   tokenCheck_counterChange_4 = validSource_4_valid ? 3'h1 : 3'h7;
  assign tokenCheck_4 = ~(tokenCheck_counter_4[2]);
  assign laneRequestSourceWire_4_ready = tokenCheck_4;
  assign queue_4_enq_valid = validSink_4_valid;
  assign queue_4_enq_bits_instructionIndex = validSink_4_bits_instructionIndex;
  assign queue_4_enq_bits_decodeResult_orderReduce = validSink_4_bits_decodeResult_orderReduce;
  assign queue_4_enq_bits_decodeResult_floatMul = validSink_4_bits_decodeResult_floatMul;
  assign queue_4_enq_bits_decodeResult_fpExecutionType = validSink_4_bits_decodeResult_fpExecutionType;
  assign queue_4_enq_bits_decodeResult_float = validSink_4_bits_decodeResult_float;
  assign queue_4_enq_bits_decodeResult_specialSlot = validSink_4_bits_decodeResult_specialSlot;
  assign queue_4_enq_bits_decodeResult_topUop = validSink_4_bits_decodeResult_topUop;
  assign queue_4_enq_bits_decodeResult_popCount = validSink_4_bits_decodeResult_popCount;
  assign queue_4_enq_bits_decodeResult_ffo = validSink_4_bits_decodeResult_ffo;
  assign queue_4_enq_bits_decodeResult_average = validSink_4_bits_decodeResult_average;
  assign queue_4_enq_bits_decodeResult_reverse = validSink_4_bits_decodeResult_reverse;
  assign queue_4_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_4_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_4_enq_bits_decodeResult_scheduler = validSink_4_bits_decodeResult_scheduler;
  assign queue_4_enq_bits_decodeResult_sReadVD = validSink_4_bits_decodeResult_sReadVD;
  assign queue_4_enq_bits_decodeResult_vtype = validSink_4_bits_decodeResult_vtype;
  assign queue_4_enq_bits_decodeResult_sWrite = validSink_4_bits_decodeResult_sWrite;
  assign queue_4_enq_bits_decodeResult_crossRead = validSink_4_bits_decodeResult_crossRead;
  assign queue_4_enq_bits_decodeResult_crossWrite = validSink_4_bits_decodeResult_crossWrite;
  assign queue_4_enq_bits_decodeResult_maskUnit = validSink_4_bits_decodeResult_maskUnit;
  assign queue_4_enq_bits_decodeResult_special = validSink_4_bits_decodeResult_special;
  assign queue_4_enq_bits_decodeResult_saturate = validSink_4_bits_decodeResult_saturate;
  assign queue_4_enq_bits_decodeResult_vwmacc = validSink_4_bits_decodeResult_vwmacc;
  assign queue_4_enq_bits_decodeResult_readOnly = validSink_4_bits_decodeResult_readOnly;
  assign queue_4_enq_bits_decodeResult_maskSource = validSink_4_bits_decodeResult_maskSource;
  assign queue_4_enq_bits_decodeResult_maskDestination = validSink_4_bits_decodeResult_maskDestination;
  assign queue_4_enq_bits_decodeResult_maskLogic = validSink_4_bits_decodeResult_maskLogic;
  assign queue_4_enq_bits_decodeResult_uop = validSink_4_bits_decodeResult_uop;
  assign queue_4_enq_bits_decodeResult_iota = validSink_4_bits_decodeResult_iota;
  assign queue_4_enq_bits_decodeResult_mv = validSink_4_bits_decodeResult_mv;
  assign queue_4_enq_bits_decodeResult_extend = validSink_4_bits_decodeResult_extend;
  assign queue_4_enq_bits_decodeResult_unOrderWrite = validSink_4_bits_decodeResult_unOrderWrite;
  assign queue_4_enq_bits_decodeResult_compress = validSink_4_bits_decodeResult_compress;
  assign queue_4_enq_bits_decodeResult_gather16 = validSink_4_bits_decodeResult_gather16;
  assign queue_4_enq_bits_decodeResult_gather = validSink_4_bits_decodeResult_gather;
  assign queue_4_enq_bits_decodeResult_slid = validSink_4_bits_decodeResult_slid;
  assign queue_4_enq_bits_decodeResult_targetRd = validSink_4_bits_decodeResult_targetRd;
  assign queue_4_enq_bits_decodeResult_widenReduce = validSink_4_bits_decodeResult_widenReduce;
  assign queue_4_enq_bits_decodeResult_red = validSink_4_bits_decodeResult_red;
  assign queue_4_enq_bits_decodeResult_nr = validSink_4_bits_decodeResult_nr;
  assign queue_4_enq_bits_decodeResult_itype = validSink_4_bits_decodeResult_itype;
  assign queue_4_enq_bits_decodeResult_unsigned1 = validSink_4_bits_decodeResult_unsigned1;
  assign queue_4_enq_bits_decodeResult_unsigned0 = validSink_4_bits_decodeResult_unsigned0;
  assign queue_4_enq_bits_decodeResult_other = validSink_4_bits_decodeResult_other;
  assign queue_4_enq_bits_decodeResult_multiCycle = validSink_4_bits_decodeResult_multiCycle;
  assign queue_4_enq_bits_decodeResult_divider = validSink_4_bits_decodeResult_divider;
  assign queue_4_enq_bits_decodeResult_multiplier = validSink_4_bits_decodeResult_multiplier;
  assign queue_4_enq_bits_decodeResult_shift = validSink_4_bits_decodeResult_shift;
  assign queue_4_enq_bits_decodeResult_adder = validSink_4_bits_decodeResult_adder;
  assign queue_4_enq_bits_decodeResult_logic = validSink_4_bits_decodeResult_logic;
  assign queue_4_enq_bits_loadStore = validSink_4_bits_loadStore;
  assign queue_4_enq_bits_issueInst = validSink_4_bits_issueInst;
  assign queue_4_enq_bits_store = validSink_4_bits_store;
  assign queue_4_enq_bits_special = validSink_4_bits_special;
  assign queue_4_enq_bits_lsWholeReg = validSink_4_bits_lsWholeReg;
  assign queue_4_enq_bits_vs1 = validSink_4_bits_vs1;
  assign queue_4_enq_bits_vs2 = validSink_4_bits_vs2;
  assign queue_4_enq_bits_vd = validSink_4_bits_vd;
  assign queue_4_enq_bits_loadStoreEEW = validSink_4_bits_loadStoreEEW;
  assign queue_4_enq_bits_mask = validSink_4_bits_mask;
  assign queue_4_enq_bits_segment = validSink_4_bits_segment;
  assign queue_4_enq_bits_readFromScalar = validSink_4_bits_readFromScalar;
  assign queue_4_enq_bits_csrInterface_vl = validSink_4_bits_csrInterface_vl;
  assign queue_4_enq_bits_csrInterface_vStart = validSink_4_bits_csrInterface_vStart;
  assign queue_4_enq_bits_csrInterface_vlmul = validSink_4_bits_csrInterface_vlmul;
  assign queue_4_enq_bits_csrInterface_vSew = validSink_4_bits_csrInterface_vSew;
  assign queue_4_enq_bits_csrInterface_vxrm = validSink_4_bits_csrInterface_vxrm;
  assign queue_4_enq_bits_csrInterface_vta = validSink_4_bits_csrInterface_vta;
  assign queue_4_enq_bits_csrInterface_vma = validSink_4_bits_csrInterface_vma;
  reg          shifterReg_4_0_valid;
  assign validSink_4_valid = shifterReg_4_0_valid;
  reg  [2:0]   shifterReg_4_0_bits_instructionIndex;
  assign validSink_4_bits_instructionIndex = shifterReg_4_0_bits_instructionIndex;
  reg          shifterReg_4_0_bits_decodeResult_orderReduce;
  assign validSink_4_bits_decodeResult_orderReduce = shifterReg_4_0_bits_decodeResult_orderReduce;
  reg          shifterReg_4_0_bits_decodeResult_floatMul;
  assign validSink_4_bits_decodeResult_floatMul = shifterReg_4_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_4_0_bits_decodeResult_fpExecutionType;
  assign validSink_4_bits_decodeResult_fpExecutionType = shifterReg_4_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_4_0_bits_decodeResult_float;
  assign validSink_4_bits_decodeResult_float = shifterReg_4_0_bits_decodeResult_float;
  reg          shifterReg_4_0_bits_decodeResult_specialSlot;
  assign validSink_4_bits_decodeResult_specialSlot = shifterReg_4_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_4_0_bits_decodeResult_topUop;
  assign validSink_4_bits_decodeResult_topUop = shifterReg_4_0_bits_decodeResult_topUop;
  reg          shifterReg_4_0_bits_decodeResult_popCount;
  assign validSink_4_bits_decodeResult_popCount = shifterReg_4_0_bits_decodeResult_popCount;
  reg          shifterReg_4_0_bits_decodeResult_ffo;
  assign validSink_4_bits_decodeResult_ffo = shifterReg_4_0_bits_decodeResult_ffo;
  reg          shifterReg_4_0_bits_decodeResult_average;
  assign validSink_4_bits_decodeResult_average = shifterReg_4_0_bits_decodeResult_average;
  reg          shifterReg_4_0_bits_decodeResult_reverse;
  assign validSink_4_bits_decodeResult_reverse = shifterReg_4_0_bits_decodeResult_reverse;
  reg          shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_4_bits_decodeResult_dontNeedExecuteInLane = shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_4_0_bits_decodeResult_scheduler;
  assign validSink_4_bits_decodeResult_scheduler = shifterReg_4_0_bits_decodeResult_scheduler;
  reg          shifterReg_4_0_bits_decodeResult_sReadVD;
  assign validSink_4_bits_decodeResult_sReadVD = shifterReg_4_0_bits_decodeResult_sReadVD;
  reg          shifterReg_4_0_bits_decodeResult_vtype;
  assign validSink_4_bits_decodeResult_vtype = shifterReg_4_0_bits_decodeResult_vtype;
  reg          shifterReg_4_0_bits_decodeResult_sWrite;
  assign validSink_4_bits_decodeResult_sWrite = shifterReg_4_0_bits_decodeResult_sWrite;
  reg          shifterReg_4_0_bits_decodeResult_crossRead;
  assign validSink_4_bits_decodeResult_crossRead = shifterReg_4_0_bits_decodeResult_crossRead;
  reg          shifterReg_4_0_bits_decodeResult_crossWrite;
  assign validSink_4_bits_decodeResult_crossWrite = shifterReg_4_0_bits_decodeResult_crossWrite;
  reg          shifterReg_4_0_bits_decodeResult_maskUnit;
  assign validSink_4_bits_decodeResult_maskUnit = shifterReg_4_0_bits_decodeResult_maskUnit;
  reg          shifterReg_4_0_bits_decodeResult_special;
  assign validSink_4_bits_decodeResult_special = shifterReg_4_0_bits_decodeResult_special;
  reg          shifterReg_4_0_bits_decodeResult_saturate;
  assign validSink_4_bits_decodeResult_saturate = shifterReg_4_0_bits_decodeResult_saturate;
  reg          shifterReg_4_0_bits_decodeResult_vwmacc;
  assign validSink_4_bits_decodeResult_vwmacc = shifterReg_4_0_bits_decodeResult_vwmacc;
  reg          shifterReg_4_0_bits_decodeResult_readOnly;
  assign validSink_4_bits_decodeResult_readOnly = shifterReg_4_0_bits_decodeResult_readOnly;
  reg          shifterReg_4_0_bits_decodeResult_maskSource;
  assign validSink_4_bits_decodeResult_maskSource = shifterReg_4_0_bits_decodeResult_maskSource;
  reg          shifterReg_4_0_bits_decodeResult_maskDestination;
  assign validSink_4_bits_decodeResult_maskDestination = shifterReg_4_0_bits_decodeResult_maskDestination;
  reg          shifterReg_4_0_bits_decodeResult_maskLogic;
  assign validSink_4_bits_decodeResult_maskLogic = shifterReg_4_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_4_0_bits_decodeResult_uop;
  assign validSink_4_bits_decodeResult_uop = shifterReg_4_0_bits_decodeResult_uop;
  reg          shifterReg_4_0_bits_decodeResult_iota;
  assign validSink_4_bits_decodeResult_iota = shifterReg_4_0_bits_decodeResult_iota;
  reg          shifterReg_4_0_bits_decodeResult_mv;
  assign validSink_4_bits_decodeResult_mv = shifterReg_4_0_bits_decodeResult_mv;
  reg          shifterReg_4_0_bits_decodeResult_extend;
  assign validSink_4_bits_decodeResult_extend = shifterReg_4_0_bits_decodeResult_extend;
  reg          shifterReg_4_0_bits_decodeResult_unOrderWrite;
  assign validSink_4_bits_decodeResult_unOrderWrite = shifterReg_4_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_4_0_bits_decodeResult_compress;
  assign validSink_4_bits_decodeResult_compress = shifterReg_4_0_bits_decodeResult_compress;
  reg          shifterReg_4_0_bits_decodeResult_gather16;
  assign validSink_4_bits_decodeResult_gather16 = shifterReg_4_0_bits_decodeResult_gather16;
  reg          shifterReg_4_0_bits_decodeResult_gather;
  assign validSink_4_bits_decodeResult_gather = shifterReg_4_0_bits_decodeResult_gather;
  reg          shifterReg_4_0_bits_decodeResult_slid;
  assign validSink_4_bits_decodeResult_slid = shifterReg_4_0_bits_decodeResult_slid;
  reg          shifterReg_4_0_bits_decodeResult_targetRd;
  assign validSink_4_bits_decodeResult_targetRd = shifterReg_4_0_bits_decodeResult_targetRd;
  reg          shifterReg_4_0_bits_decodeResult_widenReduce;
  assign validSink_4_bits_decodeResult_widenReduce = shifterReg_4_0_bits_decodeResult_widenReduce;
  reg          shifterReg_4_0_bits_decodeResult_red;
  assign validSink_4_bits_decodeResult_red = shifterReg_4_0_bits_decodeResult_red;
  reg          shifterReg_4_0_bits_decodeResult_nr;
  assign validSink_4_bits_decodeResult_nr = shifterReg_4_0_bits_decodeResult_nr;
  reg          shifterReg_4_0_bits_decodeResult_itype;
  assign validSink_4_bits_decodeResult_itype = shifterReg_4_0_bits_decodeResult_itype;
  reg          shifterReg_4_0_bits_decodeResult_unsigned1;
  assign validSink_4_bits_decodeResult_unsigned1 = shifterReg_4_0_bits_decodeResult_unsigned1;
  reg          shifterReg_4_0_bits_decodeResult_unsigned0;
  assign validSink_4_bits_decodeResult_unsigned0 = shifterReg_4_0_bits_decodeResult_unsigned0;
  reg          shifterReg_4_0_bits_decodeResult_other;
  assign validSink_4_bits_decodeResult_other = shifterReg_4_0_bits_decodeResult_other;
  reg          shifterReg_4_0_bits_decodeResult_multiCycle;
  assign validSink_4_bits_decodeResult_multiCycle = shifterReg_4_0_bits_decodeResult_multiCycle;
  reg          shifterReg_4_0_bits_decodeResult_divider;
  assign validSink_4_bits_decodeResult_divider = shifterReg_4_0_bits_decodeResult_divider;
  reg          shifterReg_4_0_bits_decodeResult_multiplier;
  assign validSink_4_bits_decodeResult_multiplier = shifterReg_4_0_bits_decodeResult_multiplier;
  reg          shifterReg_4_0_bits_decodeResult_shift;
  assign validSink_4_bits_decodeResult_shift = shifterReg_4_0_bits_decodeResult_shift;
  reg          shifterReg_4_0_bits_decodeResult_adder;
  assign validSink_4_bits_decodeResult_adder = shifterReg_4_0_bits_decodeResult_adder;
  reg          shifterReg_4_0_bits_decodeResult_logic;
  assign validSink_4_bits_decodeResult_logic = shifterReg_4_0_bits_decodeResult_logic;
  reg          shifterReg_4_0_bits_loadStore;
  assign validSink_4_bits_loadStore = shifterReg_4_0_bits_loadStore;
  reg          shifterReg_4_0_bits_issueInst;
  assign validSink_4_bits_issueInst = shifterReg_4_0_bits_issueInst;
  reg          shifterReg_4_0_bits_store;
  assign validSink_4_bits_store = shifterReg_4_0_bits_store;
  reg          shifterReg_4_0_bits_special;
  assign validSink_4_bits_special = shifterReg_4_0_bits_special;
  reg          shifterReg_4_0_bits_lsWholeReg;
  assign validSink_4_bits_lsWholeReg = shifterReg_4_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_4_0_bits_vs1;
  assign validSink_4_bits_vs1 = shifterReg_4_0_bits_vs1;
  reg  [4:0]   shifterReg_4_0_bits_vs2;
  assign validSink_4_bits_vs2 = shifterReg_4_0_bits_vs2;
  reg  [4:0]   shifterReg_4_0_bits_vd;
  assign validSink_4_bits_vd = shifterReg_4_0_bits_vd;
  reg  [1:0]   shifterReg_4_0_bits_loadStoreEEW;
  assign validSink_4_bits_loadStoreEEW = shifterReg_4_0_bits_loadStoreEEW;
  reg          shifterReg_4_0_bits_mask;
  assign validSink_4_bits_mask = shifterReg_4_0_bits_mask;
  reg  [2:0]   shifterReg_4_0_bits_segment;
  assign validSink_4_bits_segment = shifterReg_4_0_bits_segment;
  reg  [31:0]  shifterReg_4_0_bits_readFromScalar;
  assign validSink_4_bits_readFromScalar = shifterReg_4_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_4_0_bits_csrInterface_vl;
  assign validSink_4_bits_csrInterface_vl = shifterReg_4_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_4_0_bits_csrInterface_vStart;
  assign validSink_4_bits_csrInterface_vStart = shifterReg_4_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_4_0_bits_csrInterface_vlmul;
  assign validSink_4_bits_csrInterface_vlmul = shifterReg_4_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_4_0_bits_csrInterface_vSew;
  assign validSink_4_bits_csrInterface_vSew = shifterReg_4_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_4_0_bits_csrInterface_vxrm;
  assign validSink_4_bits_csrInterface_vxrm = shifterReg_4_0_bits_csrInterface_vxrm;
  reg          shifterReg_4_0_bits_csrInterface_vta;
  assign validSink_4_bits_csrInterface_vta = shifterReg_4_0_bits_csrInterface_vta;
  reg          shifterReg_4_0_bits_csrInterface_vma;
  assign validSink_4_bits_csrInterface_vma = shifterReg_4_0_bits_csrInterface_vma;
  wire         shifterValid_4 = shifterReg_4_0_valid | validSource_4_valid;
  wire         validSink_5_valid;
  wire [2:0]   validSink_5_bits_instructionIndex;
  wire         validSink_5_bits_decodeResult_orderReduce;
  wire         validSink_5_bits_decodeResult_floatMul;
  wire [1:0]   validSink_5_bits_decodeResult_fpExecutionType;
  wire         validSink_5_bits_decodeResult_float;
  wire         validSink_5_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_5_bits_decodeResult_topUop;
  wire         validSink_5_bits_decodeResult_popCount;
  wire         validSink_5_bits_decodeResult_ffo;
  wire         validSink_5_bits_decodeResult_average;
  wire         validSink_5_bits_decodeResult_reverse;
  wire         validSink_5_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_5_bits_decodeResult_scheduler;
  wire         validSink_5_bits_decodeResult_sReadVD;
  wire         validSink_5_bits_decodeResult_vtype;
  wire         validSink_5_bits_decodeResult_sWrite;
  wire         validSink_5_bits_decodeResult_crossRead;
  wire         validSink_5_bits_decodeResult_crossWrite;
  wire         validSink_5_bits_decodeResult_maskUnit;
  wire         validSink_5_bits_decodeResult_special;
  wire         validSink_5_bits_decodeResult_saturate;
  wire         validSink_5_bits_decodeResult_vwmacc;
  wire         validSink_5_bits_decodeResult_readOnly;
  wire         validSink_5_bits_decodeResult_maskSource;
  wire         validSink_5_bits_decodeResult_maskDestination;
  wire         validSink_5_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_5_bits_decodeResult_uop;
  wire         validSink_5_bits_decodeResult_iota;
  wire         validSink_5_bits_decodeResult_mv;
  wire         validSink_5_bits_decodeResult_extend;
  wire         validSink_5_bits_decodeResult_unOrderWrite;
  wire         validSink_5_bits_decodeResult_compress;
  wire         validSink_5_bits_decodeResult_gather16;
  wire         validSink_5_bits_decodeResult_gather;
  wire         validSink_5_bits_decodeResult_slid;
  wire         validSink_5_bits_decodeResult_targetRd;
  wire         validSink_5_bits_decodeResult_widenReduce;
  wire         validSink_5_bits_decodeResult_red;
  wire         validSink_5_bits_decodeResult_nr;
  wire         validSink_5_bits_decodeResult_itype;
  wire         validSink_5_bits_decodeResult_unsigned1;
  wire         validSink_5_bits_decodeResult_unsigned0;
  wire         validSink_5_bits_decodeResult_other;
  wire         validSink_5_bits_decodeResult_multiCycle;
  wire         validSink_5_bits_decodeResult_divider;
  wire         validSink_5_bits_decodeResult_multiplier;
  wire         validSink_5_bits_decodeResult_shift;
  wire         validSink_5_bits_decodeResult_adder;
  wire         validSink_5_bits_decodeResult_logic;
  wire         validSink_5_bits_loadStore;
  wire         validSink_5_bits_issueInst;
  wire         validSink_5_bits_store;
  wire         validSink_5_bits_special;
  wire         validSink_5_bits_lsWholeReg;
  wire [4:0]   validSink_5_bits_vs1;
  wire [4:0]   validSink_5_bits_vs2;
  wire [4:0]   validSink_5_bits_vd;
  wire [1:0]   validSink_5_bits_loadStoreEEW;
  wire         validSink_5_bits_mask;
  wire [2:0]   validSink_5_bits_segment;
  wire [31:0]  validSink_5_bits_readFromScalar;
  wire [11:0]  validSink_5_bits_csrInterface_vl;
  wire [11:0]  validSink_5_bits_csrInterface_vStart;
  wire [2:0]   validSink_5_bits_csrInterface_vlmul;
  wire [1:0]   validSink_5_bits_csrInterface_vSew;
  wire [1:0]   validSink_5_bits_csrInterface_vxrm;
  wire         validSink_5_bits_csrInterface_vta;
  wire         validSink_5_bits_csrInterface_vma;
  wire         laneRequestSinkWire_5_valid = queue_5_deq_valid;
  wire [2:0]   laneRequestSinkWire_5_bits_instructionIndex = queue_5_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_5_bits_decodeResult_orderReduce = queue_5_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_5_bits_decodeResult_floatMul = queue_5_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_5_bits_decodeResult_fpExecutionType = queue_5_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_5_bits_decodeResult_float = queue_5_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_5_bits_decodeResult_specialSlot = queue_5_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_5_bits_decodeResult_topUop = queue_5_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_5_bits_decodeResult_popCount = queue_5_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_5_bits_decodeResult_ffo = queue_5_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_5_bits_decodeResult_average = queue_5_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_5_bits_decodeResult_reverse = queue_5_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_5_bits_decodeResult_dontNeedExecuteInLane = queue_5_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_5_bits_decodeResult_scheduler = queue_5_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_5_bits_decodeResult_sReadVD = queue_5_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_5_bits_decodeResult_vtype = queue_5_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_5_bits_decodeResult_sWrite = queue_5_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_crossRead = queue_5_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_5_bits_decodeResult_crossWrite = queue_5_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskUnit = queue_5_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_5_bits_decodeResult_special = queue_5_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_5_bits_decodeResult_saturate = queue_5_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_5_bits_decodeResult_vwmacc = queue_5_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_5_bits_decodeResult_readOnly = queue_5_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskSource = queue_5_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskDestination = queue_5_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskLogic = queue_5_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_5_bits_decodeResult_uop = queue_5_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_5_bits_decodeResult_iota = queue_5_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_5_bits_decodeResult_mv = queue_5_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_5_bits_decodeResult_extend = queue_5_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_5_bits_decodeResult_unOrderWrite = queue_5_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_compress = queue_5_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_5_bits_decodeResult_gather16 = queue_5_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_5_bits_decodeResult_gather = queue_5_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_5_bits_decodeResult_slid = queue_5_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_5_bits_decodeResult_targetRd = queue_5_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_5_bits_decodeResult_widenReduce = queue_5_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_5_bits_decodeResult_red = queue_5_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_5_bits_decodeResult_nr = queue_5_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_5_bits_decodeResult_itype = queue_5_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_5_bits_decodeResult_unsigned1 = queue_5_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_5_bits_decodeResult_unsigned0 = queue_5_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_5_bits_decodeResult_other = queue_5_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_5_bits_decodeResult_multiCycle = queue_5_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_5_bits_decodeResult_divider = queue_5_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_5_bits_decodeResult_multiplier = queue_5_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_5_bits_decodeResult_shift = queue_5_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_5_bits_decodeResult_adder = queue_5_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_5_bits_decodeResult_logic = queue_5_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_5_bits_loadStore = queue_5_deq_bits_loadStore;
  wire         laneRequestSinkWire_5_bits_issueInst = queue_5_deq_bits_issueInst;
  wire         laneRequestSinkWire_5_bits_store = queue_5_deq_bits_store;
  wire         laneRequestSinkWire_5_bits_special = queue_5_deq_bits_special;
  wire         laneRequestSinkWire_5_bits_lsWholeReg = queue_5_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_5_bits_vs1 = queue_5_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_5_bits_vs2 = queue_5_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_5_bits_vd = queue_5_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_5_bits_loadStoreEEW = queue_5_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_5_bits_mask = queue_5_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_5_bits_segment = queue_5_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_5_bits_readFromScalar = queue_5_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_5_bits_csrInterface_vl = queue_5_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_5_bits_csrInterface_vStart = queue_5_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_5_bits_csrInterface_vlmul = queue_5_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_5_bits_csrInterface_vSew = queue_5_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_5_bits_csrInterface_vxrm = queue_5_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_5_bits_csrInterface_vta = queue_5_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_5_bits_csrInterface_vma = queue_5_deq_bits_csrInterface_vma;
  wire [1:0]   queue_5_enq_bits_csrInterface_vxrm;
  wire         queue_5_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_15 = {queue_5_enq_bits_csrInterface_vxrm, queue_5_enq_bits_csrInterface_vta};
  wire         queue_5_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_15 = {queue_dataIn_lo_hi_15, queue_5_enq_bits_csrInterface_vma};
  wire [2:0]   queue_5_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_5_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_15 = {queue_5_enq_bits_csrInterface_vlmul, queue_5_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_5_enq_bits_csrInterface_vl;
  wire [11:0]  queue_5_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_15 = {queue_5_enq_bits_csrInterface_vl, queue_5_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_15 = {queue_dataIn_hi_hi_15, queue_dataIn_hi_lo_15};
  wire         queue_5_enq_bits_decodeResult_shift;
  wire         queue_5_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_5 = {queue_5_enq_bits_decodeResult_shift, queue_5_enq_bits_decodeResult_adder};
  wire         queue_5_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_5 = {queue_dataIn_lo_lo_lo_lo_hi_5, queue_5_enq_bits_decodeResult_logic};
  wire         queue_5_enq_bits_decodeResult_multiCycle;
  wire         queue_5_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_multiCycle, queue_5_enq_bits_decodeResult_divider};
  wire         queue_5_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_5 = {queue_dataIn_lo_lo_lo_hi_hi_5, queue_5_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_5 = {queue_dataIn_lo_lo_lo_hi_5, queue_dataIn_lo_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_unsigned1;
  wire         queue_5_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_unsigned1, queue_5_enq_bits_decodeResult_unsigned0};
  wire         queue_5_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_5 = {queue_dataIn_lo_lo_hi_lo_hi_5, queue_5_enq_bits_decodeResult_other};
  wire         queue_5_enq_bits_decodeResult_red;
  wire         queue_5_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_red, queue_5_enq_bits_decodeResult_nr};
  wire         queue_5_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_5 = {queue_dataIn_lo_lo_hi_hi_hi_5, queue_5_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_10 = {queue_dataIn_lo_lo_hi_hi_5, queue_dataIn_lo_lo_hi_lo_5};
  wire [11:0]  queue_dataIn_lo_lo_10 = {queue_dataIn_lo_lo_hi_10, queue_dataIn_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_slid;
  wire         queue_5_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_5 = {queue_5_enq_bits_decodeResult_slid, queue_5_enq_bits_decodeResult_targetRd};
  wire         queue_5_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_5 = {queue_dataIn_lo_hi_lo_lo_hi_5, queue_5_enq_bits_decodeResult_widenReduce};
  wire         queue_5_enq_bits_decodeResult_compress;
  wire         queue_5_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_compress, queue_5_enq_bits_decodeResult_gather16};
  wire         queue_5_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_5 = {queue_dataIn_lo_hi_lo_hi_hi_5, queue_5_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_10 = {queue_dataIn_lo_hi_lo_hi_5, queue_dataIn_lo_hi_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_mv;
  wire         queue_5_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_mv, queue_5_enq_bits_decodeResult_extend};
  wire         queue_5_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_5 = {queue_dataIn_lo_hi_hi_lo_hi_5, queue_5_enq_bits_decodeResult_unOrderWrite};
  wire         queue_5_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_5_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_maskLogic, queue_5_enq_bits_decodeResult_uop};
  wire         queue_5_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_5 = {queue_dataIn_lo_hi_hi_hi_hi_5, queue_5_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_10 = {queue_dataIn_lo_hi_hi_hi_5, queue_dataIn_lo_hi_hi_lo_5};
  wire [14:0]  queue_dataIn_lo_hi_16 = {queue_dataIn_lo_hi_hi_10, queue_dataIn_lo_hi_lo_10};
  wire [26:0]  queue_dataIn_lo_16 = {queue_dataIn_lo_hi_16, queue_dataIn_lo_lo_10};
  wire         queue_5_enq_bits_decodeResult_readOnly;
  wire         queue_5_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_5 = {queue_5_enq_bits_decodeResult_readOnly, queue_5_enq_bits_decodeResult_maskSource};
  wire         queue_5_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_5 = {queue_dataIn_hi_lo_lo_lo_hi_5, queue_5_enq_bits_decodeResult_maskDestination};
  wire         queue_5_enq_bits_decodeResult_special;
  wire         queue_5_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_special, queue_5_enq_bits_decodeResult_saturate};
  wire         queue_5_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_5 = {queue_dataIn_hi_lo_lo_hi_hi_5, queue_5_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_10 = {queue_dataIn_hi_lo_lo_hi_5, queue_dataIn_hi_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_crossRead;
  wire         queue_5_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_crossRead, queue_5_enq_bits_decodeResult_crossWrite};
  wire         queue_5_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_5 = {queue_dataIn_hi_lo_hi_lo_hi_5, queue_5_enq_bits_decodeResult_maskUnit};
  wire         queue_5_enq_bits_decodeResult_sReadVD;
  wire         queue_5_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_sReadVD, queue_5_enq_bits_decodeResult_vtype};
  wire         queue_5_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_5 = {queue_dataIn_hi_lo_hi_hi_hi_5, queue_5_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_10 = {queue_dataIn_hi_lo_hi_hi_5, queue_dataIn_hi_lo_hi_lo_5};
  wire [11:0]  queue_dataIn_hi_lo_16 = {queue_dataIn_hi_lo_hi_10, queue_dataIn_hi_lo_lo_10};
  wire         queue_5_enq_bits_decodeResult_reverse;
  wire         queue_5_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_5 = {queue_5_enq_bits_decodeResult_reverse, queue_5_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_5_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_5 = {queue_dataIn_hi_hi_lo_lo_hi_5, queue_5_enq_bits_decodeResult_scheduler};
  wire         queue_5_enq_bits_decodeResult_popCount;
  wire         queue_5_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_popCount, queue_5_enq_bits_decodeResult_ffo};
  wire         queue_5_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_5 = {queue_dataIn_hi_hi_lo_hi_hi_5, queue_5_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_10 = {queue_dataIn_hi_hi_lo_hi_5, queue_dataIn_hi_hi_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_float;
  wire         queue_5_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_float, queue_5_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_5_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_5 = {queue_dataIn_hi_hi_hi_lo_hi_5, queue_5_enq_bits_decodeResult_topUop};
  wire         queue_5_enq_bits_decodeResult_orderReduce;
  wire         queue_5_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_orderReduce, queue_5_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_5_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_5 = {queue_dataIn_hi_hi_hi_hi_hi_5, queue_5_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_10 = {queue_dataIn_hi_hi_hi_hi_5, queue_dataIn_hi_hi_hi_lo_5};
  wire [16:0]  queue_dataIn_hi_hi_16 = {queue_dataIn_hi_hi_hi_10, queue_dataIn_hi_hi_lo_10};
  wire [28:0]  queue_dataIn_hi_16 = {queue_dataIn_hi_hi_16, queue_dataIn_hi_lo_16};
  wire [2:0]   queue_5_enq_bits_segment;
  wire [31:0]  queue_5_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_11 = {queue_5_enq_bits_segment, queue_5_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_11 = {queue_dataIn_lo_lo_hi_11, queue_dataIn_hi_15, queue_dataIn_lo_15};
  wire [1:0]   queue_5_enq_bits_loadStoreEEW;
  wire         queue_5_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_11 = {queue_5_enq_bits_loadStoreEEW, queue_5_enq_bits_mask};
  wire [4:0]   queue_5_enq_bits_vs2;
  wire [4:0]   queue_5_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_11 = {queue_5_enq_bits_vs2, queue_5_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_17 = {queue_dataIn_lo_hi_hi_11, queue_dataIn_lo_hi_lo_11};
  wire [80:0]  queue_dataIn_lo_17 = {queue_dataIn_lo_hi_17, queue_dataIn_lo_lo_11};
  wire         queue_5_enq_bits_lsWholeReg;
  wire [4:0]   queue_5_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_11 = {queue_5_enq_bits_lsWholeReg, queue_5_enq_bits_vs1};
  wire         queue_5_enq_bits_store;
  wire         queue_5_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_11 = {queue_5_enq_bits_store, queue_5_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_17 = {queue_dataIn_hi_lo_hi_11, queue_dataIn_hi_lo_lo_11};
  wire         queue_5_enq_bits_loadStore;
  wire         queue_5_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_11 = {queue_5_enq_bits_loadStore, queue_5_enq_bits_issueInst};
  wire [2:0]   queue_5_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_11 = {queue_5_enq_bits_instructionIndex, queue_dataIn_hi_16, queue_dataIn_lo_16};
  wire [60:0]  queue_dataIn_hi_hi_17 = {queue_dataIn_hi_hi_hi_11, queue_dataIn_hi_hi_lo_11};
  wire [68:0]  queue_dataIn_hi_17 = {queue_dataIn_hi_hi_17, queue_dataIn_hi_lo_17};
  wire [149:0] queue_dataIn_5 = {queue_dataIn_hi_17, queue_dataIn_lo_17};
  wire         queue_dataOut_5_csrInterface_vma = _queue_fifo_5_data_out[0];
  wire         queue_dataOut_5_csrInterface_vta = _queue_fifo_5_data_out[1];
  wire [1:0]   queue_dataOut_5_csrInterface_vxrm = _queue_fifo_5_data_out[3:2];
  wire [1:0]   queue_dataOut_5_csrInterface_vSew = _queue_fifo_5_data_out[5:4];
  wire [2:0]   queue_dataOut_5_csrInterface_vlmul = _queue_fifo_5_data_out[8:6];
  wire [11:0]  queue_dataOut_5_csrInterface_vStart = _queue_fifo_5_data_out[20:9];
  wire [11:0]  queue_dataOut_5_csrInterface_vl = _queue_fifo_5_data_out[32:21];
  wire [31:0]  queue_dataOut_5_readFromScalar = _queue_fifo_5_data_out[64:33];
  wire [2:0]   queue_dataOut_5_segment = _queue_fifo_5_data_out[67:65];
  wire         queue_dataOut_5_mask = _queue_fifo_5_data_out[68];
  wire [1:0]   queue_dataOut_5_loadStoreEEW = _queue_fifo_5_data_out[70:69];
  wire [4:0]   queue_dataOut_5_vd = _queue_fifo_5_data_out[75:71];
  wire [4:0]   queue_dataOut_5_vs2 = _queue_fifo_5_data_out[80:76];
  wire [4:0]   queue_dataOut_5_vs1 = _queue_fifo_5_data_out[85:81];
  wire         queue_dataOut_5_lsWholeReg = _queue_fifo_5_data_out[86];
  wire         queue_dataOut_5_special = _queue_fifo_5_data_out[87];
  wire         queue_dataOut_5_store = _queue_fifo_5_data_out[88];
  wire         queue_dataOut_5_issueInst = _queue_fifo_5_data_out[89];
  wire         queue_dataOut_5_loadStore = _queue_fifo_5_data_out[90];
  wire         queue_dataOut_5_decodeResult_logic = _queue_fifo_5_data_out[91];
  wire         queue_dataOut_5_decodeResult_adder = _queue_fifo_5_data_out[92];
  wire         queue_dataOut_5_decodeResult_shift = _queue_fifo_5_data_out[93];
  wire         queue_dataOut_5_decodeResult_multiplier = _queue_fifo_5_data_out[94];
  wire         queue_dataOut_5_decodeResult_divider = _queue_fifo_5_data_out[95];
  wire         queue_dataOut_5_decodeResult_multiCycle = _queue_fifo_5_data_out[96];
  wire         queue_dataOut_5_decodeResult_other = _queue_fifo_5_data_out[97];
  wire         queue_dataOut_5_decodeResult_unsigned0 = _queue_fifo_5_data_out[98];
  wire         queue_dataOut_5_decodeResult_unsigned1 = _queue_fifo_5_data_out[99];
  wire         queue_dataOut_5_decodeResult_itype = _queue_fifo_5_data_out[100];
  wire         queue_dataOut_5_decodeResult_nr = _queue_fifo_5_data_out[101];
  wire         queue_dataOut_5_decodeResult_red = _queue_fifo_5_data_out[102];
  wire         queue_dataOut_5_decodeResult_widenReduce = _queue_fifo_5_data_out[103];
  wire         queue_dataOut_5_decodeResult_targetRd = _queue_fifo_5_data_out[104];
  wire         queue_dataOut_5_decodeResult_slid = _queue_fifo_5_data_out[105];
  wire         queue_dataOut_5_decodeResult_gather = _queue_fifo_5_data_out[106];
  wire         queue_dataOut_5_decodeResult_gather16 = _queue_fifo_5_data_out[107];
  wire         queue_dataOut_5_decodeResult_compress = _queue_fifo_5_data_out[108];
  wire         queue_dataOut_5_decodeResult_unOrderWrite = _queue_fifo_5_data_out[109];
  wire         queue_dataOut_5_decodeResult_extend = _queue_fifo_5_data_out[110];
  wire         queue_dataOut_5_decodeResult_mv = _queue_fifo_5_data_out[111];
  wire         queue_dataOut_5_decodeResult_iota = _queue_fifo_5_data_out[112];
  wire [3:0]   queue_dataOut_5_decodeResult_uop = _queue_fifo_5_data_out[116:113];
  wire         queue_dataOut_5_decodeResult_maskLogic = _queue_fifo_5_data_out[117];
  wire         queue_dataOut_5_decodeResult_maskDestination = _queue_fifo_5_data_out[118];
  wire         queue_dataOut_5_decodeResult_maskSource = _queue_fifo_5_data_out[119];
  wire         queue_dataOut_5_decodeResult_readOnly = _queue_fifo_5_data_out[120];
  wire         queue_dataOut_5_decodeResult_vwmacc = _queue_fifo_5_data_out[121];
  wire         queue_dataOut_5_decodeResult_saturate = _queue_fifo_5_data_out[122];
  wire         queue_dataOut_5_decodeResult_special = _queue_fifo_5_data_out[123];
  wire         queue_dataOut_5_decodeResult_maskUnit = _queue_fifo_5_data_out[124];
  wire         queue_dataOut_5_decodeResult_crossWrite = _queue_fifo_5_data_out[125];
  wire         queue_dataOut_5_decodeResult_crossRead = _queue_fifo_5_data_out[126];
  wire         queue_dataOut_5_decodeResult_sWrite = _queue_fifo_5_data_out[127];
  wire         queue_dataOut_5_decodeResult_vtype = _queue_fifo_5_data_out[128];
  wire         queue_dataOut_5_decodeResult_sReadVD = _queue_fifo_5_data_out[129];
  wire         queue_dataOut_5_decodeResult_scheduler = _queue_fifo_5_data_out[130];
  wire         queue_dataOut_5_decodeResult_dontNeedExecuteInLane = _queue_fifo_5_data_out[131];
  wire         queue_dataOut_5_decodeResult_reverse = _queue_fifo_5_data_out[132];
  wire         queue_dataOut_5_decodeResult_average = _queue_fifo_5_data_out[133];
  wire         queue_dataOut_5_decodeResult_ffo = _queue_fifo_5_data_out[134];
  wire         queue_dataOut_5_decodeResult_popCount = _queue_fifo_5_data_out[135];
  wire [4:0]   queue_dataOut_5_decodeResult_topUop = _queue_fifo_5_data_out[140:136];
  wire         queue_dataOut_5_decodeResult_specialSlot = _queue_fifo_5_data_out[141];
  wire         queue_dataOut_5_decodeResult_float = _queue_fifo_5_data_out[142];
  wire [1:0]   queue_dataOut_5_decodeResult_fpExecutionType = _queue_fifo_5_data_out[144:143];
  wire         queue_dataOut_5_decodeResult_floatMul = _queue_fifo_5_data_out[145];
  wire         queue_dataOut_5_decodeResult_orderReduce = _queue_fifo_5_data_out[146];
  wire [2:0]   queue_dataOut_5_instructionIndex = _queue_fifo_5_data_out[149:147];
  wire         queue_5_enq_ready = ~_queue_fifo_5_full;
  wire         queue_5_enq_valid;
  assign queue_5_deq_valid = ~_queue_fifo_5_empty | queue_5_enq_valid;
  assign queue_5_deq_bits_instructionIndex = _queue_fifo_5_empty ? queue_5_enq_bits_instructionIndex : queue_dataOut_5_instructionIndex;
  assign queue_5_deq_bits_decodeResult_orderReduce = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_orderReduce : queue_dataOut_5_decodeResult_orderReduce;
  assign queue_5_deq_bits_decodeResult_floatMul = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_floatMul : queue_dataOut_5_decodeResult_floatMul;
  assign queue_5_deq_bits_decodeResult_fpExecutionType = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_fpExecutionType : queue_dataOut_5_decodeResult_fpExecutionType;
  assign queue_5_deq_bits_decodeResult_float = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_float : queue_dataOut_5_decodeResult_float;
  assign queue_5_deq_bits_decodeResult_specialSlot = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_specialSlot : queue_dataOut_5_decodeResult_specialSlot;
  assign queue_5_deq_bits_decodeResult_topUop = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_topUop : queue_dataOut_5_decodeResult_topUop;
  assign queue_5_deq_bits_decodeResult_popCount = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_popCount : queue_dataOut_5_decodeResult_popCount;
  assign queue_5_deq_bits_decodeResult_ffo = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_ffo : queue_dataOut_5_decodeResult_ffo;
  assign queue_5_deq_bits_decodeResult_average = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_average : queue_dataOut_5_decodeResult_average;
  assign queue_5_deq_bits_decodeResult_reverse = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_reverse : queue_dataOut_5_decodeResult_reverse;
  assign queue_5_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_5_decodeResult_dontNeedExecuteInLane;
  assign queue_5_deq_bits_decodeResult_scheduler = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_scheduler : queue_dataOut_5_decodeResult_scheduler;
  assign queue_5_deq_bits_decodeResult_sReadVD = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_sReadVD : queue_dataOut_5_decodeResult_sReadVD;
  assign queue_5_deq_bits_decodeResult_vtype = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_vtype : queue_dataOut_5_decodeResult_vtype;
  assign queue_5_deq_bits_decodeResult_sWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_sWrite : queue_dataOut_5_decodeResult_sWrite;
  assign queue_5_deq_bits_decodeResult_crossRead = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_crossRead : queue_dataOut_5_decodeResult_crossRead;
  assign queue_5_deq_bits_decodeResult_crossWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_crossWrite : queue_dataOut_5_decodeResult_crossWrite;
  assign queue_5_deq_bits_decodeResult_maskUnit = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskUnit : queue_dataOut_5_decodeResult_maskUnit;
  assign queue_5_deq_bits_decodeResult_special = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_special : queue_dataOut_5_decodeResult_special;
  assign queue_5_deq_bits_decodeResult_saturate = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_saturate : queue_dataOut_5_decodeResult_saturate;
  assign queue_5_deq_bits_decodeResult_vwmacc = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_vwmacc : queue_dataOut_5_decodeResult_vwmacc;
  assign queue_5_deq_bits_decodeResult_readOnly = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_readOnly : queue_dataOut_5_decodeResult_readOnly;
  assign queue_5_deq_bits_decodeResult_maskSource = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskSource : queue_dataOut_5_decodeResult_maskSource;
  assign queue_5_deq_bits_decodeResult_maskDestination = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskDestination : queue_dataOut_5_decodeResult_maskDestination;
  assign queue_5_deq_bits_decodeResult_maskLogic = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskLogic : queue_dataOut_5_decodeResult_maskLogic;
  assign queue_5_deq_bits_decodeResult_uop = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_uop : queue_dataOut_5_decodeResult_uop;
  assign queue_5_deq_bits_decodeResult_iota = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_iota : queue_dataOut_5_decodeResult_iota;
  assign queue_5_deq_bits_decodeResult_mv = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_mv : queue_dataOut_5_decodeResult_mv;
  assign queue_5_deq_bits_decodeResult_extend = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_extend : queue_dataOut_5_decodeResult_extend;
  assign queue_5_deq_bits_decodeResult_unOrderWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unOrderWrite : queue_dataOut_5_decodeResult_unOrderWrite;
  assign queue_5_deq_bits_decodeResult_compress = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_compress : queue_dataOut_5_decodeResult_compress;
  assign queue_5_deq_bits_decodeResult_gather16 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_gather16 : queue_dataOut_5_decodeResult_gather16;
  assign queue_5_deq_bits_decodeResult_gather = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_gather : queue_dataOut_5_decodeResult_gather;
  assign queue_5_deq_bits_decodeResult_slid = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_slid : queue_dataOut_5_decodeResult_slid;
  assign queue_5_deq_bits_decodeResult_targetRd = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_targetRd : queue_dataOut_5_decodeResult_targetRd;
  assign queue_5_deq_bits_decodeResult_widenReduce = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_widenReduce : queue_dataOut_5_decodeResult_widenReduce;
  assign queue_5_deq_bits_decodeResult_red = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_red : queue_dataOut_5_decodeResult_red;
  assign queue_5_deq_bits_decodeResult_nr = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_nr : queue_dataOut_5_decodeResult_nr;
  assign queue_5_deq_bits_decodeResult_itype = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_itype : queue_dataOut_5_decodeResult_itype;
  assign queue_5_deq_bits_decodeResult_unsigned1 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unsigned1 : queue_dataOut_5_decodeResult_unsigned1;
  assign queue_5_deq_bits_decodeResult_unsigned0 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unsigned0 : queue_dataOut_5_decodeResult_unsigned0;
  assign queue_5_deq_bits_decodeResult_other = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_other : queue_dataOut_5_decodeResult_other;
  assign queue_5_deq_bits_decodeResult_multiCycle = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_multiCycle : queue_dataOut_5_decodeResult_multiCycle;
  assign queue_5_deq_bits_decodeResult_divider = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_divider : queue_dataOut_5_decodeResult_divider;
  assign queue_5_deq_bits_decodeResult_multiplier = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_multiplier : queue_dataOut_5_decodeResult_multiplier;
  assign queue_5_deq_bits_decodeResult_shift = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_shift : queue_dataOut_5_decodeResult_shift;
  assign queue_5_deq_bits_decodeResult_adder = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_adder : queue_dataOut_5_decodeResult_adder;
  assign queue_5_deq_bits_decodeResult_logic = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_logic : queue_dataOut_5_decodeResult_logic;
  assign queue_5_deq_bits_loadStore = _queue_fifo_5_empty ? queue_5_enq_bits_loadStore : queue_dataOut_5_loadStore;
  assign queue_5_deq_bits_issueInst = _queue_fifo_5_empty ? queue_5_enq_bits_issueInst : queue_dataOut_5_issueInst;
  assign queue_5_deq_bits_store = _queue_fifo_5_empty ? queue_5_enq_bits_store : queue_dataOut_5_store;
  assign queue_5_deq_bits_special = _queue_fifo_5_empty ? queue_5_enq_bits_special : queue_dataOut_5_special;
  assign queue_5_deq_bits_lsWholeReg = _queue_fifo_5_empty ? queue_5_enq_bits_lsWholeReg : queue_dataOut_5_lsWholeReg;
  assign queue_5_deq_bits_vs1 = _queue_fifo_5_empty ? queue_5_enq_bits_vs1 : queue_dataOut_5_vs1;
  assign queue_5_deq_bits_vs2 = _queue_fifo_5_empty ? queue_5_enq_bits_vs2 : queue_dataOut_5_vs2;
  assign queue_5_deq_bits_vd = _queue_fifo_5_empty ? queue_5_enq_bits_vd : queue_dataOut_5_vd;
  assign queue_5_deq_bits_loadStoreEEW = _queue_fifo_5_empty ? queue_5_enq_bits_loadStoreEEW : queue_dataOut_5_loadStoreEEW;
  assign queue_5_deq_bits_mask = _queue_fifo_5_empty ? queue_5_enq_bits_mask : queue_dataOut_5_mask;
  assign queue_5_deq_bits_segment = _queue_fifo_5_empty ? queue_5_enq_bits_segment : queue_dataOut_5_segment;
  assign queue_5_deq_bits_readFromScalar = _queue_fifo_5_empty ? queue_5_enq_bits_readFromScalar : queue_dataOut_5_readFromScalar;
  assign queue_5_deq_bits_csrInterface_vl = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vl : queue_dataOut_5_csrInterface_vl;
  assign queue_5_deq_bits_csrInterface_vStart = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vStart : queue_dataOut_5_csrInterface_vStart;
  assign queue_5_deq_bits_csrInterface_vlmul = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vlmul : queue_dataOut_5_csrInterface_vlmul;
  assign queue_5_deq_bits_csrInterface_vSew = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vSew : queue_dataOut_5_csrInterface_vSew;
  assign queue_5_deq_bits_csrInterface_vxrm = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vxrm : queue_dataOut_5_csrInterface_vxrm;
  assign queue_5_deq_bits_csrInterface_vta = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vta : queue_dataOut_5_csrInterface_vta;
  assign queue_5_deq_bits_csrInterface_vma = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vma : queue_dataOut_5_csrInterface_vma;
  wire         laneVec_5_laneRequest_bits_issueInst = laneRequestSinkWire_5_ready & laneRequestSinkWire_5_valid;
  reg          releasePipe_pipe_v_5;
  wire         releasePipe_pipe_out_5_valid = releasePipe_pipe_v_5;
  wire         laneRequestSourceWire_5_ready;
  wire         validSource_5_valid = laneRequestSourceWire_5_ready & laneRequestSourceWire_5_valid;
  reg  [2:0]   tokenCheck_counter_5;
  wire [2:0]   tokenCheck_counterChange_5 = validSource_5_valid ? 3'h1 : 3'h7;
  assign tokenCheck_5 = ~(tokenCheck_counter_5[2]);
  assign laneRequestSourceWire_5_ready = tokenCheck_5;
  assign queue_5_enq_valid = validSink_5_valid;
  assign queue_5_enq_bits_instructionIndex = validSink_5_bits_instructionIndex;
  assign queue_5_enq_bits_decodeResult_orderReduce = validSink_5_bits_decodeResult_orderReduce;
  assign queue_5_enq_bits_decodeResult_floatMul = validSink_5_bits_decodeResult_floatMul;
  assign queue_5_enq_bits_decodeResult_fpExecutionType = validSink_5_bits_decodeResult_fpExecutionType;
  assign queue_5_enq_bits_decodeResult_float = validSink_5_bits_decodeResult_float;
  assign queue_5_enq_bits_decodeResult_specialSlot = validSink_5_bits_decodeResult_specialSlot;
  assign queue_5_enq_bits_decodeResult_topUop = validSink_5_bits_decodeResult_topUop;
  assign queue_5_enq_bits_decodeResult_popCount = validSink_5_bits_decodeResult_popCount;
  assign queue_5_enq_bits_decodeResult_ffo = validSink_5_bits_decodeResult_ffo;
  assign queue_5_enq_bits_decodeResult_average = validSink_5_bits_decodeResult_average;
  assign queue_5_enq_bits_decodeResult_reverse = validSink_5_bits_decodeResult_reverse;
  assign queue_5_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_5_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_5_enq_bits_decodeResult_scheduler = validSink_5_bits_decodeResult_scheduler;
  assign queue_5_enq_bits_decodeResult_sReadVD = validSink_5_bits_decodeResult_sReadVD;
  assign queue_5_enq_bits_decodeResult_vtype = validSink_5_bits_decodeResult_vtype;
  assign queue_5_enq_bits_decodeResult_sWrite = validSink_5_bits_decodeResult_sWrite;
  assign queue_5_enq_bits_decodeResult_crossRead = validSink_5_bits_decodeResult_crossRead;
  assign queue_5_enq_bits_decodeResult_crossWrite = validSink_5_bits_decodeResult_crossWrite;
  assign queue_5_enq_bits_decodeResult_maskUnit = validSink_5_bits_decodeResult_maskUnit;
  assign queue_5_enq_bits_decodeResult_special = validSink_5_bits_decodeResult_special;
  assign queue_5_enq_bits_decodeResult_saturate = validSink_5_bits_decodeResult_saturate;
  assign queue_5_enq_bits_decodeResult_vwmacc = validSink_5_bits_decodeResult_vwmacc;
  assign queue_5_enq_bits_decodeResult_readOnly = validSink_5_bits_decodeResult_readOnly;
  assign queue_5_enq_bits_decodeResult_maskSource = validSink_5_bits_decodeResult_maskSource;
  assign queue_5_enq_bits_decodeResult_maskDestination = validSink_5_bits_decodeResult_maskDestination;
  assign queue_5_enq_bits_decodeResult_maskLogic = validSink_5_bits_decodeResult_maskLogic;
  assign queue_5_enq_bits_decodeResult_uop = validSink_5_bits_decodeResult_uop;
  assign queue_5_enq_bits_decodeResult_iota = validSink_5_bits_decodeResult_iota;
  assign queue_5_enq_bits_decodeResult_mv = validSink_5_bits_decodeResult_mv;
  assign queue_5_enq_bits_decodeResult_extend = validSink_5_bits_decodeResult_extend;
  assign queue_5_enq_bits_decodeResult_unOrderWrite = validSink_5_bits_decodeResult_unOrderWrite;
  assign queue_5_enq_bits_decodeResult_compress = validSink_5_bits_decodeResult_compress;
  assign queue_5_enq_bits_decodeResult_gather16 = validSink_5_bits_decodeResult_gather16;
  assign queue_5_enq_bits_decodeResult_gather = validSink_5_bits_decodeResult_gather;
  assign queue_5_enq_bits_decodeResult_slid = validSink_5_bits_decodeResult_slid;
  assign queue_5_enq_bits_decodeResult_targetRd = validSink_5_bits_decodeResult_targetRd;
  assign queue_5_enq_bits_decodeResult_widenReduce = validSink_5_bits_decodeResult_widenReduce;
  assign queue_5_enq_bits_decodeResult_red = validSink_5_bits_decodeResult_red;
  assign queue_5_enq_bits_decodeResult_nr = validSink_5_bits_decodeResult_nr;
  assign queue_5_enq_bits_decodeResult_itype = validSink_5_bits_decodeResult_itype;
  assign queue_5_enq_bits_decodeResult_unsigned1 = validSink_5_bits_decodeResult_unsigned1;
  assign queue_5_enq_bits_decodeResult_unsigned0 = validSink_5_bits_decodeResult_unsigned0;
  assign queue_5_enq_bits_decodeResult_other = validSink_5_bits_decodeResult_other;
  assign queue_5_enq_bits_decodeResult_multiCycle = validSink_5_bits_decodeResult_multiCycle;
  assign queue_5_enq_bits_decodeResult_divider = validSink_5_bits_decodeResult_divider;
  assign queue_5_enq_bits_decodeResult_multiplier = validSink_5_bits_decodeResult_multiplier;
  assign queue_5_enq_bits_decodeResult_shift = validSink_5_bits_decodeResult_shift;
  assign queue_5_enq_bits_decodeResult_adder = validSink_5_bits_decodeResult_adder;
  assign queue_5_enq_bits_decodeResult_logic = validSink_5_bits_decodeResult_logic;
  assign queue_5_enq_bits_loadStore = validSink_5_bits_loadStore;
  assign queue_5_enq_bits_issueInst = validSink_5_bits_issueInst;
  assign queue_5_enq_bits_store = validSink_5_bits_store;
  assign queue_5_enq_bits_special = validSink_5_bits_special;
  assign queue_5_enq_bits_lsWholeReg = validSink_5_bits_lsWholeReg;
  assign queue_5_enq_bits_vs1 = validSink_5_bits_vs1;
  assign queue_5_enq_bits_vs2 = validSink_5_bits_vs2;
  assign queue_5_enq_bits_vd = validSink_5_bits_vd;
  assign queue_5_enq_bits_loadStoreEEW = validSink_5_bits_loadStoreEEW;
  assign queue_5_enq_bits_mask = validSink_5_bits_mask;
  assign queue_5_enq_bits_segment = validSink_5_bits_segment;
  assign queue_5_enq_bits_readFromScalar = validSink_5_bits_readFromScalar;
  assign queue_5_enq_bits_csrInterface_vl = validSink_5_bits_csrInterface_vl;
  assign queue_5_enq_bits_csrInterface_vStart = validSink_5_bits_csrInterface_vStart;
  assign queue_5_enq_bits_csrInterface_vlmul = validSink_5_bits_csrInterface_vlmul;
  assign queue_5_enq_bits_csrInterface_vSew = validSink_5_bits_csrInterface_vSew;
  assign queue_5_enq_bits_csrInterface_vxrm = validSink_5_bits_csrInterface_vxrm;
  assign queue_5_enq_bits_csrInterface_vta = validSink_5_bits_csrInterface_vta;
  assign queue_5_enq_bits_csrInterface_vma = validSink_5_bits_csrInterface_vma;
  reg          shifterReg_5_0_valid;
  assign validSink_5_valid = shifterReg_5_0_valid;
  reg  [2:0]   shifterReg_5_0_bits_instructionIndex;
  assign validSink_5_bits_instructionIndex = shifterReg_5_0_bits_instructionIndex;
  reg          shifterReg_5_0_bits_decodeResult_orderReduce;
  assign validSink_5_bits_decodeResult_orderReduce = shifterReg_5_0_bits_decodeResult_orderReduce;
  reg          shifterReg_5_0_bits_decodeResult_floatMul;
  assign validSink_5_bits_decodeResult_floatMul = shifterReg_5_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_5_0_bits_decodeResult_fpExecutionType;
  assign validSink_5_bits_decodeResult_fpExecutionType = shifterReg_5_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_5_0_bits_decodeResult_float;
  assign validSink_5_bits_decodeResult_float = shifterReg_5_0_bits_decodeResult_float;
  reg          shifterReg_5_0_bits_decodeResult_specialSlot;
  assign validSink_5_bits_decodeResult_specialSlot = shifterReg_5_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_5_0_bits_decodeResult_topUop;
  assign validSink_5_bits_decodeResult_topUop = shifterReg_5_0_bits_decodeResult_topUop;
  reg          shifterReg_5_0_bits_decodeResult_popCount;
  assign validSink_5_bits_decodeResult_popCount = shifterReg_5_0_bits_decodeResult_popCount;
  reg          shifterReg_5_0_bits_decodeResult_ffo;
  assign validSink_5_bits_decodeResult_ffo = shifterReg_5_0_bits_decodeResult_ffo;
  reg          shifterReg_5_0_bits_decodeResult_average;
  assign validSink_5_bits_decodeResult_average = shifterReg_5_0_bits_decodeResult_average;
  reg          shifterReg_5_0_bits_decodeResult_reverse;
  assign validSink_5_bits_decodeResult_reverse = shifterReg_5_0_bits_decodeResult_reverse;
  reg          shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_5_bits_decodeResult_dontNeedExecuteInLane = shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_5_0_bits_decodeResult_scheduler;
  assign validSink_5_bits_decodeResult_scheduler = shifterReg_5_0_bits_decodeResult_scheduler;
  reg          shifterReg_5_0_bits_decodeResult_sReadVD;
  assign validSink_5_bits_decodeResult_sReadVD = shifterReg_5_0_bits_decodeResult_sReadVD;
  reg          shifterReg_5_0_bits_decodeResult_vtype;
  assign validSink_5_bits_decodeResult_vtype = shifterReg_5_0_bits_decodeResult_vtype;
  reg          shifterReg_5_0_bits_decodeResult_sWrite;
  assign validSink_5_bits_decodeResult_sWrite = shifterReg_5_0_bits_decodeResult_sWrite;
  reg          shifterReg_5_0_bits_decodeResult_crossRead;
  assign validSink_5_bits_decodeResult_crossRead = shifterReg_5_0_bits_decodeResult_crossRead;
  reg          shifterReg_5_0_bits_decodeResult_crossWrite;
  assign validSink_5_bits_decodeResult_crossWrite = shifterReg_5_0_bits_decodeResult_crossWrite;
  reg          shifterReg_5_0_bits_decodeResult_maskUnit;
  assign validSink_5_bits_decodeResult_maskUnit = shifterReg_5_0_bits_decodeResult_maskUnit;
  reg          shifterReg_5_0_bits_decodeResult_special;
  assign validSink_5_bits_decodeResult_special = shifterReg_5_0_bits_decodeResult_special;
  reg          shifterReg_5_0_bits_decodeResult_saturate;
  assign validSink_5_bits_decodeResult_saturate = shifterReg_5_0_bits_decodeResult_saturate;
  reg          shifterReg_5_0_bits_decodeResult_vwmacc;
  assign validSink_5_bits_decodeResult_vwmacc = shifterReg_5_0_bits_decodeResult_vwmacc;
  reg          shifterReg_5_0_bits_decodeResult_readOnly;
  assign validSink_5_bits_decodeResult_readOnly = shifterReg_5_0_bits_decodeResult_readOnly;
  reg          shifterReg_5_0_bits_decodeResult_maskSource;
  assign validSink_5_bits_decodeResult_maskSource = shifterReg_5_0_bits_decodeResult_maskSource;
  reg          shifterReg_5_0_bits_decodeResult_maskDestination;
  assign validSink_5_bits_decodeResult_maskDestination = shifterReg_5_0_bits_decodeResult_maskDestination;
  reg          shifterReg_5_0_bits_decodeResult_maskLogic;
  assign validSink_5_bits_decodeResult_maskLogic = shifterReg_5_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_5_0_bits_decodeResult_uop;
  assign validSink_5_bits_decodeResult_uop = shifterReg_5_0_bits_decodeResult_uop;
  reg          shifterReg_5_0_bits_decodeResult_iota;
  assign validSink_5_bits_decodeResult_iota = shifterReg_5_0_bits_decodeResult_iota;
  reg          shifterReg_5_0_bits_decodeResult_mv;
  assign validSink_5_bits_decodeResult_mv = shifterReg_5_0_bits_decodeResult_mv;
  reg          shifterReg_5_0_bits_decodeResult_extend;
  assign validSink_5_bits_decodeResult_extend = shifterReg_5_0_bits_decodeResult_extend;
  reg          shifterReg_5_0_bits_decodeResult_unOrderWrite;
  assign validSink_5_bits_decodeResult_unOrderWrite = shifterReg_5_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_5_0_bits_decodeResult_compress;
  assign validSink_5_bits_decodeResult_compress = shifterReg_5_0_bits_decodeResult_compress;
  reg          shifterReg_5_0_bits_decodeResult_gather16;
  assign validSink_5_bits_decodeResult_gather16 = shifterReg_5_0_bits_decodeResult_gather16;
  reg          shifterReg_5_0_bits_decodeResult_gather;
  assign validSink_5_bits_decodeResult_gather = shifterReg_5_0_bits_decodeResult_gather;
  reg          shifterReg_5_0_bits_decodeResult_slid;
  assign validSink_5_bits_decodeResult_slid = shifterReg_5_0_bits_decodeResult_slid;
  reg          shifterReg_5_0_bits_decodeResult_targetRd;
  assign validSink_5_bits_decodeResult_targetRd = shifterReg_5_0_bits_decodeResult_targetRd;
  reg          shifterReg_5_0_bits_decodeResult_widenReduce;
  assign validSink_5_bits_decodeResult_widenReduce = shifterReg_5_0_bits_decodeResult_widenReduce;
  reg          shifterReg_5_0_bits_decodeResult_red;
  assign validSink_5_bits_decodeResult_red = shifterReg_5_0_bits_decodeResult_red;
  reg          shifterReg_5_0_bits_decodeResult_nr;
  assign validSink_5_bits_decodeResult_nr = shifterReg_5_0_bits_decodeResult_nr;
  reg          shifterReg_5_0_bits_decodeResult_itype;
  assign validSink_5_bits_decodeResult_itype = shifterReg_5_0_bits_decodeResult_itype;
  reg          shifterReg_5_0_bits_decodeResult_unsigned1;
  assign validSink_5_bits_decodeResult_unsigned1 = shifterReg_5_0_bits_decodeResult_unsigned1;
  reg          shifterReg_5_0_bits_decodeResult_unsigned0;
  assign validSink_5_bits_decodeResult_unsigned0 = shifterReg_5_0_bits_decodeResult_unsigned0;
  reg          shifterReg_5_0_bits_decodeResult_other;
  assign validSink_5_bits_decodeResult_other = shifterReg_5_0_bits_decodeResult_other;
  reg          shifterReg_5_0_bits_decodeResult_multiCycle;
  assign validSink_5_bits_decodeResult_multiCycle = shifterReg_5_0_bits_decodeResult_multiCycle;
  reg          shifterReg_5_0_bits_decodeResult_divider;
  assign validSink_5_bits_decodeResult_divider = shifterReg_5_0_bits_decodeResult_divider;
  reg          shifterReg_5_0_bits_decodeResult_multiplier;
  assign validSink_5_bits_decodeResult_multiplier = shifterReg_5_0_bits_decodeResult_multiplier;
  reg          shifterReg_5_0_bits_decodeResult_shift;
  assign validSink_5_bits_decodeResult_shift = shifterReg_5_0_bits_decodeResult_shift;
  reg          shifterReg_5_0_bits_decodeResult_adder;
  assign validSink_5_bits_decodeResult_adder = shifterReg_5_0_bits_decodeResult_adder;
  reg          shifterReg_5_0_bits_decodeResult_logic;
  assign validSink_5_bits_decodeResult_logic = shifterReg_5_0_bits_decodeResult_logic;
  reg          shifterReg_5_0_bits_loadStore;
  assign validSink_5_bits_loadStore = shifterReg_5_0_bits_loadStore;
  reg          shifterReg_5_0_bits_issueInst;
  assign validSink_5_bits_issueInst = shifterReg_5_0_bits_issueInst;
  reg          shifterReg_5_0_bits_store;
  assign validSink_5_bits_store = shifterReg_5_0_bits_store;
  reg          shifterReg_5_0_bits_special;
  assign validSink_5_bits_special = shifterReg_5_0_bits_special;
  reg          shifterReg_5_0_bits_lsWholeReg;
  assign validSink_5_bits_lsWholeReg = shifterReg_5_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_5_0_bits_vs1;
  assign validSink_5_bits_vs1 = shifterReg_5_0_bits_vs1;
  reg  [4:0]   shifterReg_5_0_bits_vs2;
  assign validSink_5_bits_vs2 = shifterReg_5_0_bits_vs2;
  reg  [4:0]   shifterReg_5_0_bits_vd;
  assign validSink_5_bits_vd = shifterReg_5_0_bits_vd;
  reg  [1:0]   shifterReg_5_0_bits_loadStoreEEW;
  assign validSink_5_bits_loadStoreEEW = shifterReg_5_0_bits_loadStoreEEW;
  reg          shifterReg_5_0_bits_mask;
  assign validSink_5_bits_mask = shifterReg_5_0_bits_mask;
  reg  [2:0]   shifterReg_5_0_bits_segment;
  assign validSink_5_bits_segment = shifterReg_5_0_bits_segment;
  reg  [31:0]  shifterReg_5_0_bits_readFromScalar;
  assign validSink_5_bits_readFromScalar = shifterReg_5_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_5_0_bits_csrInterface_vl;
  assign validSink_5_bits_csrInterface_vl = shifterReg_5_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_5_0_bits_csrInterface_vStart;
  assign validSink_5_bits_csrInterface_vStart = shifterReg_5_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_5_0_bits_csrInterface_vlmul;
  assign validSink_5_bits_csrInterface_vlmul = shifterReg_5_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_5_0_bits_csrInterface_vSew;
  assign validSink_5_bits_csrInterface_vSew = shifterReg_5_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_5_0_bits_csrInterface_vxrm;
  assign validSink_5_bits_csrInterface_vxrm = shifterReg_5_0_bits_csrInterface_vxrm;
  reg          shifterReg_5_0_bits_csrInterface_vta;
  assign validSink_5_bits_csrInterface_vta = shifterReg_5_0_bits_csrInterface_vta;
  reg          shifterReg_5_0_bits_csrInterface_vma;
  assign validSink_5_bits_csrInterface_vma = shifterReg_5_0_bits_csrInterface_vma;
  wire         shifterValid_5 = shifterReg_5_0_valid | validSource_5_valid;
  wire         validSink_6_valid;
  wire [2:0]   validSink_6_bits_instructionIndex;
  wire         validSink_6_bits_decodeResult_orderReduce;
  wire         validSink_6_bits_decodeResult_floatMul;
  wire [1:0]   validSink_6_bits_decodeResult_fpExecutionType;
  wire         validSink_6_bits_decodeResult_float;
  wire         validSink_6_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_6_bits_decodeResult_topUop;
  wire         validSink_6_bits_decodeResult_popCount;
  wire         validSink_6_bits_decodeResult_ffo;
  wire         validSink_6_bits_decodeResult_average;
  wire         validSink_6_bits_decodeResult_reverse;
  wire         validSink_6_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_6_bits_decodeResult_scheduler;
  wire         validSink_6_bits_decodeResult_sReadVD;
  wire         validSink_6_bits_decodeResult_vtype;
  wire         validSink_6_bits_decodeResult_sWrite;
  wire         validSink_6_bits_decodeResult_crossRead;
  wire         validSink_6_bits_decodeResult_crossWrite;
  wire         validSink_6_bits_decodeResult_maskUnit;
  wire         validSink_6_bits_decodeResult_special;
  wire         validSink_6_bits_decodeResult_saturate;
  wire         validSink_6_bits_decodeResult_vwmacc;
  wire         validSink_6_bits_decodeResult_readOnly;
  wire         validSink_6_bits_decodeResult_maskSource;
  wire         validSink_6_bits_decodeResult_maskDestination;
  wire         validSink_6_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_6_bits_decodeResult_uop;
  wire         validSink_6_bits_decodeResult_iota;
  wire         validSink_6_bits_decodeResult_mv;
  wire         validSink_6_bits_decodeResult_extend;
  wire         validSink_6_bits_decodeResult_unOrderWrite;
  wire         validSink_6_bits_decodeResult_compress;
  wire         validSink_6_bits_decodeResult_gather16;
  wire         validSink_6_bits_decodeResult_gather;
  wire         validSink_6_bits_decodeResult_slid;
  wire         validSink_6_bits_decodeResult_targetRd;
  wire         validSink_6_bits_decodeResult_widenReduce;
  wire         validSink_6_bits_decodeResult_red;
  wire         validSink_6_bits_decodeResult_nr;
  wire         validSink_6_bits_decodeResult_itype;
  wire         validSink_6_bits_decodeResult_unsigned1;
  wire         validSink_6_bits_decodeResult_unsigned0;
  wire         validSink_6_bits_decodeResult_other;
  wire         validSink_6_bits_decodeResult_multiCycle;
  wire         validSink_6_bits_decodeResult_divider;
  wire         validSink_6_bits_decodeResult_multiplier;
  wire         validSink_6_bits_decodeResult_shift;
  wire         validSink_6_bits_decodeResult_adder;
  wire         validSink_6_bits_decodeResult_logic;
  wire         validSink_6_bits_loadStore;
  wire         validSink_6_bits_issueInst;
  wire         validSink_6_bits_store;
  wire         validSink_6_bits_special;
  wire         validSink_6_bits_lsWholeReg;
  wire [4:0]   validSink_6_bits_vs1;
  wire [4:0]   validSink_6_bits_vs2;
  wire [4:0]   validSink_6_bits_vd;
  wire [1:0]   validSink_6_bits_loadStoreEEW;
  wire         validSink_6_bits_mask;
  wire [2:0]   validSink_6_bits_segment;
  wire [31:0]  validSink_6_bits_readFromScalar;
  wire [11:0]  validSink_6_bits_csrInterface_vl;
  wire [11:0]  validSink_6_bits_csrInterface_vStart;
  wire [2:0]   validSink_6_bits_csrInterface_vlmul;
  wire [1:0]   validSink_6_bits_csrInterface_vSew;
  wire [1:0]   validSink_6_bits_csrInterface_vxrm;
  wire         validSink_6_bits_csrInterface_vta;
  wire         validSink_6_bits_csrInterface_vma;
  wire         laneRequestSinkWire_6_valid = queue_6_deq_valid;
  wire [2:0]   laneRequestSinkWire_6_bits_instructionIndex = queue_6_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_6_bits_decodeResult_orderReduce = queue_6_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_6_bits_decodeResult_floatMul = queue_6_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_6_bits_decodeResult_fpExecutionType = queue_6_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_6_bits_decodeResult_float = queue_6_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_6_bits_decodeResult_specialSlot = queue_6_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_6_bits_decodeResult_topUop = queue_6_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_6_bits_decodeResult_popCount = queue_6_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_6_bits_decodeResult_ffo = queue_6_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_6_bits_decodeResult_average = queue_6_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_6_bits_decodeResult_reverse = queue_6_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_6_bits_decodeResult_dontNeedExecuteInLane = queue_6_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_6_bits_decodeResult_scheduler = queue_6_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_6_bits_decodeResult_sReadVD = queue_6_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_6_bits_decodeResult_vtype = queue_6_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_6_bits_decodeResult_sWrite = queue_6_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_crossRead = queue_6_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_6_bits_decodeResult_crossWrite = queue_6_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskUnit = queue_6_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_6_bits_decodeResult_special = queue_6_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_6_bits_decodeResult_saturate = queue_6_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_6_bits_decodeResult_vwmacc = queue_6_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_6_bits_decodeResult_readOnly = queue_6_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskSource = queue_6_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskDestination = queue_6_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskLogic = queue_6_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_6_bits_decodeResult_uop = queue_6_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_6_bits_decodeResult_iota = queue_6_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_6_bits_decodeResult_mv = queue_6_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_6_bits_decodeResult_extend = queue_6_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_6_bits_decodeResult_unOrderWrite = queue_6_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_compress = queue_6_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_6_bits_decodeResult_gather16 = queue_6_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_6_bits_decodeResult_gather = queue_6_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_6_bits_decodeResult_slid = queue_6_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_6_bits_decodeResult_targetRd = queue_6_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_6_bits_decodeResult_widenReduce = queue_6_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_6_bits_decodeResult_red = queue_6_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_6_bits_decodeResult_nr = queue_6_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_6_bits_decodeResult_itype = queue_6_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_6_bits_decodeResult_unsigned1 = queue_6_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_6_bits_decodeResult_unsigned0 = queue_6_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_6_bits_decodeResult_other = queue_6_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_6_bits_decodeResult_multiCycle = queue_6_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_6_bits_decodeResult_divider = queue_6_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_6_bits_decodeResult_multiplier = queue_6_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_6_bits_decodeResult_shift = queue_6_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_6_bits_decodeResult_adder = queue_6_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_6_bits_decodeResult_logic = queue_6_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_6_bits_loadStore = queue_6_deq_bits_loadStore;
  wire         laneRequestSinkWire_6_bits_issueInst = queue_6_deq_bits_issueInst;
  wire         laneRequestSinkWire_6_bits_store = queue_6_deq_bits_store;
  wire         laneRequestSinkWire_6_bits_special = queue_6_deq_bits_special;
  wire         laneRequestSinkWire_6_bits_lsWholeReg = queue_6_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_6_bits_vs1 = queue_6_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_6_bits_vs2 = queue_6_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_6_bits_vd = queue_6_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_6_bits_loadStoreEEW = queue_6_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_6_bits_mask = queue_6_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_6_bits_segment = queue_6_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_6_bits_readFromScalar = queue_6_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_6_bits_csrInterface_vl = queue_6_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_6_bits_csrInterface_vStart = queue_6_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_6_bits_csrInterface_vlmul = queue_6_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_6_bits_csrInterface_vSew = queue_6_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_6_bits_csrInterface_vxrm = queue_6_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_6_bits_csrInterface_vta = queue_6_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_6_bits_csrInterface_vma = queue_6_deq_bits_csrInterface_vma;
  wire [1:0]   queue_6_enq_bits_csrInterface_vxrm;
  wire         queue_6_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_18 = {queue_6_enq_bits_csrInterface_vxrm, queue_6_enq_bits_csrInterface_vta};
  wire         queue_6_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_18 = {queue_dataIn_lo_hi_18, queue_6_enq_bits_csrInterface_vma};
  wire [2:0]   queue_6_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_6_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_18 = {queue_6_enq_bits_csrInterface_vlmul, queue_6_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_6_enq_bits_csrInterface_vl;
  wire [11:0]  queue_6_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_18 = {queue_6_enq_bits_csrInterface_vl, queue_6_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_18 = {queue_dataIn_hi_hi_18, queue_dataIn_hi_lo_18};
  wire         queue_6_enq_bits_decodeResult_shift;
  wire         queue_6_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_6 = {queue_6_enq_bits_decodeResult_shift, queue_6_enq_bits_decodeResult_adder};
  wire         queue_6_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_6 = {queue_dataIn_lo_lo_lo_lo_hi_6, queue_6_enq_bits_decodeResult_logic};
  wire         queue_6_enq_bits_decodeResult_multiCycle;
  wire         queue_6_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_multiCycle, queue_6_enq_bits_decodeResult_divider};
  wire         queue_6_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_6 = {queue_dataIn_lo_lo_lo_hi_hi_6, queue_6_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_6 = {queue_dataIn_lo_lo_lo_hi_6, queue_dataIn_lo_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_unsigned1;
  wire         queue_6_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_unsigned1, queue_6_enq_bits_decodeResult_unsigned0};
  wire         queue_6_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_6 = {queue_dataIn_lo_lo_hi_lo_hi_6, queue_6_enq_bits_decodeResult_other};
  wire         queue_6_enq_bits_decodeResult_red;
  wire         queue_6_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_red, queue_6_enq_bits_decodeResult_nr};
  wire         queue_6_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_6 = {queue_dataIn_lo_lo_hi_hi_hi_6, queue_6_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_12 = {queue_dataIn_lo_lo_hi_hi_6, queue_dataIn_lo_lo_hi_lo_6};
  wire [11:0]  queue_dataIn_lo_lo_12 = {queue_dataIn_lo_lo_hi_12, queue_dataIn_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_slid;
  wire         queue_6_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_6 = {queue_6_enq_bits_decodeResult_slid, queue_6_enq_bits_decodeResult_targetRd};
  wire         queue_6_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_6 = {queue_dataIn_lo_hi_lo_lo_hi_6, queue_6_enq_bits_decodeResult_widenReduce};
  wire         queue_6_enq_bits_decodeResult_compress;
  wire         queue_6_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_compress, queue_6_enq_bits_decodeResult_gather16};
  wire         queue_6_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_6 = {queue_dataIn_lo_hi_lo_hi_hi_6, queue_6_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_12 = {queue_dataIn_lo_hi_lo_hi_6, queue_dataIn_lo_hi_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_mv;
  wire         queue_6_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_mv, queue_6_enq_bits_decodeResult_extend};
  wire         queue_6_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_6 = {queue_dataIn_lo_hi_hi_lo_hi_6, queue_6_enq_bits_decodeResult_unOrderWrite};
  wire         queue_6_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_6_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_maskLogic, queue_6_enq_bits_decodeResult_uop};
  wire         queue_6_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_6 = {queue_dataIn_lo_hi_hi_hi_hi_6, queue_6_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_12 = {queue_dataIn_lo_hi_hi_hi_6, queue_dataIn_lo_hi_hi_lo_6};
  wire [14:0]  queue_dataIn_lo_hi_19 = {queue_dataIn_lo_hi_hi_12, queue_dataIn_lo_hi_lo_12};
  wire [26:0]  queue_dataIn_lo_19 = {queue_dataIn_lo_hi_19, queue_dataIn_lo_lo_12};
  wire         queue_6_enq_bits_decodeResult_readOnly;
  wire         queue_6_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_6 = {queue_6_enq_bits_decodeResult_readOnly, queue_6_enq_bits_decodeResult_maskSource};
  wire         queue_6_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_6 = {queue_dataIn_hi_lo_lo_lo_hi_6, queue_6_enq_bits_decodeResult_maskDestination};
  wire         queue_6_enq_bits_decodeResult_special;
  wire         queue_6_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_special, queue_6_enq_bits_decodeResult_saturate};
  wire         queue_6_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_6 = {queue_dataIn_hi_lo_lo_hi_hi_6, queue_6_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_12 = {queue_dataIn_hi_lo_lo_hi_6, queue_dataIn_hi_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_crossRead;
  wire         queue_6_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_crossRead, queue_6_enq_bits_decodeResult_crossWrite};
  wire         queue_6_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_6 = {queue_dataIn_hi_lo_hi_lo_hi_6, queue_6_enq_bits_decodeResult_maskUnit};
  wire         queue_6_enq_bits_decodeResult_sReadVD;
  wire         queue_6_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_sReadVD, queue_6_enq_bits_decodeResult_vtype};
  wire         queue_6_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_6 = {queue_dataIn_hi_lo_hi_hi_hi_6, queue_6_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_12 = {queue_dataIn_hi_lo_hi_hi_6, queue_dataIn_hi_lo_hi_lo_6};
  wire [11:0]  queue_dataIn_hi_lo_19 = {queue_dataIn_hi_lo_hi_12, queue_dataIn_hi_lo_lo_12};
  wire         queue_6_enq_bits_decodeResult_reverse;
  wire         queue_6_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_6 = {queue_6_enq_bits_decodeResult_reverse, queue_6_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_6_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_6 = {queue_dataIn_hi_hi_lo_lo_hi_6, queue_6_enq_bits_decodeResult_scheduler};
  wire         queue_6_enq_bits_decodeResult_popCount;
  wire         queue_6_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_popCount, queue_6_enq_bits_decodeResult_ffo};
  wire         queue_6_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_6 = {queue_dataIn_hi_hi_lo_hi_hi_6, queue_6_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_12 = {queue_dataIn_hi_hi_lo_hi_6, queue_dataIn_hi_hi_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_float;
  wire         queue_6_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_float, queue_6_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_6_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_6 = {queue_dataIn_hi_hi_hi_lo_hi_6, queue_6_enq_bits_decodeResult_topUop};
  wire         queue_6_enq_bits_decodeResult_orderReduce;
  wire         queue_6_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_orderReduce, queue_6_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_6_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_6 = {queue_dataIn_hi_hi_hi_hi_hi_6, queue_6_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_12 = {queue_dataIn_hi_hi_hi_hi_6, queue_dataIn_hi_hi_hi_lo_6};
  wire [16:0]  queue_dataIn_hi_hi_19 = {queue_dataIn_hi_hi_hi_12, queue_dataIn_hi_hi_lo_12};
  wire [28:0]  queue_dataIn_hi_19 = {queue_dataIn_hi_hi_19, queue_dataIn_hi_lo_19};
  wire [2:0]   queue_6_enq_bits_segment;
  wire [31:0]  queue_6_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_13 = {queue_6_enq_bits_segment, queue_6_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_13 = {queue_dataIn_lo_lo_hi_13, queue_dataIn_hi_18, queue_dataIn_lo_18};
  wire [1:0]   queue_6_enq_bits_loadStoreEEW;
  wire         queue_6_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_13 = {queue_6_enq_bits_loadStoreEEW, queue_6_enq_bits_mask};
  wire [4:0]   queue_6_enq_bits_vs2;
  wire [4:0]   queue_6_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_13 = {queue_6_enq_bits_vs2, queue_6_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_20 = {queue_dataIn_lo_hi_hi_13, queue_dataIn_lo_hi_lo_13};
  wire [80:0]  queue_dataIn_lo_20 = {queue_dataIn_lo_hi_20, queue_dataIn_lo_lo_13};
  wire         queue_6_enq_bits_lsWholeReg;
  wire [4:0]   queue_6_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_13 = {queue_6_enq_bits_lsWholeReg, queue_6_enq_bits_vs1};
  wire         queue_6_enq_bits_store;
  wire         queue_6_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_13 = {queue_6_enq_bits_store, queue_6_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_20 = {queue_dataIn_hi_lo_hi_13, queue_dataIn_hi_lo_lo_13};
  wire         queue_6_enq_bits_loadStore;
  wire         queue_6_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_13 = {queue_6_enq_bits_loadStore, queue_6_enq_bits_issueInst};
  wire [2:0]   queue_6_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_13 = {queue_6_enq_bits_instructionIndex, queue_dataIn_hi_19, queue_dataIn_lo_19};
  wire [60:0]  queue_dataIn_hi_hi_20 = {queue_dataIn_hi_hi_hi_13, queue_dataIn_hi_hi_lo_13};
  wire [68:0]  queue_dataIn_hi_20 = {queue_dataIn_hi_hi_20, queue_dataIn_hi_lo_20};
  wire [149:0] queue_dataIn_6 = {queue_dataIn_hi_20, queue_dataIn_lo_20};
  wire         queue_dataOut_6_csrInterface_vma = _queue_fifo_6_data_out[0];
  wire         queue_dataOut_6_csrInterface_vta = _queue_fifo_6_data_out[1];
  wire [1:0]   queue_dataOut_6_csrInterface_vxrm = _queue_fifo_6_data_out[3:2];
  wire [1:0]   queue_dataOut_6_csrInterface_vSew = _queue_fifo_6_data_out[5:4];
  wire [2:0]   queue_dataOut_6_csrInterface_vlmul = _queue_fifo_6_data_out[8:6];
  wire [11:0]  queue_dataOut_6_csrInterface_vStart = _queue_fifo_6_data_out[20:9];
  wire [11:0]  queue_dataOut_6_csrInterface_vl = _queue_fifo_6_data_out[32:21];
  wire [31:0]  queue_dataOut_6_readFromScalar = _queue_fifo_6_data_out[64:33];
  wire [2:0]   queue_dataOut_6_segment = _queue_fifo_6_data_out[67:65];
  wire         queue_dataOut_6_mask = _queue_fifo_6_data_out[68];
  wire [1:0]   queue_dataOut_6_loadStoreEEW = _queue_fifo_6_data_out[70:69];
  wire [4:0]   queue_dataOut_6_vd = _queue_fifo_6_data_out[75:71];
  wire [4:0]   queue_dataOut_6_vs2 = _queue_fifo_6_data_out[80:76];
  wire [4:0]   queue_dataOut_6_vs1 = _queue_fifo_6_data_out[85:81];
  wire         queue_dataOut_6_lsWholeReg = _queue_fifo_6_data_out[86];
  wire         queue_dataOut_6_special = _queue_fifo_6_data_out[87];
  wire         queue_dataOut_6_store = _queue_fifo_6_data_out[88];
  wire         queue_dataOut_6_issueInst = _queue_fifo_6_data_out[89];
  wire         queue_dataOut_6_loadStore = _queue_fifo_6_data_out[90];
  wire         queue_dataOut_6_decodeResult_logic = _queue_fifo_6_data_out[91];
  wire         queue_dataOut_6_decodeResult_adder = _queue_fifo_6_data_out[92];
  wire         queue_dataOut_6_decodeResult_shift = _queue_fifo_6_data_out[93];
  wire         queue_dataOut_6_decodeResult_multiplier = _queue_fifo_6_data_out[94];
  wire         queue_dataOut_6_decodeResult_divider = _queue_fifo_6_data_out[95];
  wire         queue_dataOut_6_decodeResult_multiCycle = _queue_fifo_6_data_out[96];
  wire         queue_dataOut_6_decodeResult_other = _queue_fifo_6_data_out[97];
  wire         queue_dataOut_6_decodeResult_unsigned0 = _queue_fifo_6_data_out[98];
  wire         queue_dataOut_6_decodeResult_unsigned1 = _queue_fifo_6_data_out[99];
  wire         queue_dataOut_6_decodeResult_itype = _queue_fifo_6_data_out[100];
  wire         queue_dataOut_6_decodeResult_nr = _queue_fifo_6_data_out[101];
  wire         queue_dataOut_6_decodeResult_red = _queue_fifo_6_data_out[102];
  wire         queue_dataOut_6_decodeResult_widenReduce = _queue_fifo_6_data_out[103];
  wire         queue_dataOut_6_decodeResult_targetRd = _queue_fifo_6_data_out[104];
  wire         queue_dataOut_6_decodeResult_slid = _queue_fifo_6_data_out[105];
  wire         queue_dataOut_6_decodeResult_gather = _queue_fifo_6_data_out[106];
  wire         queue_dataOut_6_decodeResult_gather16 = _queue_fifo_6_data_out[107];
  wire         queue_dataOut_6_decodeResult_compress = _queue_fifo_6_data_out[108];
  wire         queue_dataOut_6_decodeResult_unOrderWrite = _queue_fifo_6_data_out[109];
  wire         queue_dataOut_6_decodeResult_extend = _queue_fifo_6_data_out[110];
  wire         queue_dataOut_6_decodeResult_mv = _queue_fifo_6_data_out[111];
  wire         queue_dataOut_6_decodeResult_iota = _queue_fifo_6_data_out[112];
  wire [3:0]   queue_dataOut_6_decodeResult_uop = _queue_fifo_6_data_out[116:113];
  wire         queue_dataOut_6_decodeResult_maskLogic = _queue_fifo_6_data_out[117];
  wire         queue_dataOut_6_decodeResult_maskDestination = _queue_fifo_6_data_out[118];
  wire         queue_dataOut_6_decodeResult_maskSource = _queue_fifo_6_data_out[119];
  wire         queue_dataOut_6_decodeResult_readOnly = _queue_fifo_6_data_out[120];
  wire         queue_dataOut_6_decodeResult_vwmacc = _queue_fifo_6_data_out[121];
  wire         queue_dataOut_6_decodeResult_saturate = _queue_fifo_6_data_out[122];
  wire         queue_dataOut_6_decodeResult_special = _queue_fifo_6_data_out[123];
  wire         queue_dataOut_6_decodeResult_maskUnit = _queue_fifo_6_data_out[124];
  wire         queue_dataOut_6_decodeResult_crossWrite = _queue_fifo_6_data_out[125];
  wire         queue_dataOut_6_decodeResult_crossRead = _queue_fifo_6_data_out[126];
  wire         queue_dataOut_6_decodeResult_sWrite = _queue_fifo_6_data_out[127];
  wire         queue_dataOut_6_decodeResult_vtype = _queue_fifo_6_data_out[128];
  wire         queue_dataOut_6_decodeResult_sReadVD = _queue_fifo_6_data_out[129];
  wire         queue_dataOut_6_decodeResult_scheduler = _queue_fifo_6_data_out[130];
  wire         queue_dataOut_6_decodeResult_dontNeedExecuteInLane = _queue_fifo_6_data_out[131];
  wire         queue_dataOut_6_decodeResult_reverse = _queue_fifo_6_data_out[132];
  wire         queue_dataOut_6_decodeResult_average = _queue_fifo_6_data_out[133];
  wire         queue_dataOut_6_decodeResult_ffo = _queue_fifo_6_data_out[134];
  wire         queue_dataOut_6_decodeResult_popCount = _queue_fifo_6_data_out[135];
  wire [4:0]   queue_dataOut_6_decodeResult_topUop = _queue_fifo_6_data_out[140:136];
  wire         queue_dataOut_6_decodeResult_specialSlot = _queue_fifo_6_data_out[141];
  wire         queue_dataOut_6_decodeResult_float = _queue_fifo_6_data_out[142];
  wire [1:0]   queue_dataOut_6_decodeResult_fpExecutionType = _queue_fifo_6_data_out[144:143];
  wire         queue_dataOut_6_decodeResult_floatMul = _queue_fifo_6_data_out[145];
  wire         queue_dataOut_6_decodeResult_orderReduce = _queue_fifo_6_data_out[146];
  wire [2:0]   queue_dataOut_6_instructionIndex = _queue_fifo_6_data_out[149:147];
  wire         queue_6_enq_ready = ~_queue_fifo_6_full;
  wire         queue_6_enq_valid;
  assign queue_6_deq_valid = ~_queue_fifo_6_empty | queue_6_enq_valid;
  assign queue_6_deq_bits_instructionIndex = _queue_fifo_6_empty ? queue_6_enq_bits_instructionIndex : queue_dataOut_6_instructionIndex;
  assign queue_6_deq_bits_decodeResult_orderReduce = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_orderReduce : queue_dataOut_6_decodeResult_orderReduce;
  assign queue_6_deq_bits_decodeResult_floatMul = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_floatMul : queue_dataOut_6_decodeResult_floatMul;
  assign queue_6_deq_bits_decodeResult_fpExecutionType = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_fpExecutionType : queue_dataOut_6_decodeResult_fpExecutionType;
  assign queue_6_deq_bits_decodeResult_float = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_float : queue_dataOut_6_decodeResult_float;
  assign queue_6_deq_bits_decodeResult_specialSlot = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_specialSlot : queue_dataOut_6_decodeResult_specialSlot;
  assign queue_6_deq_bits_decodeResult_topUop = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_topUop : queue_dataOut_6_decodeResult_topUop;
  assign queue_6_deq_bits_decodeResult_popCount = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_popCount : queue_dataOut_6_decodeResult_popCount;
  assign queue_6_deq_bits_decodeResult_ffo = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_ffo : queue_dataOut_6_decodeResult_ffo;
  assign queue_6_deq_bits_decodeResult_average = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_average : queue_dataOut_6_decodeResult_average;
  assign queue_6_deq_bits_decodeResult_reverse = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_reverse : queue_dataOut_6_decodeResult_reverse;
  assign queue_6_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_6_decodeResult_dontNeedExecuteInLane;
  assign queue_6_deq_bits_decodeResult_scheduler = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_scheduler : queue_dataOut_6_decodeResult_scheduler;
  assign queue_6_deq_bits_decodeResult_sReadVD = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_sReadVD : queue_dataOut_6_decodeResult_sReadVD;
  assign queue_6_deq_bits_decodeResult_vtype = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_vtype : queue_dataOut_6_decodeResult_vtype;
  assign queue_6_deq_bits_decodeResult_sWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_sWrite : queue_dataOut_6_decodeResult_sWrite;
  assign queue_6_deq_bits_decodeResult_crossRead = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_crossRead : queue_dataOut_6_decodeResult_crossRead;
  assign queue_6_deq_bits_decodeResult_crossWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_crossWrite : queue_dataOut_6_decodeResult_crossWrite;
  assign queue_6_deq_bits_decodeResult_maskUnit = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskUnit : queue_dataOut_6_decodeResult_maskUnit;
  assign queue_6_deq_bits_decodeResult_special = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_special : queue_dataOut_6_decodeResult_special;
  assign queue_6_deq_bits_decodeResult_saturate = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_saturate : queue_dataOut_6_decodeResult_saturate;
  assign queue_6_deq_bits_decodeResult_vwmacc = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_vwmacc : queue_dataOut_6_decodeResult_vwmacc;
  assign queue_6_deq_bits_decodeResult_readOnly = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_readOnly : queue_dataOut_6_decodeResult_readOnly;
  assign queue_6_deq_bits_decodeResult_maskSource = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskSource : queue_dataOut_6_decodeResult_maskSource;
  assign queue_6_deq_bits_decodeResult_maskDestination = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskDestination : queue_dataOut_6_decodeResult_maskDestination;
  assign queue_6_deq_bits_decodeResult_maskLogic = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskLogic : queue_dataOut_6_decodeResult_maskLogic;
  assign queue_6_deq_bits_decodeResult_uop = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_uop : queue_dataOut_6_decodeResult_uop;
  assign queue_6_deq_bits_decodeResult_iota = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_iota : queue_dataOut_6_decodeResult_iota;
  assign queue_6_deq_bits_decodeResult_mv = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_mv : queue_dataOut_6_decodeResult_mv;
  assign queue_6_deq_bits_decodeResult_extend = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_extend : queue_dataOut_6_decodeResult_extend;
  assign queue_6_deq_bits_decodeResult_unOrderWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unOrderWrite : queue_dataOut_6_decodeResult_unOrderWrite;
  assign queue_6_deq_bits_decodeResult_compress = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_compress : queue_dataOut_6_decodeResult_compress;
  assign queue_6_deq_bits_decodeResult_gather16 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_gather16 : queue_dataOut_6_decodeResult_gather16;
  assign queue_6_deq_bits_decodeResult_gather = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_gather : queue_dataOut_6_decodeResult_gather;
  assign queue_6_deq_bits_decodeResult_slid = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_slid : queue_dataOut_6_decodeResult_slid;
  assign queue_6_deq_bits_decodeResult_targetRd = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_targetRd : queue_dataOut_6_decodeResult_targetRd;
  assign queue_6_deq_bits_decodeResult_widenReduce = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_widenReduce : queue_dataOut_6_decodeResult_widenReduce;
  assign queue_6_deq_bits_decodeResult_red = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_red : queue_dataOut_6_decodeResult_red;
  assign queue_6_deq_bits_decodeResult_nr = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_nr : queue_dataOut_6_decodeResult_nr;
  assign queue_6_deq_bits_decodeResult_itype = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_itype : queue_dataOut_6_decodeResult_itype;
  assign queue_6_deq_bits_decodeResult_unsigned1 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unsigned1 : queue_dataOut_6_decodeResult_unsigned1;
  assign queue_6_deq_bits_decodeResult_unsigned0 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unsigned0 : queue_dataOut_6_decodeResult_unsigned0;
  assign queue_6_deq_bits_decodeResult_other = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_other : queue_dataOut_6_decodeResult_other;
  assign queue_6_deq_bits_decodeResult_multiCycle = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_multiCycle : queue_dataOut_6_decodeResult_multiCycle;
  assign queue_6_deq_bits_decodeResult_divider = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_divider : queue_dataOut_6_decodeResult_divider;
  assign queue_6_deq_bits_decodeResult_multiplier = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_multiplier : queue_dataOut_6_decodeResult_multiplier;
  assign queue_6_deq_bits_decodeResult_shift = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_shift : queue_dataOut_6_decodeResult_shift;
  assign queue_6_deq_bits_decodeResult_adder = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_adder : queue_dataOut_6_decodeResult_adder;
  assign queue_6_deq_bits_decodeResult_logic = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_logic : queue_dataOut_6_decodeResult_logic;
  assign queue_6_deq_bits_loadStore = _queue_fifo_6_empty ? queue_6_enq_bits_loadStore : queue_dataOut_6_loadStore;
  assign queue_6_deq_bits_issueInst = _queue_fifo_6_empty ? queue_6_enq_bits_issueInst : queue_dataOut_6_issueInst;
  assign queue_6_deq_bits_store = _queue_fifo_6_empty ? queue_6_enq_bits_store : queue_dataOut_6_store;
  assign queue_6_deq_bits_special = _queue_fifo_6_empty ? queue_6_enq_bits_special : queue_dataOut_6_special;
  assign queue_6_deq_bits_lsWholeReg = _queue_fifo_6_empty ? queue_6_enq_bits_lsWholeReg : queue_dataOut_6_lsWholeReg;
  assign queue_6_deq_bits_vs1 = _queue_fifo_6_empty ? queue_6_enq_bits_vs1 : queue_dataOut_6_vs1;
  assign queue_6_deq_bits_vs2 = _queue_fifo_6_empty ? queue_6_enq_bits_vs2 : queue_dataOut_6_vs2;
  assign queue_6_deq_bits_vd = _queue_fifo_6_empty ? queue_6_enq_bits_vd : queue_dataOut_6_vd;
  assign queue_6_deq_bits_loadStoreEEW = _queue_fifo_6_empty ? queue_6_enq_bits_loadStoreEEW : queue_dataOut_6_loadStoreEEW;
  assign queue_6_deq_bits_mask = _queue_fifo_6_empty ? queue_6_enq_bits_mask : queue_dataOut_6_mask;
  assign queue_6_deq_bits_segment = _queue_fifo_6_empty ? queue_6_enq_bits_segment : queue_dataOut_6_segment;
  assign queue_6_deq_bits_readFromScalar = _queue_fifo_6_empty ? queue_6_enq_bits_readFromScalar : queue_dataOut_6_readFromScalar;
  assign queue_6_deq_bits_csrInterface_vl = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vl : queue_dataOut_6_csrInterface_vl;
  assign queue_6_deq_bits_csrInterface_vStart = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vStart : queue_dataOut_6_csrInterface_vStart;
  assign queue_6_deq_bits_csrInterface_vlmul = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vlmul : queue_dataOut_6_csrInterface_vlmul;
  assign queue_6_deq_bits_csrInterface_vSew = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vSew : queue_dataOut_6_csrInterface_vSew;
  assign queue_6_deq_bits_csrInterface_vxrm = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vxrm : queue_dataOut_6_csrInterface_vxrm;
  assign queue_6_deq_bits_csrInterface_vta = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vta : queue_dataOut_6_csrInterface_vta;
  assign queue_6_deq_bits_csrInterface_vma = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vma : queue_dataOut_6_csrInterface_vma;
  wire         laneVec_6_laneRequest_bits_issueInst = laneRequestSinkWire_6_ready & laneRequestSinkWire_6_valid;
  reg          releasePipe_pipe_v_6;
  wire         releasePipe_pipe_out_6_valid = releasePipe_pipe_v_6;
  wire         laneRequestSourceWire_6_ready;
  wire         validSource_6_valid = laneRequestSourceWire_6_ready & laneRequestSourceWire_6_valid;
  reg  [2:0]   tokenCheck_counter_6;
  wire [2:0]   tokenCheck_counterChange_6 = validSource_6_valid ? 3'h1 : 3'h7;
  assign tokenCheck_6 = ~(tokenCheck_counter_6[2]);
  assign laneRequestSourceWire_6_ready = tokenCheck_6;
  assign queue_6_enq_valid = validSink_6_valid;
  assign queue_6_enq_bits_instructionIndex = validSink_6_bits_instructionIndex;
  assign queue_6_enq_bits_decodeResult_orderReduce = validSink_6_bits_decodeResult_orderReduce;
  assign queue_6_enq_bits_decodeResult_floatMul = validSink_6_bits_decodeResult_floatMul;
  assign queue_6_enq_bits_decodeResult_fpExecutionType = validSink_6_bits_decodeResult_fpExecutionType;
  assign queue_6_enq_bits_decodeResult_float = validSink_6_bits_decodeResult_float;
  assign queue_6_enq_bits_decodeResult_specialSlot = validSink_6_bits_decodeResult_specialSlot;
  assign queue_6_enq_bits_decodeResult_topUop = validSink_6_bits_decodeResult_topUop;
  assign queue_6_enq_bits_decodeResult_popCount = validSink_6_bits_decodeResult_popCount;
  assign queue_6_enq_bits_decodeResult_ffo = validSink_6_bits_decodeResult_ffo;
  assign queue_6_enq_bits_decodeResult_average = validSink_6_bits_decodeResult_average;
  assign queue_6_enq_bits_decodeResult_reverse = validSink_6_bits_decodeResult_reverse;
  assign queue_6_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_6_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_6_enq_bits_decodeResult_scheduler = validSink_6_bits_decodeResult_scheduler;
  assign queue_6_enq_bits_decodeResult_sReadVD = validSink_6_bits_decodeResult_sReadVD;
  assign queue_6_enq_bits_decodeResult_vtype = validSink_6_bits_decodeResult_vtype;
  assign queue_6_enq_bits_decodeResult_sWrite = validSink_6_bits_decodeResult_sWrite;
  assign queue_6_enq_bits_decodeResult_crossRead = validSink_6_bits_decodeResult_crossRead;
  assign queue_6_enq_bits_decodeResult_crossWrite = validSink_6_bits_decodeResult_crossWrite;
  assign queue_6_enq_bits_decodeResult_maskUnit = validSink_6_bits_decodeResult_maskUnit;
  assign queue_6_enq_bits_decodeResult_special = validSink_6_bits_decodeResult_special;
  assign queue_6_enq_bits_decodeResult_saturate = validSink_6_bits_decodeResult_saturate;
  assign queue_6_enq_bits_decodeResult_vwmacc = validSink_6_bits_decodeResult_vwmacc;
  assign queue_6_enq_bits_decodeResult_readOnly = validSink_6_bits_decodeResult_readOnly;
  assign queue_6_enq_bits_decodeResult_maskSource = validSink_6_bits_decodeResult_maskSource;
  assign queue_6_enq_bits_decodeResult_maskDestination = validSink_6_bits_decodeResult_maskDestination;
  assign queue_6_enq_bits_decodeResult_maskLogic = validSink_6_bits_decodeResult_maskLogic;
  assign queue_6_enq_bits_decodeResult_uop = validSink_6_bits_decodeResult_uop;
  assign queue_6_enq_bits_decodeResult_iota = validSink_6_bits_decodeResult_iota;
  assign queue_6_enq_bits_decodeResult_mv = validSink_6_bits_decodeResult_mv;
  assign queue_6_enq_bits_decodeResult_extend = validSink_6_bits_decodeResult_extend;
  assign queue_6_enq_bits_decodeResult_unOrderWrite = validSink_6_bits_decodeResult_unOrderWrite;
  assign queue_6_enq_bits_decodeResult_compress = validSink_6_bits_decodeResult_compress;
  assign queue_6_enq_bits_decodeResult_gather16 = validSink_6_bits_decodeResult_gather16;
  assign queue_6_enq_bits_decodeResult_gather = validSink_6_bits_decodeResult_gather;
  assign queue_6_enq_bits_decodeResult_slid = validSink_6_bits_decodeResult_slid;
  assign queue_6_enq_bits_decodeResult_targetRd = validSink_6_bits_decodeResult_targetRd;
  assign queue_6_enq_bits_decodeResult_widenReduce = validSink_6_bits_decodeResult_widenReduce;
  assign queue_6_enq_bits_decodeResult_red = validSink_6_bits_decodeResult_red;
  assign queue_6_enq_bits_decodeResult_nr = validSink_6_bits_decodeResult_nr;
  assign queue_6_enq_bits_decodeResult_itype = validSink_6_bits_decodeResult_itype;
  assign queue_6_enq_bits_decodeResult_unsigned1 = validSink_6_bits_decodeResult_unsigned1;
  assign queue_6_enq_bits_decodeResult_unsigned0 = validSink_6_bits_decodeResult_unsigned0;
  assign queue_6_enq_bits_decodeResult_other = validSink_6_bits_decodeResult_other;
  assign queue_6_enq_bits_decodeResult_multiCycle = validSink_6_bits_decodeResult_multiCycle;
  assign queue_6_enq_bits_decodeResult_divider = validSink_6_bits_decodeResult_divider;
  assign queue_6_enq_bits_decodeResult_multiplier = validSink_6_bits_decodeResult_multiplier;
  assign queue_6_enq_bits_decodeResult_shift = validSink_6_bits_decodeResult_shift;
  assign queue_6_enq_bits_decodeResult_adder = validSink_6_bits_decodeResult_adder;
  assign queue_6_enq_bits_decodeResult_logic = validSink_6_bits_decodeResult_logic;
  assign queue_6_enq_bits_loadStore = validSink_6_bits_loadStore;
  assign queue_6_enq_bits_issueInst = validSink_6_bits_issueInst;
  assign queue_6_enq_bits_store = validSink_6_bits_store;
  assign queue_6_enq_bits_special = validSink_6_bits_special;
  assign queue_6_enq_bits_lsWholeReg = validSink_6_bits_lsWholeReg;
  assign queue_6_enq_bits_vs1 = validSink_6_bits_vs1;
  assign queue_6_enq_bits_vs2 = validSink_6_bits_vs2;
  assign queue_6_enq_bits_vd = validSink_6_bits_vd;
  assign queue_6_enq_bits_loadStoreEEW = validSink_6_bits_loadStoreEEW;
  assign queue_6_enq_bits_mask = validSink_6_bits_mask;
  assign queue_6_enq_bits_segment = validSink_6_bits_segment;
  assign queue_6_enq_bits_readFromScalar = validSink_6_bits_readFromScalar;
  assign queue_6_enq_bits_csrInterface_vl = validSink_6_bits_csrInterface_vl;
  assign queue_6_enq_bits_csrInterface_vStart = validSink_6_bits_csrInterface_vStart;
  assign queue_6_enq_bits_csrInterface_vlmul = validSink_6_bits_csrInterface_vlmul;
  assign queue_6_enq_bits_csrInterface_vSew = validSink_6_bits_csrInterface_vSew;
  assign queue_6_enq_bits_csrInterface_vxrm = validSink_6_bits_csrInterface_vxrm;
  assign queue_6_enq_bits_csrInterface_vta = validSink_6_bits_csrInterface_vta;
  assign queue_6_enq_bits_csrInterface_vma = validSink_6_bits_csrInterface_vma;
  reg          shifterReg_6_0_valid;
  assign validSink_6_valid = shifterReg_6_0_valid;
  reg  [2:0]   shifterReg_6_0_bits_instructionIndex;
  assign validSink_6_bits_instructionIndex = shifterReg_6_0_bits_instructionIndex;
  reg          shifterReg_6_0_bits_decodeResult_orderReduce;
  assign validSink_6_bits_decodeResult_orderReduce = shifterReg_6_0_bits_decodeResult_orderReduce;
  reg          shifterReg_6_0_bits_decodeResult_floatMul;
  assign validSink_6_bits_decodeResult_floatMul = shifterReg_6_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_6_0_bits_decodeResult_fpExecutionType;
  assign validSink_6_bits_decodeResult_fpExecutionType = shifterReg_6_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_6_0_bits_decodeResult_float;
  assign validSink_6_bits_decodeResult_float = shifterReg_6_0_bits_decodeResult_float;
  reg          shifterReg_6_0_bits_decodeResult_specialSlot;
  assign validSink_6_bits_decodeResult_specialSlot = shifterReg_6_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_6_0_bits_decodeResult_topUop;
  assign validSink_6_bits_decodeResult_topUop = shifterReg_6_0_bits_decodeResult_topUop;
  reg          shifterReg_6_0_bits_decodeResult_popCount;
  assign validSink_6_bits_decodeResult_popCount = shifterReg_6_0_bits_decodeResult_popCount;
  reg          shifterReg_6_0_bits_decodeResult_ffo;
  assign validSink_6_bits_decodeResult_ffo = shifterReg_6_0_bits_decodeResult_ffo;
  reg          shifterReg_6_0_bits_decodeResult_average;
  assign validSink_6_bits_decodeResult_average = shifterReg_6_0_bits_decodeResult_average;
  reg          shifterReg_6_0_bits_decodeResult_reverse;
  assign validSink_6_bits_decodeResult_reverse = shifterReg_6_0_bits_decodeResult_reverse;
  reg          shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_6_bits_decodeResult_dontNeedExecuteInLane = shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_6_0_bits_decodeResult_scheduler;
  assign validSink_6_bits_decodeResult_scheduler = shifterReg_6_0_bits_decodeResult_scheduler;
  reg          shifterReg_6_0_bits_decodeResult_sReadVD;
  assign validSink_6_bits_decodeResult_sReadVD = shifterReg_6_0_bits_decodeResult_sReadVD;
  reg          shifterReg_6_0_bits_decodeResult_vtype;
  assign validSink_6_bits_decodeResult_vtype = shifterReg_6_0_bits_decodeResult_vtype;
  reg          shifterReg_6_0_bits_decodeResult_sWrite;
  assign validSink_6_bits_decodeResult_sWrite = shifterReg_6_0_bits_decodeResult_sWrite;
  reg          shifterReg_6_0_bits_decodeResult_crossRead;
  assign validSink_6_bits_decodeResult_crossRead = shifterReg_6_0_bits_decodeResult_crossRead;
  reg          shifterReg_6_0_bits_decodeResult_crossWrite;
  assign validSink_6_bits_decodeResult_crossWrite = shifterReg_6_0_bits_decodeResult_crossWrite;
  reg          shifterReg_6_0_bits_decodeResult_maskUnit;
  assign validSink_6_bits_decodeResult_maskUnit = shifterReg_6_0_bits_decodeResult_maskUnit;
  reg          shifterReg_6_0_bits_decodeResult_special;
  assign validSink_6_bits_decodeResult_special = shifterReg_6_0_bits_decodeResult_special;
  reg          shifterReg_6_0_bits_decodeResult_saturate;
  assign validSink_6_bits_decodeResult_saturate = shifterReg_6_0_bits_decodeResult_saturate;
  reg          shifterReg_6_0_bits_decodeResult_vwmacc;
  assign validSink_6_bits_decodeResult_vwmacc = shifterReg_6_0_bits_decodeResult_vwmacc;
  reg          shifterReg_6_0_bits_decodeResult_readOnly;
  assign validSink_6_bits_decodeResult_readOnly = shifterReg_6_0_bits_decodeResult_readOnly;
  reg          shifterReg_6_0_bits_decodeResult_maskSource;
  assign validSink_6_bits_decodeResult_maskSource = shifterReg_6_0_bits_decodeResult_maskSource;
  reg          shifterReg_6_0_bits_decodeResult_maskDestination;
  assign validSink_6_bits_decodeResult_maskDestination = shifterReg_6_0_bits_decodeResult_maskDestination;
  reg          shifterReg_6_0_bits_decodeResult_maskLogic;
  assign validSink_6_bits_decodeResult_maskLogic = shifterReg_6_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_6_0_bits_decodeResult_uop;
  assign validSink_6_bits_decodeResult_uop = shifterReg_6_0_bits_decodeResult_uop;
  reg          shifterReg_6_0_bits_decodeResult_iota;
  assign validSink_6_bits_decodeResult_iota = shifterReg_6_0_bits_decodeResult_iota;
  reg          shifterReg_6_0_bits_decodeResult_mv;
  assign validSink_6_bits_decodeResult_mv = shifterReg_6_0_bits_decodeResult_mv;
  reg          shifterReg_6_0_bits_decodeResult_extend;
  assign validSink_6_bits_decodeResult_extend = shifterReg_6_0_bits_decodeResult_extend;
  reg          shifterReg_6_0_bits_decodeResult_unOrderWrite;
  assign validSink_6_bits_decodeResult_unOrderWrite = shifterReg_6_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_6_0_bits_decodeResult_compress;
  assign validSink_6_bits_decodeResult_compress = shifterReg_6_0_bits_decodeResult_compress;
  reg          shifterReg_6_0_bits_decodeResult_gather16;
  assign validSink_6_bits_decodeResult_gather16 = shifterReg_6_0_bits_decodeResult_gather16;
  reg          shifterReg_6_0_bits_decodeResult_gather;
  assign validSink_6_bits_decodeResult_gather = shifterReg_6_0_bits_decodeResult_gather;
  reg          shifterReg_6_0_bits_decodeResult_slid;
  assign validSink_6_bits_decodeResult_slid = shifterReg_6_0_bits_decodeResult_slid;
  reg          shifterReg_6_0_bits_decodeResult_targetRd;
  assign validSink_6_bits_decodeResult_targetRd = shifterReg_6_0_bits_decodeResult_targetRd;
  reg          shifterReg_6_0_bits_decodeResult_widenReduce;
  assign validSink_6_bits_decodeResult_widenReduce = shifterReg_6_0_bits_decodeResult_widenReduce;
  reg          shifterReg_6_0_bits_decodeResult_red;
  assign validSink_6_bits_decodeResult_red = shifterReg_6_0_bits_decodeResult_red;
  reg          shifterReg_6_0_bits_decodeResult_nr;
  assign validSink_6_bits_decodeResult_nr = shifterReg_6_0_bits_decodeResult_nr;
  reg          shifterReg_6_0_bits_decodeResult_itype;
  assign validSink_6_bits_decodeResult_itype = shifterReg_6_0_bits_decodeResult_itype;
  reg          shifterReg_6_0_bits_decodeResult_unsigned1;
  assign validSink_6_bits_decodeResult_unsigned1 = shifterReg_6_0_bits_decodeResult_unsigned1;
  reg          shifterReg_6_0_bits_decodeResult_unsigned0;
  assign validSink_6_bits_decodeResult_unsigned0 = shifterReg_6_0_bits_decodeResult_unsigned0;
  reg          shifterReg_6_0_bits_decodeResult_other;
  assign validSink_6_bits_decodeResult_other = shifterReg_6_0_bits_decodeResult_other;
  reg          shifterReg_6_0_bits_decodeResult_multiCycle;
  assign validSink_6_bits_decodeResult_multiCycle = shifterReg_6_0_bits_decodeResult_multiCycle;
  reg          shifterReg_6_0_bits_decodeResult_divider;
  assign validSink_6_bits_decodeResult_divider = shifterReg_6_0_bits_decodeResult_divider;
  reg          shifterReg_6_0_bits_decodeResult_multiplier;
  assign validSink_6_bits_decodeResult_multiplier = shifterReg_6_0_bits_decodeResult_multiplier;
  reg          shifterReg_6_0_bits_decodeResult_shift;
  assign validSink_6_bits_decodeResult_shift = shifterReg_6_0_bits_decodeResult_shift;
  reg          shifterReg_6_0_bits_decodeResult_adder;
  assign validSink_6_bits_decodeResult_adder = shifterReg_6_0_bits_decodeResult_adder;
  reg          shifterReg_6_0_bits_decodeResult_logic;
  assign validSink_6_bits_decodeResult_logic = shifterReg_6_0_bits_decodeResult_logic;
  reg          shifterReg_6_0_bits_loadStore;
  assign validSink_6_bits_loadStore = shifterReg_6_0_bits_loadStore;
  reg          shifterReg_6_0_bits_issueInst;
  assign validSink_6_bits_issueInst = shifterReg_6_0_bits_issueInst;
  reg          shifterReg_6_0_bits_store;
  assign validSink_6_bits_store = shifterReg_6_0_bits_store;
  reg          shifterReg_6_0_bits_special;
  assign validSink_6_bits_special = shifterReg_6_0_bits_special;
  reg          shifterReg_6_0_bits_lsWholeReg;
  assign validSink_6_bits_lsWholeReg = shifterReg_6_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_6_0_bits_vs1;
  assign validSink_6_bits_vs1 = shifterReg_6_0_bits_vs1;
  reg  [4:0]   shifterReg_6_0_bits_vs2;
  assign validSink_6_bits_vs2 = shifterReg_6_0_bits_vs2;
  reg  [4:0]   shifterReg_6_0_bits_vd;
  assign validSink_6_bits_vd = shifterReg_6_0_bits_vd;
  reg  [1:0]   shifterReg_6_0_bits_loadStoreEEW;
  assign validSink_6_bits_loadStoreEEW = shifterReg_6_0_bits_loadStoreEEW;
  reg          shifterReg_6_0_bits_mask;
  assign validSink_6_bits_mask = shifterReg_6_0_bits_mask;
  reg  [2:0]   shifterReg_6_0_bits_segment;
  assign validSink_6_bits_segment = shifterReg_6_0_bits_segment;
  reg  [31:0]  shifterReg_6_0_bits_readFromScalar;
  assign validSink_6_bits_readFromScalar = shifterReg_6_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_6_0_bits_csrInterface_vl;
  assign validSink_6_bits_csrInterface_vl = shifterReg_6_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_6_0_bits_csrInterface_vStart;
  assign validSink_6_bits_csrInterface_vStart = shifterReg_6_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_6_0_bits_csrInterface_vlmul;
  assign validSink_6_bits_csrInterface_vlmul = shifterReg_6_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_6_0_bits_csrInterface_vSew;
  assign validSink_6_bits_csrInterface_vSew = shifterReg_6_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_6_0_bits_csrInterface_vxrm;
  assign validSink_6_bits_csrInterface_vxrm = shifterReg_6_0_bits_csrInterface_vxrm;
  reg          shifterReg_6_0_bits_csrInterface_vta;
  assign validSink_6_bits_csrInterface_vta = shifterReg_6_0_bits_csrInterface_vta;
  reg          shifterReg_6_0_bits_csrInterface_vma;
  assign validSink_6_bits_csrInterface_vma = shifterReg_6_0_bits_csrInterface_vma;
  wire         shifterValid_6 = shifterReg_6_0_valid | validSource_6_valid;
  wire         validSink_7_valid;
  wire [2:0]   validSink_7_bits_instructionIndex;
  wire         validSink_7_bits_decodeResult_orderReduce;
  wire         validSink_7_bits_decodeResult_floatMul;
  wire [1:0]   validSink_7_bits_decodeResult_fpExecutionType;
  wire         validSink_7_bits_decodeResult_float;
  wire         validSink_7_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_7_bits_decodeResult_topUop;
  wire         validSink_7_bits_decodeResult_popCount;
  wire         validSink_7_bits_decodeResult_ffo;
  wire         validSink_7_bits_decodeResult_average;
  wire         validSink_7_bits_decodeResult_reverse;
  wire         validSink_7_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_7_bits_decodeResult_scheduler;
  wire         validSink_7_bits_decodeResult_sReadVD;
  wire         validSink_7_bits_decodeResult_vtype;
  wire         validSink_7_bits_decodeResult_sWrite;
  wire         validSink_7_bits_decodeResult_crossRead;
  wire         validSink_7_bits_decodeResult_crossWrite;
  wire         validSink_7_bits_decodeResult_maskUnit;
  wire         validSink_7_bits_decodeResult_special;
  wire         validSink_7_bits_decodeResult_saturate;
  wire         validSink_7_bits_decodeResult_vwmacc;
  wire         validSink_7_bits_decodeResult_readOnly;
  wire         validSink_7_bits_decodeResult_maskSource;
  wire         validSink_7_bits_decodeResult_maskDestination;
  wire         validSink_7_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_7_bits_decodeResult_uop;
  wire         validSink_7_bits_decodeResult_iota;
  wire         validSink_7_bits_decodeResult_mv;
  wire         validSink_7_bits_decodeResult_extend;
  wire         validSink_7_bits_decodeResult_unOrderWrite;
  wire         validSink_7_bits_decodeResult_compress;
  wire         validSink_7_bits_decodeResult_gather16;
  wire         validSink_7_bits_decodeResult_gather;
  wire         validSink_7_bits_decodeResult_slid;
  wire         validSink_7_bits_decodeResult_targetRd;
  wire         validSink_7_bits_decodeResult_widenReduce;
  wire         validSink_7_bits_decodeResult_red;
  wire         validSink_7_bits_decodeResult_nr;
  wire         validSink_7_bits_decodeResult_itype;
  wire         validSink_7_bits_decodeResult_unsigned1;
  wire         validSink_7_bits_decodeResult_unsigned0;
  wire         validSink_7_bits_decodeResult_other;
  wire         validSink_7_bits_decodeResult_multiCycle;
  wire         validSink_7_bits_decodeResult_divider;
  wire         validSink_7_bits_decodeResult_multiplier;
  wire         validSink_7_bits_decodeResult_shift;
  wire         validSink_7_bits_decodeResult_adder;
  wire         validSink_7_bits_decodeResult_logic;
  wire         validSink_7_bits_loadStore;
  wire         validSink_7_bits_issueInst;
  wire         validSink_7_bits_store;
  wire         validSink_7_bits_special;
  wire         validSink_7_bits_lsWholeReg;
  wire [4:0]   validSink_7_bits_vs1;
  wire [4:0]   validSink_7_bits_vs2;
  wire [4:0]   validSink_7_bits_vd;
  wire [1:0]   validSink_7_bits_loadStoreEEW;
  wire         validSink_7_bits_mask;
  wire [2:0]   validSink_7_bits_segment;
  wire [31:0]  validSink_7_bits_readFromScalar;
  wire [11:0]  validSink_7_bits_csrInterface_vl;
  wire [11:0]  validSink_7_bits_csrInterface_vStart;
  wire [2:0]   validSink_7_bits_csrInterface_vlmul;
  wire [1:0]   validSink_7_bits_csrInterface_vSew;
  wire [1:0]   validSink_7_bits_csrInterface_vxrm;
  wire         validSink_7_bits_csrInterface_vta;
  wire         validSink_7_bits_csrInterface_vma;
  wire         laneRequestSinkWire_7_valid = queue_7_deq_valid;
  wire [2:0]   laneRequestSinkWire_7_bits_instructionIndex = queue_7_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_7_bits_decodeResult_orderReduce = queue_7_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_7_bits_decodeResult_floatMul = queue_7_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_7_bits_decodeResult_fpExecutionType = queue_7_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_7_bits_decodeResult_float = queue_7_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_7_bits_decodeResult_specialSlot = queue_7_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_7_bits_decodeResult_topUop = queue_7_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_7_bits_decodeResult_popCount = queue_7_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_7_bits_decodeResult_ffo = queue_7_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_7_bits_decodeResult_average = queue_7_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_7_bits_decodeResult_reverse = queue_7_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_7_bits_decodeResult_dontNeedExecuteInLane = queue_7_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_7_bits_decodeResult_scheduler = queue_7_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_7_bits_decodeResult_sReadVD = queue_7_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_7_bits_decodeResult_vtype = queue_7_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_7_bits_decodeResult_sWrite = queue_7_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_crossRead = queue_7_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_7_bits_decodeResult_crossWrite = queue_7_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskUnit = queue_7_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_7_bits_decodeResult_special = queue_7_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_7_bits_decodeResult_saturate = queue_7_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_7_bits_decodeResult_vwmacc = queue_7_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_7_bits_decodeResult_readOnly = queue_7_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskSource = queue_7_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskDestination = queue_7_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskLogic = queue_7_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_7_bits_decodeResult_uop = queue_7_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_7_bits_decodeResult_iota = queue_7_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_7_bits_decodeResult_mv = queue_7_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_7_bits_decodeResult_extend = queue_7_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_7_bits_decodeResult_unOrderWrite = queue_7_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_compress = queue_7_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_7_bits_decodeResult_gather16 = queue_7_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_7_bits_decodeResult_gather = queue_7_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_7_bits_decodeResult_slid = queue_7_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_7_bits_decodeResult_targetRd = queue_7_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_7_bits_decodeResult_widenReduce = queue_7_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_7_bits_decodeResult_red = queue_7_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_7_bits_decodeResult_nr = queue_7_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_7_bits_decodeResult_itype = queue_7_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_7_bits_decodeResult_unsigned1 = queue_7_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_7_bits_decodeResult_unsigned0 = queue_7_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_7_bits_decodeResult_other = queue_7_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_7_bits_decodeResult_multiCycle = queue_7_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_7_bits_decodeResult_divider = queue_7_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_7_bits_decodeResult_multiplier = queue_7_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_7_bits_decodeResult_shift = queue_7_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_7_bits_decodeResult_adder = queue_7_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_7_bits_decodeResult_logic = queue_7_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_7_bits_loadStore = queue_7_deq_bits_loadStore;
  wire         laneRequestSinkWire_7_bits_issueInst = queue_7_deq_bits_issueInst;
  wire         laneRequestSinkWire_7_bits_store = queue_7_deq_bits_store;
  wire         laneRequestSinkWire_7_bits_special = queue_7_deq_bits_special;
  wire         laneRequestSinkWire_7_bits_lsWholeReg = queue_7_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_7_bits_vs1 = queue_7_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_7_bits_vs2 = queue_7_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_7_bits_vd = queue_7_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_7_bits_loadStoreEEW = queue_7_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_7_bits_mask = queue_7_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_7_bits_segment = queue_7_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_7_bits_readFromScalar = queue_7_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_7_bits_csrInterface_vl = queue_7_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_7_bits_csrInterface_vStart = queue_7_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_7_bits_csrInterface_vlmul = queue_7_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_7_bits_csrInterface_vSew = queue_7_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_7_bits_csrInterface_vxrm = queue_7_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_7_bits_csrInterface_vta = queue_7_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_7_bits_csrInterface_vma = queue_7_deq_bits_csrInterface_vma;
  wire [1:0]   queue_7_enq_bits_csrInterface_vxrm;
  wire         queue_7_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_21 = {queue_7_enq_bits_csrInterface_vxrm, queue_7_enq_bits_csrInterface_vta};
  wire         queue_7_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_21 = {queue_dataIn_lo_hi_21, queue_7_enq_bits_csrInterface_vma};
  wire [2:0]   queue_7_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_7_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_21 = {queue_7_enq_bits_csrInterface_vlmul, queue_7_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_7_enq_bits_csrInterface_vl;
  wire [11:0]  queue_7_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_21 = {queue_7_enq_bits_csrInterface_vl, queue_7_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_21 = {queue_dataIn_hi_hi_21, queue_dataIn_hi_lo_21};
  wire         queue_7_enq_bits_decodeResult_shift;
  wire         queue_7_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_7 = {queue_7_enq_bits_decodeResult_shift, queue_7_enq_bits_decodeResult_adder};
  wire         queue_7_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_7 = {queue_dataIn_lo_lo_lo_lo_hi_7, queue_7_enq_bits_decodeResult_logic};
  wire         queue_7_enq_bits_decodeResult_multiCycle;
  wire         queue_7_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_multiCycle, queue_7_enq_bits_decodeResult_divider};
  wire         queue_7_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_7 = {queue_dataIn_lo_lo_lo_hi_hi_7, queue_7_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_7 = {queue_dataIn_lo_lo_lo_hi_7, queue_dataIn_lo_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_unsigned1;
  wire         queue_7_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_unsigned1, queue_7_enq_bits_decodeResult_unsigned0};
  wire         queue_7_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_7 = {queue_dataIn_lo_lo_hi_lo_hi_7, queue_7_enq_bits_decodeResult_other};
  wire         queue_7_enq_bits_decodeResult_red;
  wire         queue_7_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_red, queue_7_enq_bits_decodeResult_nr};
  wire         queue_7_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_7 = {queue_dataIn_lo_lo_hi_hi_hi_7, queue_7_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_14 = {queue_dataIn_lo_lo_hi_hi_7, queue_dataIn_lo_lo_hi_lo_7};
  wire [11:0]  queue_dataIn_lo_lo_14 = {queue_dataIn_lo_lo_hi_14, queue_dataIn_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_slid;
  wire         queue_7_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_7 = {queue_7_enq_bits_decodeResult_slid, queue_7_enq_bits_decodeResult_targetRd};
  wire         queue_7_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_7 = {queue_dataIn_lo_hi_lo_lo_hi_7, queue_7_enq_bits_decodeResult_widenReduce};
  wire         queue_7_enq_bits_decodeResult_compress;
  wire         queue_7_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_compress, queue_7_enq_bits_decodeResult_gather16};
  wire         queue_7_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_7 = {queue_dataIn_lo_hi_lo_hi_hi_7, queue_7_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_14 = {queue_dataIn_lo_hi_lo_hi_7, queue_dataIn_lo_hi_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_mv;
  wire         queue_7_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_mv, queue_7_enq_bits_decodeResult_extend};
  wire         queue_7_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_7 = {queue_dataIn_lo_hi_hi_lo_hi_7, queue_7_enq_bits_decodeResult_unOrderWrite};
  wire         queue_7_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_7_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_maskLogic, queue_7_enq_bits_decodeResult_uop};
  wire         queue_7_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_7 = {queue_dataIn_lo_hi_hi_hi_hi_7, queue_7_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_14 = {queue_dataIn_lo_hi_hi_hi_7, queue_dataIn_lo_hi_hi_lo_7};
  wire [14:0]  queue_dataIn_lo_hi_22 = {queue_dataIn_lo_hi_hi_14, queue_dataIn_lo_hi_lo_14};
  wire [26:0]  queue_dataIn_lo_22 = {queue_dataIn_lo_hi_22, queue_dataIn_lo_lo_14};
  wire         queue_7_enq_bits_decodeResult_readOnly;
  wire         queue_7_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_7 = {queue_7_enq_bits_decodeResult_readOnly, queue_7_enq_bits_decodeResult_maskSource};
  wire         queue_7_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_7 = {queue_dataIn_hi_lo_lo_lo_hi_7, queue_7_enq_bits_decodeResult_maskDestination};
  wire         queue_7_enq_bits_decodeResult_special;
  wire         queue_7_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_special, queue_7_enq_bits_decodeResult_saturate};
  wire         queue_7_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_7 = {queue_dataIn_hi_lo_lo_hi_hi_7, queue_7_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_14 = {queue_dataIn_hi_lo_lo_hi_7, queue_dataIn_hi_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_crossRead;
  wire         queue_7_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_crossRead, queue_7_enq_bits_decodeResult_crossWrite};
  wire         queue_7_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_7 = {queue_dataIn_hi_lo_hi_lo_hi_7, queue_7_enq_bits_decodeResult_maskUnit};
  wire         queue_7_enq_bits_decodeResult_sReadVD;
  wire         queue_7_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_sReadVD, queue_7_enq_bits_decodeResult_vtype};
  wire         queue_7_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_7 = {queue_dataIn_hi_lo_hi_hi_hi_7, queue_7_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_14 = {queue_dataIn_hi_lo_hi_hi_7, queue_dataIn_hi_lo_hi_lo_7};
  wire [11:0]  queue_dataIn_hi_lo_22 = {queue_dataIn_hi_lo_hi_14, queue_dataIn_hi_lo_lo_14};
  wire         queue_7_enq_bits_decodeResult_reverse;
  wire         queue_7_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_7 = {queue_7_enq_bits_decodeResult_reverse, queue_7_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_7_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_7 = {queue_dataIn_hi_hi_lo_lo_hi_7, queue_7_enq_bits_decodeResult_scheduler};
  wire         queue_7_enq_bits_decodeResult_popCount;
  wire         queue_7_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_popCount, queue_7_enq_bits_decodeResult_ffo};
  wire         queue_7_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_7 = {queue_dataIn_hi_hi_lo_hi_hi_7, queue_7_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_14 = {queue_dataIn_hi_hi_lo_hi_7, queue_dataIn_hi_hi_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_float;
  wire         queue_7_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_float, queue_7_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_7_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_7 = {queue_dataIn_hi_hi_hi_lo_hi_7, queue_7_enq_bits_decodeResult_topUop};
  wire         queue_7_enq_bits_decodeResult_orderReduce;
  wire         queue_7_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_orderReduce, queue_7_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_7_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_7 = {queue_dataIn_hi_hi_hi_hi_hi_7, queue_7_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_14 = {queue_dataIn_hi_hi_hi_hi_7, queue_dataIn_hi_hi_hi_lo_7};
  wire [16:0]  queue_dataIn_hi_hi_22 = {queue_dataIn_hi_hi_hi_14, queue_dataIn_hi_hi_lo_14};
  wire [28:0]  queue_dataIn_hi_22 = {queue_dataIn_hi_hi_22, queue_dataIn_hi_lo_22};
  wire [2:0]   queue_7_enq_bits_segment;
  wire [31:0]  queue_7_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_15 = {queue_7_enq_bits_segment, queue_7_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_15 = {queue_dataIn_lo_lo_hi_15, queue_dataIn_hi_21, queue_dataIn_lo_21};
  wire [1:0]   queue_7_enq_bits_loadStoreEEW;
  wire         queue_7_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_15 = {queue_7_enq_bits_loadStoreEEW, queue_7_enq_bits_mask};
  wire [4:0]   queue_7_enq_bits_vs2;
  wire [4:0]   queue_7_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_15 = {queue_7_enq_bits_vs2, queue_7_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_23 = {queue_dataIn_lo_hi_hi_15, queue_dataIn_lo_hi_lo_15};
  wire [80:0]  queue_dataIn_lo_23 = {queue_dataIn_lo_hi_23, queue_dataIn_lo_lo_15};
  wire         queue_7_enq_bits_lsWholeReg;
  wire [4:0]   queue_7_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_15 = {queue_7_enq_bits_lsWholeReg, queue_7_enq_bits_vs1};
  wire         queue_7_enq_bits_store;
  wire         queue_7_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_15 = {queue_7_enq_bits_store, queue_7_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_23 = {queue_dataIn_hi_lo_hi_15, queue_dataIn_hi_lo_lo_15};
  wire         queue_7_enq_bits_loadStore;
  wire         queue_7_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_15 = {queue_7_enq_bits_loadStore, queue_7_enq_bits_issueInst};
  wire [2:0]   queue_7_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_15 = {queue_7_enq_bits_instructionIndex, queue_dataIn_hi_22, queue_dataIn_lo_22};
  wire [60:0]  queue_dataIn_hi_hi_23 = {queue_dataIn_hi_hi_hi_15, queue_dataIn_hi_hi_lo_15};
  wire [68:0]  queue_dataIn_hi_23 = {queue_dataIn_hi_hi_23, queue_dataIn_hi_lo_23};
  wire [149:0] queue_dataIn_7 = {queue_dataIn_hi_23, queue_dataIn_lo_23};
  wire         queue_dataOut_7_csrInterface_vma = _queue_fifo_7_data_out[0];
  wire         queue_dataOut_7_csrInterface_vta = _queue_fifo_7_data_out[1];
  wire [1:0]   queue_dataOut_7_csrInterface_vxrm = _queue_fifo_7_data_out[3:2];
  wire [1:0]   queue_dataOut_7_csrInterface_vSew = _queue_fifo_7_data_out[5:4];
  wire [2:0]   queue_dataOut_7_csrInterface_vlmul = _queue_fifo_7_data_out[8:6];
  wire [11:0]  queue_dataOut_7_csrInterface_vStart = _queue_fifo_7_data_out[20:9];
  wire [11:0]  queue_dataOut_7_csrInterface_vl = _queue_fifo_7_data_out[32:21];
  wire [31:0]  queue_dataOut_7_readFromScalar = _queue_fifo_7_data_out[64:33];
  wire [2:0]   queue_dataOut_7_segment = _queue_fifo_7_data_out[67:65];
  wire         queue_dataOut_7_mask = _queue_fifo_7_data_out[68];
  wire [1:0]   queue_dataOut_7_loadStoreEEW = _queue_fifo_7_data_out[70:69];
  wire [4:0]   queue_dataOut_7_vd = _queue_fifo_7_data_out[75:71];
  wire [4:0]   queue_dataOut_7_vs2 = _queue_fifo_7_data_out[80:76];
  wire [4:0]   queue_dataOut_7_vs1 = _queue_fifo_7_data_out[85:81];
  wire         queue_dataOut_7_lsWholeReg = _queue_fifo_7_data_out[86];
  wire         queue_dataOut_7_special = _queue_fifo_7_data_out[87];
  wire         queue_dataOut_7_store = _queue_fifo_7_data_out[88];
  wire         queue_dataOut_7_issueInst = _queue_fifo_7_data_out[89];
  wire         queue_dataOut_7_loadStore = _queue_fifo_7_data_out[90];
  wire         queue_dataOut_7_decodeResult_logic = _queue_fifo_7_data_out[91];
  wire         queue_dataOut_7_decodeResult_adder = _queue_fifo_7_data_out[92];
  wire         queue_dataOut_7_decodeResult_shift = _queue_fifo_7_data_out[93];
  wire         queue_dataOut_7_decodeResult_multiplier = _queue_fifo_7_data_out[94];
  wire         queue_dataOut_7_decodeResult_divider = _queue_fifo_7_data_out[95];
  wire         queue_dataOut_7_decodeResult_multiCycle = _queue_fifo_7_data_out[96];
  wire         queue_dataOut_7_decodeResult_other = _queue_fifo_7_data_out[97];
  wire         queue_dataOut_7_decodeResult_unsigned0 = _queue_fifo_7_data_out[98];
  wire         queue_dataOut_7_decodeResult_unsigned1 = _queue_fifo_7_data_out[99];
  wire         queue_dataOut_7_decodeResult_itype = _queue_fifo_7_data_out[100];
  wire         queue_dataOut_7_decodeResult_nr = _queue_fifo_7_data_out[101];
  wire         queue_dataOut_7_decodeResult_red = _queue_fifo_7_data_out[102];
  wire         queue_dataOut_7_decodeResult_widenReduce = _queue_fifo_7_data_out[103];
  wire         queue_dataOut_7_decodeResult_targetRd = _queue_fifo_7_data_out[104];
  wire         queue_dataOut_7_decodeResult_slid = _queue_fifo_7_data_out[105];
  wire         queue_dataOut_7_decodeResult_gather = _queue_fifo_7_data_out[106];
  wire         queue_dataOut_7_decodeResult_gather16 = _queue_fifo_7_data_out[107];
  wire         queue_dataOut_7_decodeResult_compress = _queue_fifo_7_data_out[108];
  wire         queue_dataOut_7_decodeResult_unOrderWrite = _queue_fifo_7_data_out[109];
  wire         queue_dataOut_7_decodeResult_extend = _queue_fifo_7_data_out[110];
  wire         queue_dataOut_7_decodeResult_mv = _queue_fifo_7_data_out[111];
  wire         queue_dataOut_7_decodeResult_iota = _queue_fifo_7_data_out[112];
  wire [3:0]   queue_dataOut_7_decodeResult_uop = _queue_fifo_7_data_out[116:113];
  wire         queue_dataOut_7_decodeResult_maskLogic = _queue_fifo_7_data_out[117];
  wire         queue_dataOut_7_decodeResult_maskDestination = _queue_fifo_7_data_out[118];
  wire         queue_dataOut_7_decodeResult_maskSource = _queue_fifo_7_data_out[119];
  wire         queue_dataOut_7_decodeResult_readOnly = _queue_fifo_7_data_out[120];
  wire         queue_dataOut_7_decodeResult_vwmacc = _queue_fifo_7_data_out[121];
  wire         queue_dataOut_7_decodeResult_saturate = _queue_fifo_7_data_out[122];
  wire         queue_dataOut_7_decodeResult_special = _queue_fifo_7_data_out[123];
  wire         queue_dataOut_7_decodeResult_maskUnit = _queue_fifo_7_data_out[124];
  wire         queue_dataOut_7_decodeResult_crossWrite = _queue_fifo_7_data_out[125];
  wire         queue_dataOut_7_decodeResult_crossRead = _queue_fifo_7_data_out[126];
  wire         queue_dataOut_7_decodeResult_sWrite = _queue_fifo_7_data_out[127];
  wire         queue_dataOut_7_decodeResult_vtype = _queue_fifo_7_data_out[128];
  wire         queue_dataOut_7_decodeResult_sReadVD = _queue_fifo_7_data_out[129];
  wire         queue_dataOut_7_decodeResult_scheduler = _queue_fifo_7_data_out[130];
  wire         queue_dataOut_7_decodeResult_dontNeedExecuteInLane = _queue_fifo_7_data_out[131];
  wire         queue_dataOut_7_decodeResult_reverse = _queue_fifo_7_data_out[132];
  wire         queue_dataOut_7_decodeResult_average = _queue_fifo_7_data_out[133];
  wire         queue_dataOut_7_decodeResult_ffo = _queue_fifo_7_data_out[134];
  wire         queue_dataOut_7_decodeResult_popCount = _queue_fifo_7_data_out[135];
  wire [4:0]   queue_dataOut_7_decodeResult_topUop = _queue_fifo_7_data_out[140:136];
  wire         queue_dataOut_7_decodeResult_specialSlot = _queue_fifo_7_data_out[141];
  wire         queue_dataOut_7_decodeResult_float = _queue_fifo_7_data_out[142];
  wire [1:0]   queue_dataOut_7_decodeResult_fpExecutionType = _queue_fifo_7_data_out[144:143];
  wire         queue_dataOut_7_decodeResult_floatMul = _queue_fifo_7_data_out[145];
  wire         queue_dataOut_7_decodeResult_orderReduce = _queue_fifo_7_data_out[146];
  wire [2:0]   queue_dataOut_7_instructionIndex = _queue_fifo_7_data_out[149:147];
  wire         queue_7_enq_ready = ~_queue_fifo_7_full;
  wire         queue_7_enq_valid;
  assign queue_7_deq_valid = ~_queue_fifo_7_empty | queue_7_enq_valid;
  assign queue_7_deq_bits_instructionIndex = _queue_fifo_7_empty ? queue_7_enq_bits_instructionIndex : queue_dataOut_7_instructionIndex;
  assign queue_7_deq_bits_decodeResult_orderReduce = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_orderReduce : queue_dataOut_7_decodeResult_orderReduce;
  assign queue_7_deq_bits_decodeResult_floatMul = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_floatMul : queue_dataOut_7_decodeResult_floatMul;
  assign queue_7_deq_bits_decodeResult_fpExecutionType = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_fpExecutionType : queue_dataOut_7_decodeResult_fpExecutionType;
  assign queue_7_deq_bits_decodeResult_float = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_float : queue_dataOut_7_decodeResult_float;
  assign queue_7_deq_bits_decodeResult_specialSlot = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_specialSlot : queue_dataOut_7_decodeResult_specialSlot;
  assign queue_7_deq_bits_decodeResult_topUop = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_topUop : queue_dataOut_7_decodeResult_topUop;
  assign queue_7_deq_bits_decodeResult_popCount = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_popCount : queue_dataOut_7_decodeResult_popCount;
  assign queue_7_deq_bits_decodeResult_ffo = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_ffo : queue_dataOut_7_decodeResult_ffo;
  assign queue_7_deq_bits_decodeResult_average = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_average : queue_dataOut_7_decodeResult_average;
  assign queue_7_deq_bits_decodeResult_reverse = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_reverse : queue_dataOut_7_decodeResult_reverse;
  assign queue_7_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_7_decodeResult_dontNeedExecuteInLane;
  assign queue_7_deq_bits_decodeResult_scheduler = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_scheduler : queue_dataOut_7_decodeResult_scheduler;
  assign queue_7_deq_bits_decodeResult_sReadVD = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_sReadVD : queue_dataOut_7_decodeResult_sReadVD;
  assign queue_7_deq_bits_decodeResult_vtype = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_vtype : queue_dataOut_7_decodeResult_vtype;
  assign queue_7_deq_bits_decodeResult_sWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_sWrite : queue_dataOut_7_decodeResult_sWrite;
  assign queue_7_deq_bits_decodeResult_crossRead = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_crossRead : queue_dataOut_7_decodeResult_crossRead;
  assign queue_7_deq_bits_decodeResult_crossWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_crossWrite : queue_dataOut_7_decodeResult_crossWrite;
  assign queue_7_deq_bits_decodeResult_maskUnit = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskUnit : queue_dataOut_7_decodeResult_maskUnit;
  assign queue_7_deq_bits_decodeResult_special = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_special : queue_dataOut_7_decodeResult_special;
  assign queue_7_deq_bits_decodeResult_saturate = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_saturate : queue_dataOut_7_decodeResult_saturate;
  assign queue_7_deq_bits_decodeResult_vwmacc = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_vwmacc : queue_dataOut_7_decodeResult_vwmacc;
  assign queue_7_deq_bits_decodeResult_readOnly = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_readOnly : queue_dataOut_7_decodeResult_readOnly;
  assign queue_7_deq_bits_decodeResult_maskSource = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskSource : queue_dataOut_7_decodeResult_maskSource;
  assign queue_7_deq_bits_decodeResult_maskDestination = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskDestination : queue_dataOut_7_decodeResult_maskDestination;
  assign queue_7_deq_bits_decodeResult_maskLogic = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskLogic : queue_dataOut_7_decodeResult_maskLogic;
  assign queue_7_deq_bits_decodeResult_uop = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_uop : queue_dataOut_7_decodeResult_uop;
  assign queue_7_deq_bits_decodeResult_iota = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_iota : queue_dataOut_7_decodeResult_iota;
  assign queue_7_deq_bits_decodeResult_mv = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_mv : queue_dataOut_7_decodeResult_mv;
  assign queue_7_deq_bits_decodeResult_extend = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_extend : queue_dataOut_7_decodeResult_extend;
  assign queue_7_deq_bits_decodeResult_unOrderWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unOrderWrite : queue_dataOut_7_decodeResult_unOrderWrite;
  assign queue_7_deq_bits_decodeResult_compress = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_compress : queue_dataOut_7_decodeResult_compress;
  assign queue_7_deq_bits_decodeResult_gather16 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_gather16 : queue_dataOut_7_decodeResult_gather16;
  assign queue_7_deq_bits_decodeResult_gather = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_gather : queue_dataOut_7_decodeResult_gather;
  assign queue_7_deq_bits_decodeResult_slid = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_slid : queue_dataOut_7_decodeResult_slid;
  assign queue_7_deq_bits_decodeResult_targetRd = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_targetRd : queue_dataOut_7_decodeResult_targetRd;
  assign queue_7_deq_bits_decodeResult_widenReduce = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_widenReduce : queue_dataOut_7_decodeResult_widenReduce;
  assign queue_7_deq_bits_decodeResult_red = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_red : queue_dataOut_7_decodeResult_red;
  assign queue_7_deq_bits_decodeResult_nr = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_nr : queue_dataOut_7_decodeResult_nr;
  assign queue_7_deq_bits_decodeResult_itype = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_itype : queue_dataOut_7_decodeResult_itype;
  assign queue_7_deq_bits_decodeResult_unsigned1 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unsigned1 : queue_dataOut_7_decodeResult_unsigned1;
  assign queue_7_deq_bits_decodeResult_unsigned0 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unsigned0 : queue_dataOut_7_decodeResult_unsigned0;
  assign queue_7_deq_bits_decodeResult_other = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_other : queue_dataOut_7_decodeResult_other;
  assign queue_7_deq_bits_decodeResult_multiCycle = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_multiCycle : queue_dataOut_7_decodeResult_multiCycle;
  assign queue_7_deq_bits_decodeResult_divider = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_divider : queue_dataOut_7_decodeResult_divider;
  assign queue_7_deq_bits_decodeResult_multiplier = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_multiplier : queue_dataOut_7_decodeResult_multiplier;
  assign queue_7_deq_bits_decodeResult_shift = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_shift : queue_dataOut_7_decodeResult_shift;
  assign queue_7_deq_bits_decodeResult_adder = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_adder : queue_dataOut_7_decodeResult_adder;
  assign queue_7_deq_bits_decodeResult_logic = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_logic : queue_dataOut_7_decodeResult_logic;
  assign queue_7_deq_bits_loadStore = _queue_fifo_7_empty ? queue_7_enq_bits_loadStore : queue_dataOut_7_loadStore;
  assign queue_7_deq_bits_issueInst = _queue_fifo_7_empty ? queue_7_enq_bits_issueInst : queue_dataOut_7_issueInst;
  assign queue_7_deq_bits_store = _queue_fifo_7_empty ? queue_7_enq_bits_store : queue_dataOut_7_store;
  assign queue_7_deq_bits_special = _queue_fifo_7_empty ? queue_7_enq_bits_special : queue_dataOut_7_special;
  assign queue_7_deq_bits_lsWholeReg = _queue_fifo_7_empty ? queue_7_enq_bits_lsWholeReg : queue_dataOut_7_lsWholeReg;
  assign queue_7_deq_bits_vs1 = _queue_fifo_7_empty ? queue_7_enq_bits_vs1 : queue_dataOut_7_vs1;
  assign queue_7_deq_bits_vs2 = _queue_fifo_7_empty ? queue_7_enq_bits_vs2 : queue_dataOut_7_vs2;
  assign queue_7_deq_bits_vd = _queue_fifo_7_empty ? queue_7_enq_bits_vd : queue_dataOut_7_vd;
  assign queue_7_deq_bits_loadStoreEEW = _queue_fifo_7_empty ? queue_7_enq_bits_loadStoreEEW : queue_dataOut_7_loadStoreEEW;
  assign queue_7_deq_bits_mask = _queue_fifo_7_empty ? queue_7_enq_bits_mask : queue_dataOut_7_mask;
  assign queue_7_deq_bits_segment = _queue_fifo_7_empty ? queue_7_enq_bits_segment : queue_dataOut_7_segment;
  assign queue_7_deq_bits_readFromScalar = _queue_fifo_7_empty ? queue_7_enq_bits_readFromScalar : queue_dataOut_7_readFromScalar;
  assign queue_7_deq_bits_csrInterface_vl = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vl : queue_dataOut_7_csrInterface_vl;
  assign queue_7_deq_bits_csrInterface_vStart = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vStart : queue_dataOut_7_csrInterface_vStart;
  assign queue_7_deq_bits_csrInterface_vlmul = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vlmul : queue_dataOut_7_csrInterface_vlmul;
  assign queue_7_deq_bits_csrInterface_vSew = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vSew : queue_dataOut_7_csrInterface_vSew;
  assign queue_7_deq_bits_csrInterface_vxrm = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vxrm : queue_dataOut_7_csrInterface_vxrm;
  assign queue_7_deq_bits_csrInterface_vta = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vta : queue_dataOut_7_csrInterface_vta;
  assign queue_7_deq_bits_csrInterface_vma = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vma : queue_dataOut_7_csrInterface_vma;
  wire         laneVec_7_laneRequest_bits_issueInst = laneRequestSinkWire_7_ready & laneRequestSinkWire_7_valid;
  reg          releasePipe_pipe_v_7;
  wire         releasePipe_pipe_out_7_valid = releasePipe_pipe_v_7;
  wire         laneRequestSourceWire_7_ready;
  wire         validSource_7_valid = laneRequestSourceWire_7_ready & laneRequestSourceWire_7_valid;
  reg  [2:0]   tokenCheck_counter_7;
  wire [2:0]   tokenCheck_counterChange_7 = validSource_7_valid ? 3'h1 : 3'h7;
  assign tokenCheck_7 = ~(tokenCheck_counter_7[2]);
  assign laneRequestSourceWire_7_ready = tokenCheck_7;
  assign queue_7_enq_valid = validSink_7_valid;
  assign queue_7_enq_bits_instructionIndex = validSink_7_bits_instructionIndex;
  assign queue_7_enq_bits_decodeResult_orderReduce = validSink_7_bits_decodeResult_orderReduce;
  assign queue_7_enq_bits_decodeResult_floatMul = validSink_7_bits_decodeResult_floatMul;
  assign queue_7_enq_bits_decodeResult_fpExecutionType = validSink_7_bits_decodeResult_fpExecutionType;
  assign queue_7_enq_bits_decodeResult_float = validSink_7_bits_decodeResult_float;
  assign queue_7_enq_bits_decodeResult_specialSlot = validSink_7_bits_decodeResult_specialSlot;
  assign queue_7_enq_bits_decodeResult_topUop = validSink_7_bits_decodeResult_topUop;
  assign queue_7_enq_bits_decodeResult_popCount = validSink_7_bits_decodeResult_popCount;
  assign queue_7_enq_bits_decodeResult_ffo = validSink_7_bits_decodeResult_ffo;
  assign queue_7_enq_bits_decodeResult_average = validSink_7_bits_decodeResult_average;
  assign queue_7_enq_bits_decodeResult_reverse = validSink_7_bits_decodeResult_reverse;
  assign queue_7_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_7_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_7_enq_bits_decodeResult_scheduler = validSink_7_bits_decodeResult_scheduler;
  assign queue_7_enq_bits_decodeResult_sReadVD = validSink_7_bits_decodeResult_sReadVD;
  assign queue_7_enq_bits_decodeResult_vtype = validSink_7_bits_decodeResult_vtype;
  assign queue_7_enq_bits_decodeResult_sWrite = validSink_7_bits_decodeResult_sWrite;
  assign queue_7_enq_bits_decodeResult_crossRead = validSink_7_bits_decodeResult_crossRead;
  assign queue_7_enq_bits_decodeResult_crossWrite = validSink_7_bits_decodeResult_crossWrite;
  assign queue_7_enq_bits_decodeResult_maskUnit = validSink_7_bits_decodeResult_maskUnit;
  assign queue_7_enq_bits_decodeResult_special = validSink_7_bits_decodeResult_special;
  assign queue_7_enq_bits_decodeResult_saturate = validSink_7_bits_decodeResult_saturate;
  assign queue_7_enq_bits_decodeResult_vwmacc = validSink_7_bits_decodeResult_vwmacc;
  assign queue_7_enq_bits_decodeResult_readOnly = validSink_7_bits_decodeResult_readOnly;
  assign queue_7_enq_bits_decodeResult_maskSource = validSink_7_bits_decodeResult_maskSource;
  assign queue_7_enq_bits_decodeResult_maskDestination = validSink_7_bits_decodeResult_maskDestination;
  assign queue_7_enq_bits_decodeResult_maskLogic = validSink_7_bits_decodeResult_maskLogic;
  assign queue_7_enq_bits_decodeResult_uop = validSink_7_bits_decodeResult_uop;
  assign queue_7_enq_bits_decodeResult_iota = validSink_7_bits_decodeResult_iota;
  assign queue_7_enq_bits_decodeResult_mv = validSink_7_bits_decodeResult_mv;
  assign queue_7_enq_bits_decodeResult_extend = validSink_7_bits_decodeResult_extend;
  assign queue_7_enq_bits_decodeResult_unOrderWrite = validSink_7_bits_decodeResult_unOrderWrite;
  assign queue_7_enq_bits_decodeResult_compress = validSink_7_bits_decodeResult_compress;
  assign queue_7_enq_bits_decodeResult_gather16 = validSink_7_bits_decodeResult_gather16;
  assign queue_7_enq_bits_decodeResult_gather = validSink_7_bits_decodeResult_gather;
  assign queue_7_enq_bits_decodeResult_slid = validSink_7_bits_decodeResult_slid;
  assign queue_7_enq_bits_decodeResult_targetRd = validSink_7_bits_decodeResult_targetRd;
  assign queue_7_enq_bits_decodeResult_widenReduce = validSink_7_bits_decodeResult_widenReduce;
  assign queue_7_enq_bits_decodeResult_red = validSink_7_bits_decodeResult_red;
  assign queue_7_enq_bits_decodeResult_nr = validSink_7_bits_decodeResult_nr;
  assign queue_7_enq_bits_decodeResult_itype = validSink_7_bits_decodeResult_itype;
  assign queue_7_enq_bits_decodeResult_unsigned1 = validSink_7_bits_decodeResult_unsigned1;
  assign queue_7_enq_bits_decodeResult_unsigned0 = validSink_7_bits_decodeResult_unsigned0;
  assign queue_7_enq_bits_decodeResult_other = validSink_7_bits_decodeResult_other;
  assign queue_7_enq_bits_decodeResult_multiCycle = validSink_7_bits_decodeResult_multiCycle;
  assign queue_7_enq_bits_decodeResult_divider = validSink_7_bits_decodeResult_divider;
  assign queue_7_enq_bits_decodeResult_multiplier = validSink_7_bits_decodeResult_multiplier;
  assign queue_7_enq_bits_decodeResult_shift = validSink_7_bits_decodeResult_shift;
  assign queue_7_enq_bits_decodeResult_adder = validSink_7_bits_decodeResult_adder;
  assign queue_7_enq_bits_decodeResult_logic = validSink_7_bits_decodeResult_logic;
  assign queue_7_enq_bits_loadStore = validSink_7_bits_loadStore;
  assign queue_7_enq_bits_issueInst = validSink_7_bits_issueInst;
  assign queue_7_enq_bits_store = validSink_7_bits_store;
  assign queue_7_enq_bits_special = validSink_7_bits_special;
  assign queue_7_enq_bits_lsWholeReg = validSink_7_bits_lsWholeReg;
  assign queue_7_enq_bits_vs1 = validSink_7_bits_vs1;
  assign queue_7_enq_bits_vs2 = validSink_7_bits_vs2;
  assign queue_7_enq_bits_vd = validSink_7_bits_vd;
  assign queue_7_enq_bits_loadStoreEEW = validSink_7_bits_loadStoreEEW;
  assign queue_7_enq_bits_mask = validSink_7_bits_mask;
  assign queue_7_enq_bits_segment = validSink_7_bits_segment;
  assign queue_7_enq_bits_readFromScalar = validSink_7_bits_readFromScalar;
  assign queue_7_enq_bits_csrInterface_vl = validSink_7_bits_csrInterface_vl;
  assign queue_7_enq_bits_csrInterface_vStart = validSink_7_bits_csrInterface_vStart;
  assign queue_7_enq_bits_csrInterface_vlmul = validSink_7_bits_csrInterface_vlmul;
  assign queue_7_enq_bits_csrInterface_vSew = validSink_7_bits_csrInterface_vSew;
  assign queue_7_enq_bits_csrInterface_vxrm = validSink_7_bits_csrInterface_vxrm;
  assign queue_7_enq_bits_csrInterface_vta = validSink_7_bits_csrInterface_vta;
  assign queue_7_enq_bits_csrInterface_vma = validSink_7_bits_csrInterface_vma;
  reg          shifterReg_7_0_valid;
  assign validSink_7_valid = shifterReg_7_0_valid;
  reg  [2:0]   shifterReg_7_0_bits_instructionIndex;
  assign validSink_7_bits_instructionIndex = shifterReg_7_0_bits_instructionIndex;
  reg          shifterReg_7_0_bits_decodeResult_orderReduce;
  assign validSink_7_bits_decodeResult_orderReduce = shifterReg_7_0_bits_decodeResult_orderReduce;
  reg          shifterReg_7_0_bits_decodeResult_floatMul;
  assign validSink_7_bits_decodeResult_floatMul = shifterReg_7_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_7_0_bits_decodeResult_fpExecutionType;
  assign validSink_7_bits_decodeResult_fpExecutionType = shifterReg_7_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_7_0_bits_decodeResult_float;
  assign validSink_7_bits_decodeResult_float = shifterReg_7_0_bits_decodeResult_float;
  reg          shifterReg_7_0_bits_decodeResult_specialSlot;
  assign validSink_7_bits_decodeResult_specialSlot = shifterReg_7_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_7_0_bits_decodeResult_topUop;
  assign validSink_7_bits_decodeResult_topUop = shifterReg_7_0_bits_decodeResult_topUop;
  reg          shifterReg_7_0_bits_decodeResult_popCount;
  assign validSink_7_bits_decodeResult_popCount = shifterReg_7_0_bits_decodeResult_popCount;
  reg          shifterReg_7_0_bits_decodeResult_ffo;
  assign validSink_7_bits_decodeResult_ffo = shifterReg_7_0_bits_decodeResult_ffo;
  reg          shifterReg_7_0_bits_decodeResult_average;
  assign validSink_7_bits_decodeResult_average = shifterReg_7_0_bits_decodeResult_average;
  reg          shifterReg_7_0_bits_decodeResult_reverse;
  assign validSink_7_bits_decodeResult_reverse = shifterReg_7_0_bits_decodeResult_reverse;
  reg          shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_7_bits_decodeResult_dontNeedExecuteInLane = shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_7_0_bits_decodeResult_scheduler;
  assign validSink_7_bits_decodeResult_scheduler = shifterReg_7_0_bits_decodeResult_scheduler;
  reg          shifterReg_7_0_bits_decodeResult_sReadVD;
  assign validSink_7_bits_decodeResult_sReadVD = shifterReg_7_0_bits_decodeResult_sReadVD;
  reg          shifterReg_7_0_bits_decodeResult_vtype;
  assign validSink_7_bits_decodeResult_vtype = shifterReg_7_0_bits_decodeResult_vtype;
  reg          shifterReg_7_0_bits_decodeResult_sWrite;
  assign validSink_7_bits_decodeResult_sWrite = shifterReg_7_0_bits_decodeResult_sWrite;
  reg          shifterReg_7_0_bits_decodeResult_crossRead;
  assign validSink_7_bits_decodeResult_crossRead = shifterReg_7_0_bits_decodeResult_crossRead;
  reg          shifterReg_7_0_bits_decodeResult_crossWrite;
  assign validSink_7_bits_decodeResult_crossWrite = shifterReg_7_0_bits_decodeResult_crossWrite;
  reg          shifterReg_7_0_bits_decodeResult_maskUnit;
  assign validSink_7_bits_decodeResult_maskUnit = shifterReg_7_0_bits_decodeResult_maskUnit;
  reg          shifterReg_7_0_bits_decodeResult_special;
  assign validSink_7_bits_decodeResult_special = shifterReg_7_0_bits_decodeResult_special;
  reg          shifterReg_7_0_bits_decodeResult_saturate;
  assign validSink_7_bits_decodeResult_saturate = shifterReg_7_0_bits_decodeResult_saturate;
  reg          shifterReg_7_0_bits_decodeResult_vwmacc;
  assign validSink_7_bits_decodeResult_vwmacc = shifterReg_7_0_bits_decodeResult_vwmacc;
  reg          shifterReg_7_0_bits_decodeResult_readOnly;
  assign validSink_7_bits_decodeResult_readOnly = shifterReg_7_0_bits_decodeResult_readOnly;
  reg          shifterReg_7_0_bits_decodeResult_maskSource;
  assign validSink_7_bits_decodeResult_maskSource = shifterReg_7_0_bits_decodeResult_maskSource;
  reg          shifterReg_7_0_bits_decodeResult_maskDestination;
  assign validSink_7_bits_decodeResult_maskDestination = shifterReg_7_0_bits_decodeResult_maskDestination;
  reg          shifterReg_7_0_bits_decodeResult_maskLogic;
  assign validSink_7_bits_decodeResult_maskLogic = shifterReg_7_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_7_0_bits_decodeResult_uop;
  assign validSink_7_bits_decodeResult_uop = shifterReg_7_0_bits_decodeResult_uop;
  reg          shifterReg_7_0_bits_decodeResult_iota;
  assign validSink_7_bits_decodeResult_iota = shifterReg_7_0_bits_decodeResult_iota;
  reg          shifterReg_7_0_bits_decodeResult_mv;
  assign validSink_7_bits_decodeResult_mv = shifterReg_7_0_bits_decodeResult_mv;
  reg          shifterReg_7_0_bits_decodeResult_extend;
  assign validSink_7_bits_decodeResult_extend = shifterReg_7_0_bits_decodeResult_extend;
  reg          shifterReg_7_0_bits_decodeResult_unOrderWrite;
  assign validSink_7_bits_decodeResult_unOrderWrite = shifterReg_7_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_7_0_bits_decodeResult_compress;
  assign validSink_7_bits_decodeResult_compress = shifterReg_7_0_bits_decodeResult_compress;
  reg          shifterReg_7_0_bits_decodeResult_gather16;
  assign validSink_7_bits_decodeResult_gather16 = shifterReg_7_0_bits_decodeResult_gather16;
  reg          shifterReg_7_0_bits_decodeResult_gather;
  assign validSink_7_bits_decodeResult_gather = shifterReg_7_0_bits_decodeResult_gather;
  reg          shifterReg_7_0_bits_decodeResult_slid;
  assign validSink_7_bits_decodeResult_slid = shifterReg_7_0_bits_decodeResult_slid;
  reg          shifterReg_7_0_bits_decodeResult_targetRd;
  assign validSink_7_bits_decodeResult_targetRd = shifterReg_7_0_bits_decodeResult_targetRd;
  reg          shifterReg_7_0_bits_decodeResult_widenReduce;
  assign validSink_7_bits_decodeResult_widenReduce = shifterReg_7_0_bits_decodeResult_widenReduce;
  reg          shifterReg_7_0_bits_decodeResult_red;
  assign validSink_7_bits_decodeResult_red = shifterReg_7_0_bits_decodeResult_red;
  reg          shifterReg_7_0_bits_decodeResult_nr;
  assign validSink_7_bits_decodeResult_nr = shifterReg_7_0_bits_decodeResult_nr;
  reg          shifterReg_7_0_bits_decodeResult_itype;
  assign validSink_7_bits_decodeResult_itype = shifterReg_7_0_bits_decodeResult_itype;
  reg          shifterReg_7_0_bits_decodeResult_unsigned1;
  assign validSink_7_bits_decodeResult_unsigned1 = shifterReg_7_0_bits_decodeResult_unsigned1;
  reg          shifterReg_7_0_bits_decodeResult_unsigned0;
  assign validSink_7_bits_decodeResult_unsigned0 = shifterReg_7_0_bits_decodeResult_unsigned0;
  reg          shifterReg_7_0_bits_decodeResult_other;
  assign validSink_7_bits_decodeResult_other = shifterReg_7_0_bits_decodeResult_other;
  reg          shifterReg_7_0_bits_decodeResult_multiCycle;
  assign validSink_7_bits_decodeResult_multiCycle = shifterReg_7_0_bits_decodeResult_multiCycle;
  reg          shifterReg_7_0_bits_decodeResult_divider;
  assign validSink_7_bits_decodeResult_divider = shifterReg_7_0_bits_decodeResult_divider;
  reg          shifterReg_7_0_bits_decodeResult_multiplier;
  assign validSink_7_bits_decodeResult_multiplier = shifterReg_7_0_bits_decodeResult_multiplier;
  reg          shifterReg_7_0_bits_decodeResult_shift;
  assign validSink_7_bits_decodeResult_shift = shifterReg_7_0_bits_decodeResult_shift;
  reg          shifterReg_7_0_bits_decodeResult_adder;
  assign validSink_7_bits_decodeResult_adder = shifterReg_7_0_bits_decodeResult_adder;
  reg          shifterReg_7_0_bits_decodeResult_logic;
  assign validSink_7_bits_decodeResult_logic = shifterReg_7_0_bits_decodeResult_logic;
  reg          shifterReg_7_0_bits_loadStore;
  assign validSink_7_bits_loadStore = shifterReg_7_0_bits_loadStore;
  reg          shifterReg_7_0_bits_issueInst;
  assign validSink_7_bits_issueInst = shifterReg_7_0_bits_issueInst;
  reg          shifterReg_7_0_bits_store;
  assign validSink_7_bits_store = shifterReg_7_0_bits_store;
  reg          shifterReg_7_0_bits_special;
  assign validSink_7_bits_special = shifterReg_7_0_bits_special;
  reg          shifterReg_7_0_bits_lsWholeReg;
  assign validSink_7_bits_lsWholeReg = shifterReg_7_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_7_0_bits_vs1;
  assign validSink_7_bits_vs1 = shifterReg_7_0_bits_vs1;
  reg  [4:0]   shifterReg_7_0_bits_vs2;
  assign validSink_7_bits_vs2 = shifterReg_7_0_bits_vs2;
  reg  [4:0]   shifterReg_7_0_bits_vd;
  assign validSink_7_bits_vd = shifterReg_7_0_bits_vd;
  reg  [1:0]   shifterReg_7_0_bits_loadStoreEEW;
  assign validSink_7_bits_loadStoreEEW = shifterReg_7_0_bits_loadStoreEEW;
  reg          shifterReg_7_0_bits_mask;
  assign validSink_7_bits_mask = shifterReg_7_0_bits_mask;
  reg  [2:0]   shifterReg_7_0_bits_segment;
  assign validSink_7_bits_segment = shifterReg_7_0_bits_segment;
  reg  [31:0]  shifterReg_7_0_bits_readFromScalar;
  assign validSink_7_bits_readFromScalar = shifterReg_7_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_7_0_bits_csrInterface_vl;
  assign validSink_7_bits_csrInterface_vl = shifterReg_7_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_7_0_bits_csrInterface_vStart;
  assign validSink_7_bits_csrInterface_vStart = shifterReg_7_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_7_0_bits_csrInterface_vlmul;
  assign validSink_7_bits_csrInterface_vlmul = shifterReg_7_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_7_0_bits_csrInterface_vSew;
  assign validSink_7_bits_csrInterface_vSew = shifterReg_7_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_7_0_bits_csrInterface_vxrm;
  assign validSink_7_bits_csrInterface_vxrm = shifterReg_7_0_bits_csrInterface_vxrm;
  reg          shifterReg_7_0_bits_csrInterface_vta;
  assign validSink_7_bits_csrInterface_vta = shifterReg_7_0_bits_csrInterface_vta;
  reg          shifterReg_7_0_bits_csrInterface_vma;
  assign validSink_7_bits_csrInterface_vma = shifterReg_7_0_bits_csrInterface_vma;
  wire         shifterValid_7 = shifterReg_7_0_valid | validSource_7_valid;
  wire         validSink_8_valid;
  wire [2:0]   validSink_8_bits_instructionIndex;
  wire         validSink_8_bits_decodeResult_orderReduce;
  wire         validSink_8_bits_decodeResult_floatMul;
  wire [1:0]   validSink_8_bits_decodeResult_fpExecutionType;
  wire         validSink_8_bits_decodeResult_float;
  wire         validSink_8_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_8_bits_decodeResult_topUop;
  wire         validSink_8_bits_decodeResult_popCount;
  wire         validSink_8_bits_decodeResult_ffo;
  wire         validSink_8_bits_decodeResult_average;
  wire         validSink_8_bits_decodeResult_reverse;
  wire         validSink_8_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_8_bits_decodeResult_scheduler;
  wire         validSink_8_bits_decodeResult_sReadVD;
  wire         validSink_8_bits_decodeResult_vtype;
  wire         validSink_8_bits_decodeResult_sWrite;
  wire         validSink_8_bits_decodeResult_crossRead;
  wire         validSink_8_bits_decodeResult_crossWrite;
  wire         validSink_8_bits_decodeResult_maskUnit;
  wire         validSink_8_bits_decodeResult_special;
  wire         validSink_8_bits_decodeResult_saturate;
  wire         validSink_8_bits_decodeResult_vwmacc;
  wire         validSink_8_bits_decodeResult_readOnly;
  wire         validSink_8_bits_decodeResult_maskSource;
  wire         validSink_8_bits_decodeResult_maskDestination;
  wire         validSink_8_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_8_bits_decodeResult_uop;
  wire         validSink_8_bits_decodeResult_iota;
  wire         validSink_8_bits_decodeResult_mv;
  wire         validSink_8_bits_decodeResult_extend;
  wire         validSink_8_bits_decodeResult_unOrderWrite;
  wire         validSink_8_bits_decodeResult_compress;
  wire         validSink_8_bits_decodeResult_gather16;
  wire         validSink_8_bits_decodeResult_gather;
  wire         validSink_8_bits_decodeResult_slid;
  wire         validSink_8_bits_decodeResult_targetRd;
  wire         validSink_8_bits_decodeResult_widenReduce;
  wire         validSink_8_bits_decodeResult_red;
  wire         validSink_8_bits_decodeResult_nr;
  wire         validSink_8_bits_decodeResult_itype;
  wire         validSink_8_bits_decodeResult_unsigned1;
  wire         validSink_8_bits_decodeResult_unsigned0;
  wire         validSink_8_bits_decodeResult_other;
  wire         validSink_8_bits_decodeResult_multiCycle;
  wire         validSink_8_bits_decodeResult_divider;
  wire         validSink_8_bits_decodeResult_multiplier;
  wire         validSink_8_bits_decodeResult_shift;
  wire         validSink_8_bits_decodeResult_adder;
  wire         validSink_8_bits_decodeResult_logic;
  wire         validSink_8_bits_loadStore;
  wire         validSink_8_bits_issueInst;
  wire         validSink_8_bits_store;
  wire         validSink_8_bits_special;
  wire         validSink_8_bits_lsWholeReg;
  wire [4:0]   validSink_8_bits_vs1;
  wire [4:0]   validSink_8_bits_vs2;
  wire [4:0]   validSink_8_bits_vd;
  wire [1:0]   validSink_8_bits_loadStoreEEW;
  wire         validSink_8_bits_mask;
  wire [2:0]   validSink_8_bits_segment;
  wire [31:0]  validSink_8_bits_readFromScalar;
  wire [11:0]  validSink_8_bits_csrInterface_vl;
  wire [11:0]  validSink_8_bits_csrInterface_vStart;
  wire [2:0]   validSink_8_bits_csrInterface_vlmul;
  wire [1:0]   validSink_8_bits_csrInterface_vSew;
  wire [1:0]   validSink_8_bits_csrInterface_vxrm;
  wire         validSink_8_bits_csrInterface_vta;
  wire         validSink_8_bits_csrInterface_vma;
  wire         laneRequestSinkWire_8_valid = queue_8_deq_valid;
  wire [2:0]   laneRequestSinkWire_8_bits_instructionIndex = queue_8_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_8_bits_decodeResult_orderReduce = queue_8_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_8_bits_decodeResult_floatMul = queue_8_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_8_bits_decodeResult_fpExecutionType = queue_8_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_8_bits_decodeResult_float = queue_8_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_8_bits_decodeResult_specialSlot = queue_8_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_8_bits_decodeResult_topUop = queue_8_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_8_bits_decodeResult_popCount = queue_8_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_8_bits_decodeResult_ffo = queue_8_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_8_bits_decodeResult_average = queue_8_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_8_bits_decodeResult_reverse = queue_8_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_8_bits_decodeResult_dontNeedExecuteInLane = queue_8_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_8_bits_decodeResult_scheduler = queue_8_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_8_bits_decodeResult_sReadVD = queue_8_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_8_bits_decodeResult_vtype = queue_8_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_8_bits_decodeResult_sWrite = queue_8_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_8_bits_decodeResult_crossRead = queue_8_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_8_bits_decodeResult_crossWrite = queue_8_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_8_bits_decodeResult_maskUnit = queue_8_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_8_bits_decodeResult_special = queue_8_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_8_bits_decodeResult_saturate = queue_8_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_8_bits_decodeResult_vwmacc = queue_8_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_8_bits_decodeResult_readOnly = queue_8_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_8_bits_decodeResult_maskSource = queue_8_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_8_bits_decodeResult_maskDestination = queue_8_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_8_bits_decodeResult_maskLogic = queue_8_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_8_bits_decodeResult_uop = queue_8_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_8_bits_decodeResult_iota = queue_8_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_8_bits_decodeResult_mv = queue_8_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_8_bits_decodeResult_extend = queue_8_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_8_bits_decodeResult_unOrderWrite = queue_8_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_8_bits_decodeResult_compress = queue_8_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_8_bits_decodeResult_gather16 = queue_8_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_8_bits_decodeResult_gather = queue_8_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_8_bits_decodeResult_slid = queue_8_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_8_bits_decodeResult_targetRd = queue_8_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_8_bits_decodeResult_widenReduce = queue_8_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_8_bits_decodeResult_red = queue_8_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_8_bits_decodeResult_nr = queue_8_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_8_bits_decodeResult_itype = queue_8_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_8_bits_decodeResult_unsigned1 = queue_8_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_8_bits_decodeResult_unsigned0 = queue_8_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_8_bits_decodeResult_other = queue_8_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_8_bits_decodeResult_multiCycle = queue_8_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_8_bits_decodeResult_divider = queue_8_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_8_bits_decodeResult_multiplier = queue_8_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_8_bits_decodeResult_shift = queue_8_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_8_bits_decodeResult_adder = queue_8_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_8_bits_decodeResult_logic = queue_8_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_8_bits_loadStore = queue_8_deq_bits_loadStore;
  wire         laneRequestSinkWire_8_bits_issueInst = queue_8_deq_bits_issueInst;
  wire         laneRequestSinkWire_8_bits_store = queue_8_deq_bits_store;
  wire         laneRequestSinkWire_8_bits_special = queue_8_deq_bits_special;
  wire         laneRequestSinkWire_8_bits_lsWholeReg = queue_8_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_8_bits_vs1 = queue_8_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_8_bits_vs2 = queue_8_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_8_bits_vd = queue_8_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_8_bits_loadStoreEEW = queue_8_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_8_bits_mask = queue_8_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_8_bits_segment = queue_8_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_8_bits_readFromScalar = queue_8_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_8_bits_csrInterface_vl = queue_8_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_8_bits_csrInterface_vStart = queue_8_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_8_bits_csrInterface_vlmul = queue_8_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_8_bits_csrInterface_vSew = queue_8_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_8_bits_csrInterface_vxrm = queue_8_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_8_bits_csrInterface_vta = queue_8_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_8_bits_csrInterface_vma = queue_8_deq_bits_csrInterface_vma;
  wire [1:0]   queue_8_enq_bits_csrInterface_vxrm;
  wire         queue_8_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_24 = {queue_8_enq_bits_csrInterface_vxrm, queue_8_enq_bits_csrInterface_vta};
  wire         queue_8_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_24 = {queue_dataIn_lo_hi_24, queue_8_enq_bits_csrInterface_vma};
  wire [2:0]   queue_8_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_8_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_24 = {queue_8_enq_bits_csrInterface_vlmul, queue_8_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_8_enq_bits_csrInterface_vl;
  wire [11:0]  queue_8_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_24 = {queue_8_enq_bits_csrInterface_vl, queue_8_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_24 = {queue_dataIn_hi_hi_24, queue_dataIn_hi_lo_24};
  wire         queue_8_enq_bits_decodeResult_shift;
  wire         queue_8_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_8 = {queue_8_enq_bits_decodeResult_shift, queue_8_enq_bits_decodeResult_adder};
  wire         queue_8_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_8 = {queue_dataIn_lo_lo_lo_lo_hi_8, queue_8_enq_bits_decodeResult_logic};
  wire         queue_8_enq_bits_decodeResult_multiCycle;
  wire         queue_8_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_8 = {queue_8_enq_bits_decodeResult_multiCycle, queue_8_enq_bits_decodeResult_divider};
  wire         queue_8_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_8 = {queue_dataIn_lo_lo_lo_hi_hi_8, queue_8_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_8 = {queue_dataIn_lo_lo_lo_hi_8, queue_dataIn_lo_lo_lo_lo_8};
  wire         queue_8_enq_bits_decodeResult_unsigned1;
  wire         queue_8_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_8 = {queue_8_enq_bits_decodeResult_unsigned1, queue_8_enq_bits_decodeResult_unsigned0};
  wire         queue_8_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_8 = {queue_dataIn_lo_lo_hi_lo_hi_8, queue_8_enq_bits_decodeResult_other};
  wire         queue_8_enq_bits_decodeResult_red;
  wire         queue_8_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_8 = {queue_8_enq_bits_decodeResult_red, queue_8_enq_bits_decodeResult_nr};
  wire         queue_8_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_8 = {queue_dataIn_lo_lo_hi_hi_hi_8, queue_8_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_16 = {queue_dataIn_lo_lo_hi_hi_8, queue_dataIn_lo_lo_hi_lo_8};
  wire [11:0]  queue_dataIn_lo_lo_16 = {queue_dataIn_lo_lo_hi_16, queue_dataIn_lo_lo_lo_8};
  wire         queue_8_enq_bits_decodeResult_slid;
  wire         queue_8_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_8 = {queue_8_enq_bits_decodeResult_slid, queue_8_enq_bits_decodeResult_targetRd};
  wire         queue_8_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_8 = {queue_dataIn_lo_hi_lo_lo_hi_8, queue_8_enq_bits_decodeResult_widenReduce};
  wire         queue_8_enq_bits_decodeResult_compress;
  wire         queue_8_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_8 = {queue_8_enq_bits_decodeResult_compress, queue_8_enq_bits_decodeResult_gather16};
  wire         queue_8_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_8 = {queue_dataIn_lo_hi_lo_hi_hi_8, queue_8_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_16 = {queue_dataIn_lo_hi_lo_hi_8, queue_dataIn_lo_hi_lo_lo_8};
  wire         queue_8_enq_bits_decodeResult_mv;
  wire         queue_8_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_8 = {queue_8_enq_bits_decodeResult_mv, queue_8_enq_bits_decodeResult_extend};
  wire         queue_8_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_8 = {queue_dataIn_lo_hi_hi_lo_hi_8, queue_8_enq_bits_decodeResult_unOrderWrite};
  wire         queue_8_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_8_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_8 = {queue_8_enq_bits_decodeResult_maskLogic, queue_8_enq_bits_decodeResult_uop};
  wire         queue_8_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_8 = {queue_dataIn_lo_hi_hi_hi_hi_8, queue_8_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_16 = {queue_dataIn_lo_hi_hi_hi_8, queue_dataIn_lo_hi_hi_lo_8};
  wire [14:0]  queue_dataIn_lo_hi_25 = {queue_dataIn_lo_hi_hi_16, queue_dataIn_lo_hi_lo_16};
  wire [26:0]  queue_dataIn_lo_25 = {queue_dataIn_lo_hi_25, queue_dataIn_lo_lo_16};
  wire         queue_8_enq_bits_decodeResult_readOnly;
  wire         queue_8_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_8 = {queue_8_enq_bits_decodeResult_readOnly, queue_8_enq_bits_decodeResult_maskSource};
  wire         queue_8_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_8 = {queue_dataIn_hi_lo_lo_lo_hi_8, queue_8_enq_bits_decodeResult_maskDestination};
  wire         queue_8_enq_bits_decodeResult_special;
  wire         queue_8_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_8 = {queue_8_enq_bits_decodeResult_special, queue_8_enq_bits_decodeResult_saturate};
  wire         queue_8_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_8 = {queue_dataIn_hi_lo_lo_hi_hi_8, queue_8_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_16 = {queue_dataIn_hi_lo_lo_hi_8, queue_dataIn_hi_lo_lo_lo_8};
  wire         queue_8_enq_bits_decodeResult_crossRead;
  wire         queue_8_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_8 = {queue_8_enq_bits_decodeResult_crossRead, queue_8_enq_bits_decodeResult_crossWrite};
  wire         queue_8_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_8 = {queue_dataIn_hi_lo_hi_lo_hi_8, queue_8_enq_bits_decodeResult_maskUnit};
  wire         queue_8_enq_bits_decodeResult_sReadVD;
  wire         queue_8_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_8 = {queue_8_enq_bits_decodeResult_sReadVD, queue_8_enq_bits_decodeResult_vtype};
  wire         queue_8_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_8 = {queue_dataIn_hi_lo_hi_hi_hi_8, queue_8_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_16 = {queue_dataIn_hi_lo_hi_hi_8, queue_dataIn_hi_lo_hi_lo_8};
  wire [11:0]  queue_dataIn_hi_lo_25 = {queue_dataIn_hi_lo_hi_16, queue_dataIn_hi_lo_lo_16};
  wire         queue_8_enq_bits_decodeResult_reverse;
  wire         queue_8_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_8 = {queue_8_enq_bits_decodeResult_reverse, queue_8_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_8_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_8 = {queue_dataIn_hi_hi_lo_lo_hi_8, queue_8_enq_bits_decodeResult_scheduler};
  wire         queue_8_enq_bits_decodeResult_popCount;
  wire         queue_8_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_8 = {queue_8_enq_bits_decodeResult_popCount, queue_8_enq_bits_decodeResult_ffo};
  wire         queue_8_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_8 = {queue_dataIn_hi_hi_lo_hi_hi_8, queue_8_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_16 = {queue_dataIn_hi_hi_lo_hi_8, queue_dataIn_hi_hi_lo_lo_8};
  wire         queue_8_enq_bits_decodeResult_float;
  wire         queue_8_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_8 = {queue_8_enq_bits_decodeResult_float, queue_8_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_8_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_8 = {queue_dataIn_hi_hi_hi_lo_hi_8, queue_8_enq_bits_decodeResult_topUop};
  wire         queue_8_enq_bits_decodeResult_orderReduce;
  wire         queue_8_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_8 = {queue_8_enq_bits_decodeResult_orderReduce, queue_8_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_8_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_8 = {queue_dataIn_hi_hi_hi_hi_hi_8, queue_8_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_16 = {queue_dataIn_hi_hi_hi_hi_8, queue_dataIn_hi_hi_hi_lo_8};
  wire [16:0]  queue_dataIn_hi_hi_25 = {queue_dataIn_hi_hi_hi_16, queue_dataIn_hi_hi_lo_16};
  wire [28:0]  queue_dataIn_hi_25 = {queue_dataIn_hi_hi_25, queue_dataIn_hi_lo_25};
  wire [2:0]   queue_8_enq_bits_segment;
  wire [31:0]  queue_8_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_17 = {queue_8_enq_bits_segment, queue_8_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_17 = {queue_dataIn_lo_lo_hi_17, queue_dataIn_hi_24, queue_dataIn_lo_24};
  wire [1:0]   queue_8_enq_bits_loadStoreEEW;
  wire         queue_8_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_17 = {queue_8_enq_bits_loadStoreEEW, queue_8_enq_bits_mask};
  wire [4:0]   queue_8_enq_bits_vs2;
  wire [4:0]   queue_8_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_17 = {queue_8_enq_bits_vs2, queue_8_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_26 = {queue_dataIn_lo_hi_hi_17, queue_dataIn_lo_hi_lo_17};
  wire [80:0]  queue_dataIn_lo_26 = {queue_dataIn_lo_hi_26, queue_dataIn_lo_lo_17};
  wire         queue_8_enq_bits_lsWholeReg;
  wire [4:0]   queue_8_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_17 = {queue_8_enq_bits_lsWholeReg, queue_8_enq_bits_vs1};
  wire         queue_8_enq_bits_store;
  wire         queue_8_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_17 = {queue_8_enq_bits_store, queue_8_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_26 = {queue_dataIn_hi_lo_hi_17, queue_dataIn_hi_lo_lo_17};
  wire         queue_8_enq_bits_loadStore;
  wire         queue_8_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_17 = {queue_8_enq_bits_loadStore, queue_8_enq_bits_issueInst};
  wire [2:0]   queue_8_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_17 = {queue_8_enq_bits_instructionIndex, queue_dataIn_hi_25, queue_dataIn_lo_25};
  wire [60:0]  queue_dataIn_hi_hi_26 = {queue_dataIn_hi_hi_hi_17, queue_dataIn_hi_hi_lo_17};
  wire [68:0]  queue_dataIn_hi_26 = {queue_dataIn_hi_hi_26, queue_dataIn_hi_lo_26};
  wire [149:0] queue_dataIn_8 = {queue_dataIn_hi_26, queue_dataIn_lo_26};
  wire         queue_dataOut_8_csrInterface_vma = _queue_fifo_8_data_out[0];
  wire         queue_dataOut_8_csrInterface_vta = _queue_fifo_8_data_out[1];
  wire [1:0]   queue_dataOut_8_csrInterface_vxrm = _queue_fifo_8_data_out[3:2];
  wire [1:0]   queue_dataOut_8_csrInterface_vSew = _queue_fifo_8_data_out[5:4];
  wire [2:0]   queue_dataOut_8_csrInterface_vlmul = _queue_fifo_8_data_out[8:6];
  wire [11:0]  queue_dataOut_8_csrInterface_vStart = _queue_fifo_8_data_out[20:9];
  wire [11:0]  queue_dataOut_8_csrInterface_vl = _queue_fifo_8_data_out[32:21];
  wire [31:0]  queue_dataOut_8_readFromScalar = _queue_fifo_8_data_out[64:33];
  wire [2:0]   queue_dataOut_8_segment = _queue_fifo_8_data_out[67:65];
  wire         queue_dataOut_8_mask = _queue_fifo_8_data_out[68];
  wire [1:0]   queue_dataOut_8_loadStoreEEW = _queue_fifo_8_data_out[70:69];
  wire [4:0]   queue_dataOut_8_vd = _queue_fifo_8_data_out[75:71];
  wire [4:0]   queue_dataOut_8_vs2 = _queue_fifo_8_data_out[80:76];
  wire [4:0]   queue_dataOut_8_vs1 = _queue_fifo_8_data_out[85:81];
  wire         queue_dataOut_8_lsWholeReg = _queue_fifo_8_data_out[86];
  wire         queue_dataOut_8_special = _queue_fifo_8_data_out[87];
  wire         queue_dataOut_8_store = _queue_fifo_8_data_out[88];
  wire         queue_dataOut_8_issueInst = _queue_fifo_8_data_out[89];
  wire         queue_dataOut_8_loadStore = _queue_fifo_8_data_out[90];
  wire         queue_dataOut_8_decodeResult_logic = _queue_fifo_8_data_out[91];
  wire         queue_dataOut_8_decodeResult_adder = _queue_fifo_8_data_out[92];
  wire         queue_dataOut_8_decodeResult_shift = _queue_fifo_8_data_out[93];
  wire         queue_dataOut_8_decodeResult_multiplier = _queue_fifo_8_data_out[94];
  wire         queue_dataOut_8_decodeResult_divider = _queue_fifo_8_data_out[95];
  wire         queue_dataOut_8_decodeResult_multiCycle = _queue_fifo_8_data_out[96];
  wire         queue_dataOut_8_decodeResult_other = _queue_fifo_8_data_out[97];
  wire         queue_dataOut_8_decodeResult_unsigned0 = _queue_fifo_8_data_out[98];
  wire         queue_dataOut_8_decodeResult_unsigned1 = _queue_fifo_8_data_out[99];
  wire         queue_dataOut_8_decodeResult_itype = _queue_fifo_8_data_out[100];
  wire         queue_dataOut_8_decodeResult_nr = _queue_fifo_8_data_out[101];
  wire         queue_dataOut_8_decodeResult_red = _queue_fifo_8_data_out[102];
  wire         queue_dataOut_8_decodeResult_widenReduce = _queue_fifo_8_data_out[103];
  wire         queue_dataOut_8_decodeResult_targetRd = _queue_fifo_8_data_out[104];
  wire         queue_dataOut_8_decodeResult_slid = _queue_fifo_8_data_out[105];
  wire         queue_dataOut_8_decodeResult_gather = _queue_fifo_8_data_out[106];
  wire         queue_dataOut_8_decodeResult_gather16 = _queue_fifo_8_data_out[107];
  wire         queue_dataOut_8_decodeResult_compress = _queue_fifo_8_data_out[108];
  wire         queue_dataOut_8_decodeResult_unOrderWrite = _queue_fifo_8_data_out[109];
  wire         queue_dataOut_8_decodeResult_extend = _queue_fifo_8_data_out[110];
  wire         queue_dataOut_8_decodeResult_mv = _queue_fifo_8_data_out[111];
  wire         queue_dataOut_8_decodeResult_iota = _queue_fifo_8_data_out[112];
  wire [3:0]   queue_dataOut_8_decodeResult_uop = _queue_fifo_8_data_out[116:113];
  wire         queue_dataOut_8_decodeResult_maskLogic = _queue_fifo_8_data_out[117];
  wire         queue_dataOut_8_decodeResult_maskDestination = _queue_fifo_8_data_out[118];
  wire         queue_dataOut_8_decodeResult_maskSource = _queue_fifo_8_data_out[119];
  wire         queue_dataOut_8_decodeResult_readOnly = _queue_fifo_8_data_out[120];
  wire         queue_dataOut_8_decodeResult_vwmacc = _queue_fifo_8_data_out[121];
  wire         queue_dataOut_8_decodeResult_saturate = _queue_fifo_8_data_out[122];
  wire         queue_dataOut_8_decodeResult_special = _queue_fifo_8_data_out[123];
  wire         queue_dataOut_8_decodeResult_maskUnit = _queue_fifo_8_data_out[124];
  wire         queue_dataOut_8_decodeResult_crossWrite = _queue_fifo_8_data_out[125];
  wire         queue_dataOut_8_decodeResult_crossRead = _queue_fifo_8_data_out[126];
  wire         queue_dataOut_8_decodeResult_sWrite = _queue_fifo_8_data_out[127];
  wire         queue_dataOut_8_decodeResult_vtype = _queue_fifo_8_data_out[128];
  wire         queue_dataOut_8_decodeResult_sReadVD = _queue_fifo_8_data_out[129];
  wire         queue_dataOut_8_decodeResult_scheduler = _queue_fifo_8_data_out[130];
  wire         queue_dataOut_8_decodeResult_dontNeedExecuteInLane = _queue_fifo_8_data_out[131];
  wire         queue_dataOut_8_decodeResult_reverse = _queue_fifo_8_data_out[132];
  wire         queue_dataOut_8_decodeResult_average = _queue_fifo_8_data_out[133];
  wire         queue_dataOut_8_decodeResult_ffo = _queue_fifo_8_data_out[134];
  wire         queue_dataOut_8_decodeResult_popCount = _queue_fifo_8_data_out[135];
  wire [4:0]   queue_dataOut_8_decodeResult_topUop = _queue_fifo_8_data_out[140:136];
  wire         queue_dataOut_8_decodeResult_specialSlot = _queue_fifo_8_data_out[141];
  wire         queue_dataOut_8_decodeResult_float = _queue_fifo_8_data_out[142];
  wire [1:0]   queue_dataOut_8_decodeResult_fpExecutionType = _queue_fifo_8_data_out[144:143];
  wire         queue_dataOut_8_decodeResult_floatMul = _queue_fifo_8_data_out[145];
  wire         queue_dataOut_8_decodeResult_orderReduce = _queue_fifo_8_data_out[146];
  wire [2:0]   queue_dataOut_8_instructionIndex = _queue_fifo_8_data_out[149:147];
  wire         queue_8_enq_ready = ~_queue_fifo_8_full;
  wire         queue_8_enq_valid;
  assign queue_8_deq_valid = ~_queue_fifo_8_empty | queue_8_enq_valid;
  assign queue_8_deq_bits_instructionIndex = _queue_fifo_8_empty ? queue_8_enq_bits_instructionIndex : queue_dataOut_8_instructionIndex;
  assign queue_8_deq_bits_decodeResult_orderReduce = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_orderReduce : queue_dataOut_8_decodeResult_orderReduce;
  assign queue_8_deq_bits_decodeResult_floatMul = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_floatMul : queue_dataOut_8_decodeResult_floatMul;
  assign queue_8_deq_bits_decodeResult_fpExecutionType = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_fpExecutionType : queue_dataOut_8_decodeResult_fpExecutionType;
  assign queue_8_deq_bits_decodeResult_float = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_float : queue_dataOut_8_decodeResult_float;
  assign queue_8_deq_bits_decodeResult_specialSlot = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_specialSlot : queue_dataOut_8_decodeResult_specialSlot;
  assign queue_8_deq_bits_decodeResult_topUop = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_topUop : queue_dataOut_8_decodeResult_topUop;
  assign queue_8_deq_bits_decodeResult_popCount = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_popCount : queue_dataOut_8_decodeResult_popCount;
  assign queue_8_deq_bits_decodeResult_ffo = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_ffo : queue_dataOut_8_decodeResult_ffo;
  assign queue_8_deq_bits_decodeResult_average = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_average : queue_dataOut_8_decodeResult_average;
  assign queue_8_deq_bits_decodeResult_reverse = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_reverse : queue_dataOut_8_decodeResult_reverse;
  assign queue_8_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_8_decodeResult_dontNeedExecuteInLane;
  assign queue_8_deq_bits_decodeResult_scheduler = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_scheduler : queue_dataOut_8_decodeResult_scheduler;
  assign queue_8_deq_bits_decodeResult_sReadVD = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_sReadVD : queue_dataOut_8_decodeResult_sReadVD;
  assign queue_8_deq_bits_decodeResult_vtype = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_vtype : queue_dataOut_8_decodeResult_vtype;
  assign queue_8_deq_bits_decodeResult_sWrite = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_sWrite : queue_dataOut_8_decodeResult_sWrite;
  assign queue_8_deq_bits_decodeResult_crossRead = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_crossRead : queue_dataOut_8_decodeResult_crossRead;
  assign queue_8_deq_bits_decodeResult_crossWrite = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_crossWrite : queue_dataOut_8_decodeResult_crossWrite;
  assign queue_8_deq_bits_decodeResult_maskUnit = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_maskUnit : queue_dataOut_8_decodeResult_maskUnit;
  assign queue_8_deq_bits_decodeResult_special = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_special : queue_dataOut_8_decodeResult_special;
  assign queue_8_deq_bits_decodeResult_saturate = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_saturate : queue_dataOut_8_decodeResult_saturate;
  assign queue_8_deq_bits_decodeResult_vwmacc = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_vwmacc : queue_dataOut_8_decodeResult_vwmacc;
  assign queue_8_deq_bits_decodeResult_readOnly = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_readOnly : queue_dataOut_8_decodeResult_readOnly;
  assign queue_8_deq_bits_decodeResult_maskSource = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_maskSource : queue_dataOut_8_decodeResult_maskSource;
  assign queue_8_deq_bits_decodeResult_maskDestination = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_maskDestination : queue_dataOut_8_decodeResult_maskDestination;
  assign queue_8_deq_bits_decodeResult_maskLogic = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_maskLogic : queue_dataOut_8_decodeResult_maskLogic;
  assign queue_8_deq_bits_decodeResult_uop = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_uop : queue_dataOut_8_decodeResult_uop;
  assign queue_8_deq_bits_decodeResult_iota = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_iota : queue_dataOut_8_decodeResult_iota;
  assign queue_8_deq_bits_decodeResult_mv = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_mv : queue_dataOut_8_decodeResult_mv;
  assign queue_8_deq_bits_decodeResult_extend = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_extend : queue_dataOut_8_decodeResult_extend;
  assign queue_8_deq_bits_decodeResult_unOrderWrite = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_unOrderWrite : queue_dataOut_8_decodeResult_unOrderWrite;
  assign queue_8_deq_bits_decodeResult_compress = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_compress : queue_dataOut_8_decodeResult_compress;
  assign queue_8_deq_bits_decodeResult_gather16 = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_gather16 : queue_dataOut_8_decodeResult_gather16;
  assign queue_8_deq_bits_decodeResult_gather = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_gather : queue_dataOut_8_decodeResult_gather;
  assign queue_8_deq_bits_decodeResult_slid = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_slid : queue_dataOut_8_decodeResult_slid;
  assign queue_8_deq_bits_decodeResult_targetRd = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_targetRd : queue_dataOut_8_decodeResult_targetRd;
  assign queue_8_deq_bits_decodeResult_widenReduce = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_widenReduce : queue_dataOut_8_decodeResult_widenReduce;
  assign queue_8_deq_bits_decodeResult_red = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_red : queue_dataOut_8_decodeResult_red;
  assign queue_8_deq_bits_decodeResult_nr = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_nr : queue_dataOut_8_decodeResult_nr;
  assign queue_8_deq_bits_decodeResult_itype = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_itype : queue_dataOut_8_decodeResult_itype;
  assign queue_8_deq_bits_decodeResult_unsigned1 = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_unsigned1 : queue_dataOut_8_decodeResult_unsigned1;
  assign queue_8_deq_bits_decodeResult_unsigned0 = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_unsigned0 : queue_dataOut_8_decodeResult_unsigned0;
  assign queue_8_deq_bits_decodeResult_other = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_other : queue_dataOut_8_decodeResult_other;
  assign queue_8_deq_bits_decodeResult_multiCycle = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_multiCycle : queue_dataOut_8_decodeResult_multiCycle;
  assign queue_8_deq_bits_decodeResult_divider = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_divider : queue_dataOut_8_decodeResult_divider;
  assign queue_8_deq_bits_decodeResult_multiplier = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_multiplier : queue_dataOut_8_decodeResult_multiplier;
  assign queue_8_deq_bits_decodeResult_shift = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_shift : queue_dataOut_8_decodeResult_shift;
  assign queue_8_deq_bits_decodeResult_adder = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_adder : queue_dataOut_8_decodeResult_adder;
  assign queue_8_deq_bits_decodeResult_logic = _queue_fifo_8_empty ? queue_8_enq_bits_decodeResult_logic : queue_dataOut_8_decodeResult_logic;
  assign queue_8_deq_bits_loadStore = _queue_fifo_8_empty ? queue_8_enq_bits_loadStore : queue_dataOut_8_loadStore;
  assign queue_8_deq_bits_issueInst = _queue_fifo_8_empty ? queue_8_enq_bits_issueInst : queue_dataOut_8_issueInst;
  assign queue_8_deq_bits_store = _queue_fifo_8_empty ? queue_8_enq_bits_store : queue_dataOut_8_store;
  assign queue_8_deq_bits_special = _queue_fifo_8_empty ? queue_8_enq_bits_special : queue_dataOut_8_special;
  assign queue_8_deq_bits_lsWholeReg = _queue_fifo_8_empty ? queue_8_enq_bits_lsWholeReg : queue_dataOut_8_lsWholeReg;
  assign queue_8_deq_bits_vs1 = _queue_fifo_8_empty ? queue_8_enq_bits_vs1 : queue_dataOut_8_vs1;
  assign queue_8_deq_bits_vs2 = _queue_fifo_8_empty ? queue_8_enq_bits_vs2 : queue_dataOut_8_vs2;
  assign queue_8_deq_bits_vd = _queue_fifo_8_empty ? queue_8_enq_bits_vd : queue_dataOut_8_vd;
  assign queue_8_deq_bits_loadStoreEEW = _queue_fifo_8_empty ? queue_8_enq_bits_loadStoreEEW : queue_dataOut_8_loadStoreEEW;
  assign queue_8_deq_bits_mask = _queue_fifo_8_empty ? queue_8_enq_bits_mask : queue_dataOut_8_mask;
  assign queue_8_deq_bits_segment = _queue_fifo_8_empty ? queue_8_enq_bits_segment : queue_dataOut_8_segment;
  assign queue_8_deq_bits_readFromScalar = _queue_fifo_8_empty ? queue_8_enq_bits_readFromScalar : queue_dataOut_8_readFromScalar;
  assign queue_8_deq_bits_csrInterface_vl = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vl : queue_dataOut_8_csrInterface_vl;
  assign queue_8_deq_bits_csrInterface_vStart = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vStart : queue_dataOut_8_csrInterface_vStart;
  assign queue_8_deq_bits_csrInterface_vlmul = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vlmul : queue_dataOut_8_csrInterface_vlmul;
  assign queue_8_deq_bits_csrInterface_vSew = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vSew : queue_dataOut_8_csrInterface_vSew;
  assign queue_8_deq_bits_csrInterface_vxrm = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vxrm : queue_dataOut_8_csrInterface_vxrm;
  assign queue_8_deq_bits_csrInterface_vta = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vta : queue_dataOut_8_csrInterface_vta;
  assign queue_8_deq_bits_csrInterface_vma = _queue_fifo_8_empty ? queue_8_enq_bits_csrInterface_vma : queue_dataOut_8_csrInterface_vma;
  wire         laneVec_8_laneRequest_bits_issueInst = laneRequestSinkWire_8_ready & laneRequestSinkWire_8_valid;
  reg          releasePipe_pipe_v_8;
  wire         releasePipe_pipe_out_8_valid = releasePipe_pipe_v_8;
  wire         laneRequestSourceWire_8_ready;
  wire         validSource_8_valid = laneRequestSourceWire_8_ready & laneRequestSourceWire_8_valid;
  reg  [2:0]   tokenCheck_counter_8;
  wire [2:0]   tokenCheck_counterChange_8 = validSource_8_valid ? 3'h1 : 3'h7;
  assign tokenCheck_8 = ~(tokenCheck_counter_8[2]);
  assign laneRequestSourceWire_8_ready = tokenCheck_8;
  assign queue_8_enq_valid = validSink_8_valid;
  assign queue_8_enq_bits_instructionIndex = validSink_8_bits_instructionIndex;
  assign queue_8_enq_bits_decodeResult_orderReduce = validSink_8_bits_decodeResult_orderReduce;
  assign queue_8_enq_bits_decodeResult_floatMul = validSink_8_bits_decodeResult_floatMul;
  assign queue_8_enq_bits_decodeResult_fpExecutionType = validSink_8_bits_decodeResult_fpExecutionType;
  assign queue_8_enq_bits_decodeResult_float = validSink_8_bits_decodeResult_float;
  assign queue_8_enq_bits_decodeResult_specialSlot = validSink_8_bits_decodeResult_specialSlot;
  assign queue_8_enq_bits_decodeResult_topUop = validSink_8_bits_decodeResult_topUop;
  assign queue_8_enq_bits_decodeResult_popCount = validSink_8_bits_decodeResult_popCount;
  assign queue_8_enq_bits_decodeResult_ffo = validSink_8_bits_decodeResult_ffo;
  assign queue_8_enq_bits_decodeResult_average = validSink_8_bits_decodeResult_average;
  assign queue_8_enq_bits_decodeResult_reverse = validSink_8_bits_decodeResult_reverse;
  assign queue_8_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_8_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_8_enq_bits_decodeResult_scheduler = validSink_8_bits_decodeResult_scheduler;
  assign queue_8_enq_bits_decodeResult_sReadVD = validSink_8_bits_decodeResult_sReadVD;
  assign queue_8_enq_bits_decodeResult_vtype = validSink_8_bits_decodeResult_vtype;
  assign queue_8_enq_bits_decodeResult_sWrite = validSink_8_bits_decodeResult_sWrite;
  assign queue_8_enq_bits_decodeResult_crossRead = validSink_8_bits_decodeResult_crossRead;
  assign queue_8_enq_bits_decodeResult_crossWrite = validSink_8_bits_decodeResult_crossWrite;
  assign queue_8_enq_bits_decodeResult_maskUnit = validSink_8_bits_decodeResult_maskUnit;
  assign queue_8_enq_bits_decodeResult_special = validSink_8_bits_decodeResult_special;
  assign queue_8_enq_bits_decodeResult_saturate = validSink_8_bits_decodeResult_saturate;
  assign queue_8_enq_bits_decodeResult_vwmacc = validSink_8_bits_decodeResult_vwmacc;
  assign queue_8_enq_bits_decodeResult_readOnly = validSink_8_bits_decodeResult_readOnly;
  assign queue_8_enq_bits_decodeResult_maskSource = validSink_8_bits_decodeResult_maskSource;
  assign queue_8_enq_bits_decodeResult_maskDestination = validSink_8_bits_decodeResult_maskDestination;
  assign queue_8_enq_bits_decodeResult_maskLogic = validSink_8_bits_decodeResult_maskLogic;
  assign queue_8_enq_bits_decodeResult_uop = validSink_8_bits_decodeResult_uop;
  assign queue_8_enq_bits_decodeResult_iota = validSink_8_bits_decodeResult_iota;
  assign queue_8_enq_bits_decodeResult_mv = validSink_8_bits_decodeResult_mv;
  assign queue_8_enq_bits_decodeResult_extend = validSink_8_bits_decodeResult_extend;
  assign queue_8_enq_bits_decodeResult_unOrderWrite = validSink_8_bits_decodeResult_unOrderWrite;
  assign queue_8_enq_bits_decodeResult_compress = validSink_8_bits_decodeResult_compress;
  assign queue_8_enq_bits_decodeResult_gather16 = validSink_8_bits_decodeResult_gather16;
  assign queue_8_enq_bits_decodeResult_gather = validSink_8_bits_decodeResult_gather;
  assign queue_8_enq_bits_decodeResult_slid = validSink_8_bits_decodeResult_slid;
  assign queue_8_enq_bits_decodeResult_targetRd = validSink_8_bits_decodeResult_targetRd;
  assign queue_8_enq_bits_decodeResult_widenReduce = validSink_8_bits_decodeResult_widenReduce;
  assign queue_8_enq_bits_decodeResult_red = validSink_8_bits_decodeResult_red;
  assign queue_8_enq_bits_decodeResult_nr = validSink_8_bits_decodeResult_nr;
  assign queue_8_enq_bits_decodeResult_itype = validSink_8_bits_decodeResult_itype;
  assign queue_8_enq_bits_decodeResult_unsigned1 = validSink_8_bits_decodeResult_unsigned1;
  assign queue_8_enq_bits_decodeResult_unsigned0 = validSink_8_bits_decodeResult_unsigned0;
  assign queue_8_enq_bits_decodeResult_other = validSink_8_bits_decodeResult_other;
  assign queue_8_enq_bits_decodeResult_multiCycle = validSink_8_bits_decodeResult_multiCycle;
  assign queue_8_enq_bits_decodeResult_divider = validSink_8_bits_decodeResult_divider;
  assign queue_8_enq_bits_decodeResult_multiplier = validSink_8_bits_decodeResult_multiplier;
  assign queue_8_enq_bits_decodeResult_shift = validSink_8_bits_decodeResult_shift;
  assign queue_8_enq_bits_decodeResult_adder = validSink_8_bits_decodeResult_adder;
  assign queue_8_enq_bits_decodeResult_logic = validSink_8_bits_decodeResult_logic;
  assign queue_8_enq_bits_loadStore = validSink_8_bits_loadStore;
  assign queue_8_enq_bits_issueInst = validSink_8_bits_issueInst;
  assign queue_8_enq_bits_store = validSink_8_bits_store;
  assign queue_8_enq_bits_special = validSink_8_bits_special;
  assign queue_8_enq_bits_lsWholeReg = validSink_8_bits_lsWholeReg;
  assign queue_8_enq_bits_vs1 = validSink_8_bits_vs1;
  assign queue_8_enq_bits_vs2 = validSink_8_bits_vs2;
  assign queue_8_enq_bits_vd = validSink_8_bits_vd;
  assign queue_8_enq_bits_loadStoreEEW = validSink_8_bits_loadStoreEEW;
  assign queue_8_enq_bits_mask = validSink_8_bits_mask;
  assign queue_8_enq_bits_segment = validSink_8_bits_segment;
  assign queue_8_enq_bits_readFromScalar = validSink_8_bits_readFromScalar;
  assign queue_8_enq_bits_csrInterface_vl = validSink_8_bits_csrInterface_vl;
  assign queue_8_enq_bits_csrInterface_vStart = validSink_8_bits_csrInterface_vStart;
  assign queue_8_enq_bits_csrInterface_vlmul = validSink_8_bits_csrInterface_vlmul;
  assign queue_8_enq_bits_csrInterface_vSew = validSink_8_bits_csrInterface_vSew;
  assign queue_8_enq_bits_csrInterface_vxrm = validSink_8_bits_csrInterface_vxrm;
  assign queue_8_enq_bits_csrInterface_vta = validSink_8_bits_csrInterface_vta;
  assign queue_8_enq_bits_csrInterface_vma = validSink_8_bits_csrInterface_vma;
  reg          shifterReg_8_0_valid;
  assign validSink_8_valid = shifterReg_8_0_valid;
  reg  [2:0]   shifterReg_8_0_bits_instructionIndex;
  assign validSink_8_bits_instructionIndex = shifterReg_8_0_bits_instructionIndex;
  reg          shifterReg_8_0_bits_decodeResult_orderReduce;
  assign validSink_8_bits_decodeResult_orderReduce = shifterReg_8_0_bits_decodeResult_orderReduce;
  reg          shifterReg_8_0_bits_decodeResult_floatMul;
  assign validSink_8_bits_decodeResult_floatMul = shifterReg_8_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_8_0_bits_decodeResult_fpExecutionType;
  assign validSink_8_bits_decodeResult_fpExecutionType = shifterReg_8_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_8_0_bits_decodeResult_float;
  assign validSink_8_bits_decodeResult_float = shifterReg_8_0_bits_decodeResult_float;
  reg          shifterReg_8_0_bits_decodeResult_specialSlot;
  assign validSink_8_bits_decodeResult_specialSlot = shifterReg_8_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_8_0_bits_decodeResult_topUop;
  assign validSink_8_bits_decodeResult_topUop = shifterReg_8_0_bits_decodeResult_topUop;
  reg          shifterReg_8_0_bits_decodeResult_popCount;
  assign validSink_8_bits_decodeResult_popCount = shifterReg_8_0_bits_decodeResult_popCount;
  reg          shifterReg_8_0_bits_decodeResult_ffo;
  assign validSink_8_bits_decodeResult_ffo = shifterReg_8_0_bits_decodeResult_ffo;
  reg          shifterReg_8_0_bits_decodeResult_average;
  assign validSink_8_bits_decodeResult_average = shifterReg_8_0_bits_decodeResult_average;
  reg          shifterReg_8_0_bits_decodeResult_reverse;
  assign validSink_8_bits_decodeResult_reverse = shifterReg_8_0_bits_decodeResult_reverse;
  reg          shifterReg_8_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_8_bits_decodeResult_dontNeedExecuteInLane = shifterReg_8_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_8_0_bits_decodeResult_scheduler;
  assign validSink_8_bits_decodeResult_scheduler = shifterReg_8_0_bits_decodeResult_scheduler;
  reg          shifterReg_8_0_bits_decodeResult_sReadVD;
  assign validSink_8_bits_decodeResult_sReadVD = shifterReg_8_0_bits_decodeResult_sReadVD;
  reg          shifterReg_8_0_bits_decodeResult_vtype;
  assign validSink_8_bits_decodeResult_vtype = shifterReg_8_0_bits_decodeResult_vtype;
  reg          shifterReg_8_0_bits_decodeResult_sWrite;
  assign validSink_8_bits_decodeResult_sWrite = shifterReg_8_0_bits_decodeResult_sWrite;
  reg          shifterReg_8_0_bits_decodeResult_crossRead;
  assign validSink_8_bits_decodeResult_crossRead = shifterReg_8_0_bits_decodeResult_crossRead;
  reg          shifterReg_8_0_bits_decodeResult_crossWrite;
  assign validSink_8_bits_decodeResult_crossWrite = shifterReg_8_0_bits_decodeResult_crossWrite;
  reg          shifterReg_8_0_bits_decodeResult_maskUnit;
  assign validSink_8_bits_decodeResult_maskUnit = shifterReg_8_0_bits_decodeResult_maskUnit;
  reg          shifterReg_8_0_bits_decodeResult_special;
  assign validSink_8_bits_decodeResult_special = shifterReg_8_0_bits_decodeResult_special;
  reg          shifterReg_8_0_bits_decodeResult_saturate;
  assign validSink_8_bits_decodeResult_saturate = shifterReg_8_0_bits_decodeResult_saturate;
  reg          shifterReg_8_0_bits_decodeResult_vwmacc;
  assign validSink_8_bits_decodeResult_vwmacc = shifterReg_8_0_bits_decodeResult_vwmacc;
  reg          shifterReg_8_0_bits_decodeResult_readOnly;
  assign validSink_8_bits_decodeResult_readOnly = shifterReg_8_0_bits_decodeResult_readOnly;
  reg          shifterReg_8_0_bits_decodeResult_maskSource;
  assign validSink_8_bits_decodeResult_maskSource = shifterReg_8_0_bits_decodeResult_maskSource;
  reg          shifterReg_8_0_bits_decodeResult_maskDestination;
  assign validSink_8_bits_decodeResult_maskDestination = shifterReg_8_0_bits_decodeResult_maskDestination;
  reg          shifterReg_8_0_bits_decodeResult_maskLogic;
  assign validSink_8_bits_decodeResult_maskLogic = shifterReg_8_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_8_0_bits_decodeResult_uop;
  assign validSink_8_bits_decodeResult_uop = shifterReg_8_0_bits_decodeResult_uop;
  reg          shifterReg_8_0_bits_decodeResult_iota;
  assign validSink_8_bits_decodeResult_iota = shifterReg_8_0_bits_decodeResult_iota;
  reg          shifterReg_8_0_bits_decodeResult_mv;
  assign validSink_8_bits_decodeResult_mv = shifterReg_8_0_bits_decodeResult_mv;
  reg          shifterReg_8_0_bits_decodeResult_extend;
  assign validSink_8_bits_decodeResult_extend = shifterReg_8_0_bits_decodeResult_extend;
  reg          shifterReg_8_0_bits_decodeResult_unOrderWrite;
  assign validSink_8_bits_decodeResult_unOrderWrite = shifterReg_8_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_8_0_bits_decodeResult_compress;
  assign validSink_8_bits_decodeResult_compress = shifterReg_8_0_bits_decodeResult_compress;
  reg          shifterReg_8_0_bits_decodeResult_gather16;
  assign validSink_8_bits_decodeResult_gather16 = shifterReg_8_0_bits_decodeResult_gather16;
  reg          shifterReg_8_0_bits_decodeResult_gather;
  assign validSink_8_bits_decodeResult_gather = shifterReg_8_0_bits_decodeResult_gather;
  reg          shifterReg_8_0_bits_decodeResult_slid;
  assign validSink_8_bits_decodeResult_slid = shifterReg_8_0_bits_decodeResult_slid;
  reg          shifterReg_8_0_bits_decodeResult_targetRd;
  assign validSink_8_bits_decodeResult_targetRd = shifterReg_8_0_bits_decodeResult_targetRd;
  reg          shifterReg_8_0_bits_decodeResult_widenReduce;
  assign validSink_8_bits_decodeResult_widenReduce = shifterReg_8_0_bits_decodeResult_widenReduce;
  reg          shifterReg_8_0_bits_decodeResult_red;
  assign validSink_8_bits_decodeResult_red = shifterReg_8_0_bits_decodeResult_red;
  reg          shifterReg_8_0_bits_decodeResult_nr;
  assign validSink_8_bits_decodeResult_nr = shifterReg_8_0_bits_decodeResult_nr;
  reg          shifterReg_8_0_bits_decodeResult_itype;
  assign validSink_8_bits_decodeResult_itype = shifterReg_8_0_bits_decodeResult_itype;
  reg          shifterReg_8_0_bits_decodeResult_unsigned1;
  assign validSink_8_bits_decodeResult_unsigned1 = shifterReg_8_0_bits_decodeResult_unsigned1;
  reg          shifterReg_8_0_bits_decodeResult_unsigned0;
  assign validSink_8_bits_decodeResult_unsigned0 = shifterReg_8_0_bits_decodeResult_unsigned0;
  reg          shifterReg_8_0_bits_decodeResult_other;
  assign validSink_8_bits_decodeResult_other = shifterReg_8_0_bits_decodeResult_other;
  reg          shifterReg_8_0_bits_decodeResult_multiCycle;
  assign validSink_8_bits_decodeResult_multiCycle = shifterReg_8_0_bits_decodeResult_multiCycle;
  reg          shifterReg_8_0_bits_decodeResult_divider;
  assign validSink_8_bits_decodeResult_divider = shifterReg_8_0_bits_decodeResult_divider;
  reg          shifterReg_8_0_bits_decodeResult_multiplier;
  assign validSink_8_bits_decodeResult_multiplier = shifterReg_8_0_bits_decodeResult_multiplier;
  reg          shifterReg_8_0_bits_decodeResult_shift;
  assign validSink_8_bits_decodeResult_shift = shifterReg_8_0_bits_decodeResult_shift;
  reg          shifterReg_8_0_bits_decodeResult_adder;
  assign validSink_8_bits_decodeResult_adder = shifterReg_8_0_bits_decodeResult_adder;
  reg          shifterReg_8_0_bits_decodeResult_logic;
  assign validSink_8_bits_decodeResult_logic = shifterReg_8_0_bits_decodeResult_logic;
  reg          shifterReg_8_0_bits_loadStore;
  assign validSink_8_bits_loadStore = shifterReg_8_0_bits_loadStore;
  reg          shifterReg_8_0_bits_issueInst;
  assign validSink_8_bits_issueInst = shifterReg_8_0_bits_issueInst;
  reg          shifterReg_8_0_bits_store;
  assign validSink_8_bits_store = shifterReg_8_0_bits_store;
  reg          shifterReg_8_0_bits_special;
  assign validSink_8_bits_special = shifterReg_8_0_bits_special;
  reg          shifterReg_8_0_bits_lsWholeReg;
  assign validSink_8_bits_lsWholeReg = shifterReg_8_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_8_0_bits_vs1;
  assign validSink_8_bits_vs1 = shifterReg_8_0_bits_vs1;
  reg  [4:0]   shifterReg_8_0_bits_vs2;
  assign validSink_8_bits_vs2 = shifterReg_8_0_bits_vs2;
  reg  [4:0]   shifterReg_8_0_bits_vd;
  assign validSink_8_bits_vd = shifterReg_8_0_bits_vd;
  reg  [1:0]   shifterReg_8_0_bits_loadStoreEEW;
  assign validSink_8_bits_loadStoreEEW = shifterReg_8_0_bits_loadStoreEEW;
  reg          shifterReg_8_0_bits_mask;
  assign validSink_8_bits_mask = shifterReg_8_0_bits_mask;
  reg  [2:0]   shifterReg_8_0_bits_segment;
  assign validSink_8_bits_segment = shifterReg_8_0_bits_segment;
  reg  [31:0]  shifterReg_8_0_bits_readFromScalar;
  assign validSink_8_bits_readFromScalar = shifterReg_8_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_8_0_bits_csrInterface_vl;
  assign validSink_8_bits_csrInterface_vl = shifterReg_8_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_8_0_bits_csrInterface_vStart;
  assign validSink_8_bits_csrInterface_vStart = shifterReg_8_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_8_0_bits_csrInterface_vlmul;
  assign validSink_8_bits_csrInterface_vlmul = shifterReg_8_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_8_0_bits_csrInterface_vSew;
  assign validSink_8_bits_csrInterface_vSew = shifterReg_8_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_8_0_bits_csrInterface_vxrm;
  assign validSink_8_bits_csrInterface_vxrm = shifterReg_8_0_bits_csrInterface_vxrm;
  reg          shifterReg_8_0_bits_csrInterface_vta;
  assign validSink_8_bits_csrInterface_vta = shifterReg_8_0_bits_csrInterface_vta;
  reg          shifterReg_8_0_bits_csrInterface_vma;
  assign validSink_8_bits_csrInterface_vma = shifterReg_8_0_bits_csrInterface_vma;
  wire         shifterValid_8 = shifterReg_8_0_valid | validSource_8_valid;
  wire         validSink_9_valid;
  wire [2:0]   validSink_9_bits_instructionIndex;
  wire         validSink_9_bits_decodeResult_orderReduce;
  wire         validSink_9_bits_decodeResult_floatMul;
  wire [1:0]   validSink_9_bits_decodeResult_fpExecutionType;
  wire         validSink_9_bits_decodeResult_float;
  wire         validSink_9_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_9_bits_decodeResult_topUop;
  wire         validSink_9_bits_decodeResult_popCount;
  wire         validSink_9_bits_decodeResult_ffo;
  wire         validSink_9_bits_decodeResult_average;
  wire         validSink_9_bits_decodeResult_reverse;
  wire         validSink_9_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_9_bits_decodeResult_scheduler;
  wire         validSink_9_bits_decodeResult_sReadVD;
  wire         validSink_9_bits_decodeResult_vtype;
  wire         validSink_9_bits_decodeResult_sWrite;
  wire         validSink_9_bits_decodeResult_crossRead;
  wire         validSink_9_bits_decodeResult_crossWrite;
  wire         validSink_9_bits_decodeResult_maskUnit;
  wire         validSink_9_bits_decodeResult_special;
  wire         validSink_9_bits_decodeResult_saturate;
  wire         validSink_9_bits_decodeResult_vwmacc;
  wire         validSink_9_bits_decodeResult_readOnly;
  wire         validSink_9_bits_decodeResult_maskSource;
  wire         validSink_9_bits_decodeResult_maskDestination;
  wire         validSink_9_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_9_bits_decodeResult_uop;
  wire         validSink_9_bits_decodeResult_iota;
  wire         validSink_9_bits_decodeResult_mv;
  wire         validSink_9_bits_decodeResult_extend;
  wire         validSink_9_bits_decodeResult_unOrderWrite;
  wire         validSink_9_bits_decodeResult_compress;
  wire         validSink_9_bits_decodeResult_gather16;
  wire         validSink_9_bits_decodeResult_gather;
  wire         validSink_9_bits_decodeResult_slid;
  wire         validSink_9_bits_decodeResult_targetRd;
  wire         validSink_9_bits_decodeResult_widenReduce;
  wire         validSink_9_bits_decodeResult_red;
  wire         validSink_9_bits_decodeResult_nr;
  wire         validSink_9_bits_decodeResult_itype;
  wire         validSink_9_bits_decodeResult_unsigned1;
  wire         validSink_9_bits_decodeResult_unsigned0;
  wire         validSink_9_bits_decodeResult_other;
  wire         validSink_9_bits_decodeResult_multiCycle;
  wire         validSink_9_bits_decodeResult_divider;
  wire         validSink_9_bits_decodeResult_multiplier;
  wire         validSink_9_bits_decodeResult_shift;
  wire         validSink_9_bits_decodeResult_adder;
  wire         validSink_9_bits_decodeResult_logic;
  wire         validSink_9_bits_loadStore;
  wire         validSink_9_bits_issueInst;
  wire         validSink_9_bits_store;
  wire         validSink_9_bits_special;
  wire         validSink_9_bits_lsWholeReg;
  wire [4:0]   validSink_9_bits_vs1;
  wire [4:0]   validSink_9_bits_vs2;
  wire [4:0]   validSink_9_bits_vd;
  wire [1:0]   validSink_9_bits_loadStoreEEW;
  wire         validSink_9_bits_mask;
  wire [2:0]   validSink_9_bits_segment;
  wire [31:0]  validSink_9_bits_readFromScalar;
  wire [11:0]  validSink_9_bits_csrInterface_vl;
  wire [11:0]  validSink_9_bits_csrInterface_vStart;
  wire [2:0]   validSink_9_bits_csrInterface_vlmul;
  wire [1:0]   validSink_9_bits_csrInterface_vSew;
  wire [1:0]   validSink_9_bits_csrInterface_vxrm;
  wire         validSink_9_bits_csrInterface_vta;
  wire         validSink_9_bits_csrInterface_vma;
  wire         laneRequestSinkWire_9_valid = queue_9_deq_valid;
  wire [2:0]   laneRequestSinkWire_9_bits_instructionIndex = queue_9_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_9_bits_decodeResult_orderReduce = queue_9_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_9_bits_decodeResult_floatMul = queue_9_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_9_bits_decodeResult_fpExecutionType = queue_9_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_9_bits_decodeResult_float = queue_9_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_9_bits_decodeResult_specialSlot = queue_9_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_9_bits_decodeResult_topUop = queue_9_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_9_bits_decodeResult_popCount = queue_9_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_9_bits_decodeResult_ffo = queue_9_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_9_bits_decodeResult_average = queue_9_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_9_bits_decodeResult_reverse = queue_9_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_9_bits_decodeResult_dontNeedExecuteInLane = queue_9_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_9_bits_decodeResult_scheduler = queue_9_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_9_bits_decodeResult_sReadVD = queue_9_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_9_bits_decodeResult_vtype = queue_9_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_9_bits_decodeResult_sWrite = queue_9_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_9_bits_decodeResult_crossRead = queue_9_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_9_bits_decodeResult_crossWrite = queue_9_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_9_bits_decodeResult_maskUnit = queue_9_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_9_bits_decodeResult_special = queue_9_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_9_bits_decodeResult_saturate = queue_9_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_9_bits_decodeResult_vwmacc = queue_9_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_9_bits_decodeResult_readOnly = queue_9_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_9_bits_decodeResult_maskSource = queue_9_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_9_bits_decodeResult_maskDestination = queue_9_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_9_bits_decodeResult_maskLogic = queue_9_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_9_bits_decodeResult_uop = queue_9_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_9_bits_decodeResult_iota = queue_9_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_9_bits_decodeResult_mv = queue_9_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_9_bits_decodeResult_extend = queue_9_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_9_bits_decodeResult_unOrderWrite = queue_9_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_9_bits_decodeResult_compress = queue_9_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_9_bits_decodeResult_gather16 = queue_9_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_9_bits_decodeResult_gather = queue_9_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_9_bits_decodeResult_slid = queue_9_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_9_bits_decodeResult_targetRd = queue_9_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_9_bits_decodeResult_widenReduce = queue_9_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_9_bits_decodeResult_red = queue_9_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_9_bits_decodeResult_nr = queue_9_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_9_bits_decodeResult_itype = queue_9_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_9_bits_decodeResult_unsigned1 = queue_9_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_9_bits_decodeResult_unsigned0 = queue_9_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_9_bits_decodeResult_other = queue_9_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_9_bits_decodeResult_multiCycle = queue_9_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_9_bits_decodeResult_divider = queue_9_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_9_bits_decodeResult_multiplier = queue_9_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_9_bits_decodeResult_shift = queue_9_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_9_bits_decodeResult_adder = queue_9_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_9_bits_decodeResult_logic = queue_9_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_9_bits_loadStore = queue_9_deq_bits_loadStore;
  wire         laneRequestSinkWire_9_bits_issueInst = queue_9_deq_bits_issueInst;
  wire         laneRequestSinkWire_9_bits_store = queue_9_deq_bits_store;
  wire         laneRequestSinkWire_9_bits_special = queue_9_deq_bits_special;
  wire         laneRequestSinkWire_9_bits_lsWholeReg = queue_9_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_9_bits_vs1 = queue_9_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_9_bits_vs2 = queue_9_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_9_bits_vd = queue_9_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_9_bits_loadStoreEEW = queue_9_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_9_bits_mask = queue_9_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_9_bits_segment = queue_9_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_9_bits_readFromScalar = queue_9_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_9_bits_csrInterface_vl = queue_9_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_9_bits_csrInterface_vStart = queue_9_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_9_bits_csrInterface_vlmul = queue_9_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_9_bits_csrInterface_vSew = queue_9_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_9_bits_csrInterface_vxrm = queue_9_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_9_bits_csrInterface_vta = queue_9_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_9_bits_csrInterface_vma = queue_9_deq_bits_csrInterface_vma;
  wire [1:0]   queue_9_enq_bits_csrInterface_vxrm;
  wire         queue_9_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_27 = {queue_9_enq_bits_csrInterface_vxrm, queue_9_enq_bits_csrInterface_vta};
  wire         queue_9_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_27 = {queue_dataIn_lo_hi_27, queue_9_enq_bits_csrInterface_vma};
  wire [2:0]   queue_9_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_9_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_27 = {queue_9_enq_bits_csrInterface_vlmul, queue_9_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_9_enq_bits_csrInterface_vl;
  wire [11:0]  queue_9_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_27 = {queue_9_enq_bits_csrInterface_vl, queue_9_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_27 = {queue_dataIn_hi_hi_27, queue_dataIn_hi_lo_27};
  wire         queue_9_enq_bits_decodeResult_shift;
  wire         queue_9_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_9 = {queue_9_enq_bits_decodeResult_shift, queue_9_enq_bits_decodeResult_adder};
  wire         queue_9_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_9 = {queue_dataIn_lo_lo_lo_lo_hi_9, queue_9_enq_bits_decodeResult_logic};
  wire         queue_9_enq_bits_decodeResult_multiCycle;
  wire         queue_9_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_9 = {queue_9_enq_bits_decodeResult_multiCycle, queue_9_enq_bits_decodeResult_divider};
  wire         queue_9_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_9 = {queue_dataIn_lo_lo_lo_hi_hi_9, queue_9_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_9 = {queue_dataIn_lo_lo_lo_hi_9, queue_dataIn_lo_lo_lo_lo_9};
  wire         queue_9_enq_bits_decodeResult_unsigned1;
  wire         queue_9_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_9 = {queue_9_enq_bits_decodeResult_unsigned1, queue_9_enq_bits_decodeResult_unsigned0};
  wire         queue_9_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_9 = {queue_dataIn_lo_lo_hi_lo_hi_9, queue_9_enq_bits_decodeResult_other};
  wire         queue_9_enq_bits_decodeResult_red;
  wire         queue_9_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_9 = {queue_9_enq_bits_decodeResult_red, queue_9_enq_bits_decodeResult_nr};
  wire         queue_9_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_9 = {queue_dataIn_lo_lo_hi_hi_hi_9, queue_9_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_18 = {queue_dataIn_lo_lo_hi_hi_9, queue_dataIn_lo_lo_hi_lo_9};
  wire [11:0]  queue_dataIn_lo_lo_18 = {queue_dataIn_lo_lo_hi_18, queue_dataIn_lo_lo_lo_9};
  wire         queue_9_enq_bits_decodeResult_slid;
  wire         queue_9_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_9 = {queue_9_enq_bits_decodeResult_slid, queue_9_enq_bits_decodeResult_targetRd};
  wire         queue_9_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_9 = {queue_dataIn_lo_hi_lo_lo_hi_9, queue_9_enq_bits_decodeResult_widenReduce};
  wire         queue_9_enq_bits_decodeResult_compress;
  wire         queue_9_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_9 = {queue_9_enq_bits_decodeResult_compress, queue_9_enq_bits_decodeResult_gather16};
  wire         queue_9_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_9 = {queue_dataIn_lo_hi_lo_hi_hi_9, queue_9_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_18 = {queue_dataIn_lo_hi_lo_hi_9, queue_dataIn_lo_hi_lo_lo_9};
  wire         queue_9_enq_bits_decodeResult_mv;
  wire         queue_9_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_9 = {queue_9_enq_bits_decodeResult_mv, queue_9_enq_bits_decodeResult_extend};
  wire         queue_9_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_9 = {queue_dataIn_lo_hi_hi_lo_hi_9, queue_9_enq_bits_decodeResult_unOrderWrite};
  wire         queue_9_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_9_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_9 = {queue_9_enq_bits_decodeResult_maskLogic, queue_9_enq_bits_decodeResult_uop};
  wire         queue_9_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_9 = {queue_dataIn_lo_hi_hi_hi_hi_9, queue_9_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_18 = {queue_dataIn_lo_hi_hi_hi_9, queue_dataIn_lo_hi_hi_lo_9};
  wire [14:0]  queue_dataIn_lo_hi_28 = {queue_dataIn_lo_hi_hi_18, queue_dataIn_lo_hi_lo_18};
  wire [26:0]  queue_dataIn_lo_28 = {queue_dataIn_lo_hi_28, queue_dataIn_lo_lo_18};
  wire         queue_9_enq_bits_decodeResult_readOnly;
  wire         queue_9_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_9 = {queue_9_enq_bits_decodeResult_readOnly, queue_9_enq_bits_decodeResult_maskSource};
  wire         queue_9_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_9 = {queue_dataIn_hi_lo_lo_lo_hi_9, queue_9_enq_bits_decodeResult_maskDestination};
  wire         queue_9_enq_bits_decodeResult_special;
  wire         queue_9_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_9 = {queue_9_enq_bits_decodeResult_special, queue_9_enq_bits_decodeResult_saturate};
  wire         queue_9_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_9 = {queue_dataIn_hi_lo_lo_hi_hi_9, queue_9_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_18 = {queue_dataIn_hi_lo_lo_hi_9, queue_dataIn_hi_lo_lo_lo_9};
  wire         queue_9_enq_bits_decodeResult_crossRead;
  wire         queue_9_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_9 = {queue_9_enq_bits_decodeResult_crossRead, queue_9_enq_bits_decodeResult_crossWrite};
  wire         queue_9_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_9 = {queue_dataIn_hi_lo_hi_lo_hi_9, queue_9_enq_bits_decodeResult_maskUnit};
  wire         queue_9_enq_bits_decodeResult_sReadVD;
  wire         queue_9_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_9 = {queue_9_enq_bits_decodeResult_sReadVD, queue_9_enq_bits_decodeResult_vtype};
  wire         queue_9_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_9 = {queue_dataIn_hi_lo_hi_hi_hi_9, queue_9_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_18 = {queue_dataIn_hi_lo_hi_hi_9, queue_dataIn_hi_lo_hi_lo_9};
  wire [11:0]  queue_dataIn_hi_lo_28 = {queue_dataIn_hi_lo_hi_18, queue_dataIn_hi_lo_lo_18};
  wire         queue_9_enq_bits_decodeResult_reverse;
  wire         queue_9_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_9 = {queue_9_enq_bits_decodeResult_reverse, queue_9_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_9_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_9 = {queue_dataIn_hi_hi_lo_lo_hi_9, queue_9_enq_bits_decodeResult_scheduler};
  wire         queue_9_enq_bits_decodeResult_popCount;
  wire         queue_9_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_9 = {queue_9_enq_bits_decodeResult_popCount, queue_9_enq_bits_decodeResult_ffo};
  wire         queue_9_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_9 = {queue_dataIn_hi_hi_lo_hi_hi_9, queue_9_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_18 = {queue_dataIn_hi_hi_lo_hi_9, queue_dataIn_hi_hi_lo_lo_9};
  wire         queue_9_enq_bits_decodeResult_float;
  wire         queue_9_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_9 = {queue_9_enq_bits_decodeResult_float, queue_9_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_9_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_9 = {queue_dataIn_hi_hi_hi_lo_hi_9, queue_9_enq_bits_decodeResult_topUop};
  wire         queue_9_enq_bits_decodeResult_orderReduce;
  wire         queue_9_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_9 = {queue_9_enq_bits_decodeResult_orderReduce, queue_9_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_9_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_9 = {queue_dataIn_hi_hi_hi_hi_hi_9, queue_9_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_18 = {queue_dataIn_hi_hi_hi_hi_9, queue_dataIn_hi_hi_hi_lo_9};
  wire [16:0]  queue_dataIn_hi_hi_28 = {queue_dataIn_hi_hi_hi_18, queue_dataIn_hi_hi_lo_18};
  wire [28:0]  queue_dataIn_hi_28 = {queue_dataIn_hi_hi_28, queue_dataIn_hi_lo_28};
  wire [2:0]   queue_9_enq_bits_segment;
  wire [31:0]  queue_9_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_19 = {queue_9_enq_bits_segment, queue_9_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_19 = {queue_dataIn_lo_lo_hi_19, queue_dataIn_hi_27, queue_dataIn_lo_27};
  wire [1:0]   queue_9_enq_bits_loadStoreEEW;
  wire         queue_9_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_19 = {queue_9_enq_bits_loadStoreEEW, queue_9_enq_bits_mask};
  wire [4:0]   queue_9_enq_bits_vs2;
  wire [4:0]   queue_9_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_19 = {queue_9_enq_bits_vs2, queue_9_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_29 = {queue_dataIn_lo_hi_hi_19, queue_dataIn_lo_hi_lo_19};
  wire [80:0]  queue_dataIn_lo_29 = {queue_dataIn_lo_hi_29, queue_dataIn_lo_lo_19};
  wire         queue_9_enq_bits_lsWholeReg;
  wire [4:0]   queue_9_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_19 = {queue_9_enq_bits_lsWholeReg, queue_9_enq_bits_vs1};
  wire         queue_9_enq_bits_store;
  wire         queue_9_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_19 = {queue_9_enq_bits_store, queue_9_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_29 = {queue_dataIn_hi_lo_hi_19, queue_dataIn_hi_lo_lo_19};
  wire         queue_9_enq_bits_loadStore;
  wire         queue_9_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_19 = {queue_9_enq_bits_loadStore, queue_9_enq_bits_issueInst};
  wire [2:0]   queue_9_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_19 = {queue_9_enq_bits_instructionIndex, queue_dataIn_hi_28, queue_dataIn_lo_28};
  wire [60:0]  queue_dataIn_hi_hi_29 = {queue_dataIn_hi_hi_hi_19, queue_dataIn_hi_hi_lo_19};
  wire [68:0]  queue_dataIn_hi_29 = {queue_dataIn_hi_hi_29, queue_dataIn_hi_lo_29};
  wire [149:0] queue_dataIn_9 = {queue_dataIn_hi_29, queue_dataIn_lo_29};
  wire         queue_dataOut_9_csrInterface_vma = _queue_fifo_9_data_out[0];
  wire         queue_dataOut_9_csrInterface_vta = _queue_fifo_9_data_out[1];
  wire [1:0]   queue_dataOut_9_csrInterface_vxrm = _queue_fifo_9_data_out[3:2];
  wire [1:0]   queue_dataOut_9_csrInterface_vSew = _queue_fifo_9_data_out[5:4];
  wire [2:0]   queue_dataOut_9_csrInterface_vlmul = _queue_fifo_9_data_out[8:6];
  wire [11:0]  queue_dataOut_9_csrInterface_vStart = _queue_fifo_9_data_out[20:9];
  wire [11:0]  queue_dataOut_9_csrInterface_vl = _queue_fifo_9_data_out[32:21];
  wire [31:0]  queue_dataOut_9_readFromScalar = _queue_fifo_9_data_out[64:33];
  wire [2:0]   queue_dataOut_9_segment = _queue_fifo_9_data_out[67:65];
  wire         queue_dataOut_9_mask = _queue_fifo_9_data_out[68];
  wire [1:0]   queue_dataOut_9_loadStoreEEW = _queue_fifo_9_data_out[70:69];
  wire [4:0]   queue_dataOut_9_vd = _queue_fifo_9_data_out[75:71];
  wire [4:0]   queue_dataOut_9_vs2 = _queue_fifo_9_data_out[80:76];
  wire [4:0]   queue_dataOut_9_vs1 = _queue_fifo_9_data_out[85:81];
  wire         queue_dataOut_9_lsWholeReg = _queue_fifo_9_data_out[86];
  wire         queue_dataOut_9_special = _queue_fifo_9_data_out[87];
  wire         queue_dataOut_9_store = _queue_fifo_9_data_out[88];
  wire         queue_dataOut_9_issueInst = _queue_fifo_9_data_out[89];
  wire         queue_dataOut_9_loadStore = _queue_fifo_9_data_out[90];
  wire         queue_dataOut_9_decodeResult_logic = _queue_fifo_9_data_out[91];
  wire         queue_dataOut_9_decodeResult_adder = _queue_fifo_9_data_out[92];
  wire         queue_dataOut_9_decodeResult_shift = _queue_fifo_9_data_out[93];
  wire         queue_dataOut_9_decodeResult_multiplier = _queue_fifo_9_data_out[94];
  wire         queue_dataOut_9_decodeResult_divider = _queue_fifo_9_data_out[95];
  wire         queue_dataOut_9_decodeResult_multiCycle = _queue_fifo_9_data_out[96];
  wire         queue_dataOut_9_decodeResult_other = _queue_fifo_9_data_out[97];
  wire         queue_dataOut_9_decodeResult_unsigned0 = _queue_fifo_9_data_out[98];
  wire         queue_dataOut_9_decodeResult_unsigned1 = _queue_fifo_9_data_out[99];
  wire         queue_dataOut_9_decodeResult_itype = _queue_fifo_9_data_out[100];
  wire         queue_dataOut_9_decodeResult_nr = _queue_fifo_9_data_out[101];
  wire         queue_dataOut_9_decodeResult_red = _queue_fifo_9_data_out[102];
  wire         queue_dataOut_9_decodeResult_widenReduce = _queue_fifo_9_data_out[103];
  wire         queue_dataOut_9_decodeResult_targetRd = _queue_fifo_9_data_out[104];
  wire         queue_dataOut_9_decodeResult_slid = _queue_fifo_9_data_out[105];
  wire         queue_dataOut_9_decodeResult_gather = _queue_fifo_9_data_out[106];
  wire         queue_dataOut_9_decodeResult_gather16 = _queue_fifo_9_data_out[107];
  wire         queue_dataOut_9_decodeResult_compress = _queue_fifo_9_data_out[108];
  wire         queue_dataOut_9_decodeResult_unOrderWrite = _queue_fifo_9_data_out[109];
  wire         queue_dataOut_9_decodeResult_extend = _queue_fifo_9_data_out[110];
  wire         queue_dataOut_9_decodeResult_mv = _queue_fifo_9_data_out[111];
  wire         queue_dataOut_9_decodeResult_iota = _queue_fifo_9_data_out[112];
  wire [3:0]   queue_dataOut_9_decodeResult_uop = _queue_fifo_9_data_out[116:113];
  wire         queue_dataOut_9_decodeResult_maskLogic = _queue_fifo_9_data_out[117];
  wire         queue_dataOut_9_decodeResult_maskDestination = _queue_fifo_9_data_out[118];
  wire         queue_dataOut_9_decodeResult_maskSource = _queue_fifo_9_data_out[119];
  wire         queue_dataOut_9_decodeResult_readOnly = _queue_fifo_9_data_out[120];
  wire         queue_dataOut_9_decodeResult_vwmacc = _queue_fifo_9_data_out[121];
  wire         queue_dataOut_9_decodeResult_saturate = _queue_fifo_9_data_out[122];
  wire         queue_dataOut_9_decodeResult_special = _queue_fifo_9_data_out[123];
  wire         queue_dataOut_9_decodeResult_maskUnit = _queue_fifo_9_data_out[124];
  wire         queue_dataOut_9_decodeResult_crossWrite = _queue_fifo_9_data_out[125];
  wire         queue_dataOut_9_decodeResult_crossRead = _queue_fifo_9_data_out[126];
  wire         queue_dataOut_9_decodeResult_sWrite = _queue_fifo_9_data_out[127];
  wire         queue_dataOut_9_decodeResult_vtype = _queue_fifo_9_data_out[128];
  wire         queue_dataOut_9_decodeResult_sReadVD = _queue_fifo_9_data_out[129];
  wire         queue_dataOut_9_decodeResult_scheduler = _queue_fifo_9_data_out[130];
  wire         queue_dataOut_9_decodeResult_dontNeedExecuteInLane = _queue_fifo_9_data_out[131];
  wire         queue_dataOut_9_decodeResult_reverse = _queue_fifo_9_data_out[132];
  wire         queue_dataOut_9_decodeResult_average = _queue_fifo_9_data_out[133];
  wire         queue_dataOut_9_decodeResult_ffo = _queue_fifo_9_data_out[134];
  wire         queue_dataOut_9_decodeResult_popCount = _queue_fifo_9_data_out[135];
  wire [4:0]   queue_dataOut_9_decodeResult_topUop = _queue_fifo_9_data_out[140:136];
  wire         queue_dataOut_9_decodeResult_specialSlot = _queue_fifo_9_data_out[141];
  wire         queue_dataOut_9_decodeResult_float = _queue_fifo_9_data_out[142];
  wire [1:0]   queue_dataOut_9_decodeResult_fpExecutionType = _queue_fifo_9_data_out[144:143];
  wire         queue_dataOut_9_decodeResult_floatMul = _queue_fifo_9_data_out[145];
  wire         queue_dataOut_9_decodeResult_orderReduce = _queue_fifo_9_data_out[146];
  wire [2:0]   queue_dataOut_9_instructionIndex = _queue_fifo_9_data_out[149:147];
  wire         queue_9_enq_ready = ~_queue_fifo_9_full;
  wire         queue_9_enq_valid;
  assign queue_9_deq_valid = ~_queue_fifo_9_empty | queue_9_enq_valid;
  assign queue_9_deq_bits_instructionIndex = _queue_fifo_9_empty ? queue_9_enq_bits_instructionIndex : queue_dataOut_9_instructionIndex;
  assign queue_9_deq_bits_decodeResult_orderReduce = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_orderReduce : queue_dataOut_9_decodeResult_orderReduce;
  assign queue_9_deq_bits_decodeResult_floatMul = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_floatMul : queue_dataOut_9_decodeResult_floatMul;
  assign queue_9_deq_bits_decodeResult_fpExecutionType = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_fpExecutionType : queue_dataOut_9_decodeResult_fpExecutionType;
  assign queue_9_deq_bits_decodeResult_float = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_float : queue_dataOut_9_decodeResult_float;
  assign queue_9_deq_bits_decodeResult_specialSlot = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_specialSlot : queue_dataOut_9_decodeResult_specialSlot;
  assign queue_9_deq_bits_decodeResult_topUop = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_topUop : queue_dataOut_9_decodeResult_topUop;
  assign queue_9_deq_bits_decodeResult_popCount = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_popCount : queue_dataOut_9_decodeResult_popCount;
  assign queue_9_deq_bits_decodeResult_ffo = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_ffo : queue_dataOut_9_decodeResult_ffo;
  assign queue_9_deq_bits_decodeResult_average = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_average : queue_dataOut_9_decodeResult_average;
  assign queue_9_deq_bits_decodeResult_reverse = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_reverse : queue_dataOut_9_decodeResult_reverse;
  assign queue_9_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_9_decodeResult_dontNeedExecuteInLane;
  assign queue_9_deq_bits_decodeResult_scheduler = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_scheduler : queue_dataOut_9_decodeResult_scheduler;
  assign queue_9_deq_bits_decodeResult_sReadVD = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_sReadVD : queue_dataOut_9_decodeResult_sReadVD;
  assign queue_9_deq_bits_decodeResult_vtype = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_vtype : queue_dataOut_9_decodeResult_vtype;
  assign queue_9_deq_bits_decodeResult_sWrite = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_sWrite : queue_dataOut_9_decodeResult_sWrite;
  assign queue_9_deq_bits_decodeResult_crossRead = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_crossRead : queue_dataOut_9_decodeResult_crossRead;
  assign queue_9_deq_bits_decodeResult_crossWrite = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_crossWrite : queue_dataOut_9_decodeResult_crossWrite;
  assign queue_9_deq_bits_decodeResult_maskUnit = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_maskUnit : queue_dataOut_9_decodeResult_maskUnit;
  assign queue_9_deq_bits_decodeResult_special = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_special : queue_dataOut_9_decodeResult_special;
  assign queue_9_deq_bits_decodeResult_saturate = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_saturate : queue_dataOut_9_decodeResult_saturate;
  assign queue_9_deq_bits_decodeResult_vwmacc = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_vwmacc : queue_dataOut_9_decodeResult_vwmacc;
  assign queue_9_deq_bits_decodeResult_readOnly = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_readOnly : queue_dataOut_9_decodeResult_readOnly;
  assign queue_9_deq_bits_decodeResult_maskSource = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_maskSource : queue_dataOut_9_decodeResult_maskSource;
  assign queue_9_deq_bits_decodeResult_maskDestination = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_maskDestination : queue_dataOut_9_decodeResult_maskDestination;
  assign queue_9_deq_bits_decodeResult_maskLogic = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_maskLogic : queue_dataOut_9_decodeResult_maskLogic;
  assign queue_9_deq_bits_decodeResult_uop = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_uop : queue_dataOut_9_decodeResult_uop;
  assign queue_9_deq_bits_decodeResult_iota = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_iota : queue_dataOut_9_decodeResult_iota;
  assign queue_9_deq_bits_decodeResult_mv = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_mv : queue_dataOut_9_decodeResult_mv;
  assign queue_9_deq_bits_decodeResult_extend = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_extend : queue_dataOut_9_decodeResult_extend;
  assign queue_9_deq_bits_decodeResult_unOrderWrite = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_unOrderWrite : queue_dataOut_9_decodeResult_unOrderWrite;
  assign queue_9_deq_bits_decodeResult_compress = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_compress : queue_dataOut_9_decodeResult_compress;
  assign queue_9_deq_bits_decodeResult_gather16 = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_gather16 : queue_dataOut_9_decodeResult_gather16;
  assign queue_9_deq_bits_decodeResult_gather = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_gather : queue_dataOut_9_decodeResult_gather;
  assign queue_9_deq_bits_decodeResult_slid = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_slid : queue_dataOut_9_decodeResult_slid;
  assign queue_9_deq_bits_decodeResult_targetRd = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_targetRd : queue_dataOut_9_decodeResult_targetRd;
  assign queue_9_deq_bits_decodeResult_widenReduce = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_widenReduce : queue_dataOut_9_decodeResult_widenReduce;
  assign queue_9_deq_bits_decodeResult_red = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_red : queue_dataOut_9_decodeResult_red;
  assign queue_9_deq_bits_decodeResult_nr = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_nr : queue_dataOut_9_decodeResult_nr;
  assign queue_9_deq_bits_decodeResult_itype = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_itype : queue_dataOut_9_decodeResult_itype;
  assign queue_9_deq_bits_decodeResult_unsigned1 = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_unsigned1 : queue_dataOut_9_decodeResult_unsigned1;
  assign queue_9_deq_bits_decodeResult_unsigned0 = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_unsigned0 : queue_dataOut_9_decodeResult_unsigned0;
  assign queue_9_deq_bits_decodeResult_other = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_other : queue_dataOut_9_decodeResult_other;
  assign queue_9_deq_bits_decodeResult_multiCycle = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_multiCycle : queue_dataOut_9_decodeResult_multiCycle;
  assign queue_9_deq_bits_decodeResult_divider = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_divider : queue_dataOut_9_decodeResult_divider;
  assign queue_9_deq_bits_decodeResult_multiplier = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_multiplier : queue_dataOut_9_decodeResult_multiplier;
  assign queue_9_deq_bits_decodeResult_shift = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_shift : queue_dataOut_9_decodeResult_shift;
  assign queue_9_deq_bits_decodeResult_adder = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_adder : queue_dataOut_9_decodeResult_adder;
  assign queue_9_deq_bits_decodeResult_logic = _queue_fifo_9_empty ? queue_9_enq_bits_decodeResult_logic : queue_dataOut_9_decodeResult_logic;
  assign queue_9_deq_bits_loadStore = _queue_fifo_9_empty ? queue_9_enq_bits_loadStore : queue_dataOut_9_loadStore;
  assign queue_9_deq_bits_issueInst = _queue_fifo_9_empty ? queue_9_enq_bits_issueInst : queue_dataOut_9_issueInst;
  assign queue_9_deq_bits_store = _queue_fifo_9_empty ? queue_9_enq_bits_store : queue_dataOut_9_store;
  assign queue_9_deq_bits_special = _queue_fifo_9_empty ? queue_9_enq_bits_special : queue_dataOut_9_special;
  assign queue_9_deq_bits_lsWholeReg = _queue_fifo_9_empty ? queue_9_enq_bits_lsWholeReg : queue_dataOut_9_lsWholeReg;
  assign queue_9_deq_bits_vs1 = _queue_fifo_9_empty ? queue_9_enq_bits_vs1 : queue_dataOut_9_vs1;
  assign queue_9_deq_bits_vs2 = _queue_fifo_9_empty ? queue_9_enq_bits_vs2 : queue_dataOut_9_vs2;
  assign queue_9_deq_bits_vd = _queue_fifo_9_empty ? queue_9_enq_bits_vd : queue_dataOut_9_vd;
  assign queue_9_deq_bits_loadStoreEEW = _queue_fifo_9_empty ? queue_9_enq_bits_loadStoreEEW : queue_dataOut_9_loadStoreEEW;
  assign queue_9_deq_bits_mask = _queue_fifo_9_empty ? queue_9_enq_bits_mask : queue_dataOut_9_mask;
  assign queue_9_deq_bits_segment = _queue_fifo_9_empty ? queue_9_enq_bits_segment : queue_dataOut_9_segment;
  assign queue_9_deq_bits_readFromScalar = _queue_fifo_9_empty ? queue_9_enq_bits_readFromScalar : queue_dataOut_9_readFromScalar;
  assign queue_9_deq_bits_csrInterface_vl = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vl : queue_dataOut_9_csrInterface_vl;
  assign queue_9_deq_bits_csrInterface_vStart = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vStart : queue_dataOut_9_csrInterface_vStart;
  assign queue_9_deq_bits_csrInterface_vlmul = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vlmul : queue_dataOut_9_csrInterface_vlmul;
  assign queue_9_deq_bits_csrInterface_vSew = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vSew : queue_dataOut_9_csrInterface_vSew;
  assign queue_9_deq_bits_csrInterface_vxrm = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vxrm : queue_dataOut_9_csrInterface_vxrm;
  assign queue_9_deq_bits_csrInterface_vta = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vta : queue_dataOut_9_csrInterface_vta;
  assign queue_9_deq_bits_csrInterface_vma = _queue_fifo_9_empty ? queue_9_enq_bits_csrInterface_vma : queue_dataOut_9_csrInterface_vma;
  wire         laneVec_9_laneRequest_bits_issueInst = laneRequestSinkWire_9_ready & laneRequestSinkWire_9_valid;
  reg          releasePipe_pipe_v_9;
  wire         releasePipe_pipe_out_9_valid = releasePipe_pipe_v_9;
  wire         laneRequestSourceWire_9_ready;
  wire         validSource_9_valid = laneRequestSourceWire_9_ready & laneRequestSourceWire_9_valid;
  reg  [2:0]   tokenCheck_counter_9;
  wire [2:0]   tokenCheck_counterChange_9 = validSource_9_valid ? 3'h1 : 3'h7;
  assign tokenCheck_9 = ~(tokenCheck_counter_9[2]);
  assign laneRequestSourceWire_9_ready = tokenCheck_9;
  assign queue_9_enq_valid = validSink_9_valid;
  assign queue_9_enq_bits_instructionIndex = validSink_9_bits_instructionIndex;
  assign queue_9_enq_bits_decodeResult_orderReduce = validSink_9_bits_decodeResult_orderReduce;
  assign queue_9_enq_bits_decodeResult_floatMul = validSink_9_bits_decodeResult_floatMul;
  assign queue_9_enq_bits_decodeResult_fpExecutionType = validSink_9_bits_decodeResult_fpExecutionType;
  assign queue_9_enq_bits_decodeResult_float = validSink_9_bits_decodeResult_float;
  assign queue_9_enq_bits_decodeResult_specialSlot = validSink_9_bits_decodeResult_specialSlot;
  assign queue_9_enq_bits_decodeResult_topUop = validSink_9_bits_decodeResult_topUop;
  assign queue_9_enq_bits_decodeResult_popCount = validSink_9_bits_decodeResult_popCount;
  assign queue_9_enq_bits_decodeResult_ffo = validSink_9_bits_decodeResult_ffo;
  assign queue_9_enq_bits_decodeResult_average = validSink_9_bits_decodeResult_average;
  assign queue_9_enq_bits_decodeResult_reverse = validSink_9_bits_decodeResult_reverse;
  assign queue_9_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_9_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_9_enq_bits_decodeResult_scheduler = validSink_9_bits_decodeResult_scheduler;
  assign queue_9_enq_bits_decodeResult_sReadVD = validSink_9_bits_decodeResult_sReadVD;
  assign queue_9_enq_bits_decodeResult_vtype = validSink_9_bits_decodeResult_vtype;
  assign queue_9_enq_bits_decodeResult_sWrite = validSink_9_bits_decodeResult_sWrite;
  assign queue_9_enq_bits_decodeResult_crossRead = validSink_9_bits_decodeResult_crossRead;
  assign queue_9_enq_bits_decodeResult_crossWrite = validSink_9_bits_decodeResult_crossWrite;
  assign queue_9_enq_bits_decodeResult_maskUnit = validSink_9_bits_decodeResult_maskUnit;
  assign queue_9_enq_bits_decodeResult_special = validSink_9_bits_decodeResult_special;
  assign queue_9_enq_bits_decodeResult_saturate = validSink_9_bits_decodeResult_saturate;
  assign queue_9_enq_bits_decodeResult_vwmacc = validSink_9_bits_decodeResult_vwmacc;
  assign queue_9_enq_bits_decodeResult_readOnly = validSink_9_bits_decodeResult_readOnly;
  assign queue_9_enq_bits_decodeResult_maskSource = validSink_9_bits_decodeResult_maskSource;
  assign queue_9_enq_bits_decodeResult_maskDestination = validSink_9_bits_decodeResult_maskDestination;
  assign queue_9_enq_bits_decodeResult_maskLogic = validSink_9_bits_decodeResult_maskLogic;
  assign queue_9_enq_bits_decodeResult_uop = validSink_9_bits_decodeResult_uop;
  assign queue_9_enq_bits_decodeResult_iota = validSink_9_bits_decodeResult_iota;
  assign queue_9_enq_bits_decodeResult_mv = validSink_9_bits_decodeResult_mv;
  assign queue_9_enq_bits_decodeResult_extend = validSink_9_bits_decodeResult_extend;
  assign queue_9_enq_bits_decodeResult_unOrderWrite = validSink_9_bits_decodeResult_unOrderWrite;
  assign queue_9_enq_bits_decodeResult_compress = validSink_9_bits_decodeResult_compress;
  assign queue_9_enq_bits_decodeResult_gather16 = validSink_9_bits_decodeResult_gather16;
  assign queue_9_enq_bits_decodeResult_gather = validSink_9_bits_decodeResult_gather;
  assign queue_9_enq_bits_decodeResult_slid = validSink_9_bits_decodeResult_slid;
  assign queue_9_enq_bits_decodeResult_targetRd = validSink_9_bits_decodeResult_targetRd;
  assign queue_9_enq_bits_decodeResult_widenReduce = validSink_9_bits_decodeResult_widenReduce;
  assign queue_9_enq_bits_decodeResult_red = validSink_9_bits_decodeResult_red;
  assign queue_9_enq_bits_decodeResult_nr = validSink_9_bits_decodeResult_nr;
  assign queue_9_enq_bits_decodeResult_itype = validSink_9_bits_decodeResult_itype;
  assign queue_9_enq_bits_decodeResult_unsigned1 = validSink_9_bits_decodeResult_unsigned1;
  assign queue_9_enq_bits_decodeResult_unsigned0 = validSink_9_bits_decodeResult_unsigned0;
  assign queue_9_enq_bits_decodeResult_other = validSink_9_bits_decodeResult_other;
  assign queue_9_enq_bits_decodeResult_multiCycle = validSink_9_bits_decodeResult_multiCycle;
  assign queue_9_enq_bits_decodeResult_divider = validSink_9_bits_decodeResult_divider;
  assign queue_9_enq_bits_decodeResult_multiplier = validSink_9_bits_decodeResult_multiplier;
  assign queue_9_enq_bits_decodeResult_shift = validSink_9_bits_decodeResult_shift;
  assign queue_9_enq_bits_decodeResult_adder = validSink_9_bits_decodeResult_adder;
  assign queue_9_enq_bits_decodeResult_logic = validSink_9_bits_decodeResult_logic;
  assign queue_9_enq_bits_loadStore = validSink_9_bits_loadStore;
  assign queue_9_enq_bits_issueInst = validSink_9_bits_issueInst;
  assign queue_9_enq_bits_store = validSink_9_bits_store;
  assign queue_9_enq_bits_special = validSink_9_bits_special;
  assign queue_9_enq_bits_lsWholeReg = validSink_9_bits_lsWholeReg;
  assign queue_9_enq_bits_vs1 = validSink_9_bits_vs1;
  assign queue_9_enq_bits_vs2 = validSink_9_bits_vs2;
  assign queue_9_enq_bits_vd = validSink_9_bits_vd;
  assign queue_9_enq_bits_loadStoreEEW = validSink_9_bits_loadStoreEEW;
  assign queue_9_enq_bits_mask = validSink_9_bits_mask;
  assign queue_9_enq_bits_segment = validSink_9_bits_segment;
  assign queue_9_enq_bits_readFromScalar = validSink_9_bits_readFromScalar;
  assign queue_9_enq_bits_csrInterface_vl = validSink_9_bits_csrInterface_vl;
  assign queue_9_enq_bits_csrInterface_vStart = validSink_9_bits_csrInterface_vStart;
  assign queue_9_enq_bits_csrInterface_vlmul = validSink_9_bits_csrInterface_vlmul;
  assign queue_9_enq_bits_csrInterface_vSew = validSink_9_bits_csrInterface_vSew;
  assign queue_9_enq_bits_csrInterface_vxrm = validSink_9_bits_csrInterface_vxrm;
  assign queue_9_enq_bits_csrInterface_vta = validSink_9_bits_csrInterface_vta;
  assign queue_9_enq_bits_csrInterface_vma = validSink_9_bits_csrInterface_vma;
  reg          shifterReg_9_0_valid;
  assign validSink_9_valid = shifterReg_9_0_valid;
  reg  [2:0]   shifterReg_9_0_bits_instructionIndex;
  assign validSink_9_bits_instructionIndex = shifterReg_9_0_bits_instructionIndex;
  reg          shifterReg_9_0_bits_decodeResult_orderReduce;
  assign validSink_9_bits_decodeResult_orderReduce = shifterReg_9_0_bits_decodeResult_orderReduce;
  reg          shifterReg_9_0_bits_decodeResult_floatMul;
  assign validSink_9_bits_decodeResult_floatMul = shifterReg_9_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_9_0_bits_decodeResult_fpExecutionType;
  assign validSink_9_bits_decodeResult_fpExecutionType = shifterReg_9_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_9_0_bits_decodeResult_float;
  assign validSink_9_bits_decodeResult_float = shifterReg_9_0_bits_decodeResult_float;
  reg          shifterReg_9_0_bits_decodeResult_specialSlot;
  assign validSink_9_bits_decodeResult_specialSlot = shifterReg_9_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_9_0_bits_decodeResult_topUop;
  assign validSink_9_bits_decodeResult_topUop = shifterReg_9_0_bits_decodeResult_topUop;
  reg          shifterReg_9_0_bits_decodeResult_popCount;
  assign validSink_9_bits_decodeResult_popCount = shifterReg_9_0_bits_decodeResult_popCount;
  reg          shifterReg_9_0_bits_decodeResult_ffo;
  assign validSink_9_bits_decodeResult_ffo = shifterReg_9_0_bits_decodeResult_ffo;
  reg          shifterReg_9_0_bits_decodeResult_average;
  assign validSink_9_bits_decodeResult_average = shifterReg_9_0_bits_decodeResult_average;
  reg          shifterReg_9_0_bits_decodeResult_reverse;
  assign validSink_9_bits_decodeResult_reverse = shifterReg_9_0_bits_decodeResult_reverse;
  reg          shifterReg_9_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_9_bits_decodeResult_dontNeedExecuteInLane = shifterReg_9_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_9_0_bits_decodeResult_scheduler;
  assign validSink_9_bits_decodeResult_scheduler = shifterReg_9_0_bits_decodeResult_scheduler;
  reg          shifterReg_9_0_bits_decodeResult_sReadVD;
  assign validSink_9_bits_decodeResult_sReadVD = shifterReg_9_0_bits_decodeResult_sReadVD;
  reg          shifterReg_9_0_bits_decodeResult_vtype;
  assign validSink_9_bits_decodeResult_vtype = shifterReg_9_0_bits_decodeResult_vtype;
  reg          shifterReg_9_0_bits_decodeResult_sWrite;
  assign validSink_9_bits_decodeResult_sWrite = shifterReg_9_0_bits_decodeResult_sWrite;
  reg          shifterReg_9_0_bits_decodeResult_crossRead;
  assign validSink_9_bits_decodeResult_crossRead = shifterReg_9_0_bits_decodeResult_crossRead;
  reg          shifterReg_9_0_bits_decodeResult_crossWrite;
  assign validSink_9_bits_decodeResult_crossWrite = shifterReg_9_0_bits_decodeResult_crossWrite;
  reg          shifterReg_9_0_bits_decodeResult_maskUnit;
  assign validSink_9_bits_decodeResult_maskUnit = shifterReg_9_0_bits_decodeResult_maskUnit;
  reg          shifterReg_9_0_bits_decodeResult_special;
  assign validSink_9_bits_decodeResult_special = shifterReg_9_0_bits_decodeResult_special;
  reg          shifterReg_9_0_bits_decodeResult_saturate;
  assign validSink_9_bits_decodeResult_saturate = shifterReg_9_0_bits_decodeResult_saturate;
  reg          shifterReg_9_0_bits_decodeResult_vwmacc;
  assign validSink_9_bits_decodeResult_vwmacc = shifterReg_9_0_bits_decodeResult_vwmacc;
  reg          shifterReg_9_0_bits_decodeResult_readOnly;
  assign validSink_9_bits_decodeResult_readOnly = shifterReg_9_0_bits_decodeResult_readOnly;
  reg          shifterReg_9_0_bits_decodeResult_maskSource;
  assign validSink_9_bits_decodeResult_maskSource = shifterReg_9_0_bits_decodeResult_maskSource;
  reg          shifterReg_9_0_bits_decodeResult_maskDestination;
  assign validSink_9_bits_decodeResult_maskDestination = shifterReg_9_0_bits_decodeResult_maskDestination;
  reg          shifterReg_9_0_bits_decodeResult_maskLogic;
  assign validSink_9_bits_decodeResult_maskLogic = shifterReg_9_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_9_0_bits_decodeResult_uop;
  assign validSink_9_bits_decodeResult_uop = shifterReg_9_0_bits_decodeResult_uop;
  reg          shifterReg_9_0_bits_decodeResult_iota;
  assign validSink_9_bits_decodeResult_iota = shifterReg_9_0_bits_decodeResult_iota;
  reg          shifterReg_9_0_bits_decodeResult_mv;
  assign validSink_9_bits_decodeResult_mv = shifterReg_9_0_bits_decodeResult_mv;
  reg          shifterReg_9_0_bits_decodeResult_extend;
  assign validSink_9_bits_decodeResult_extend = shifterReg_9_0_bits_decodeResult_extend;
  reg          shifterReg_9_0_bits_decodeResult_unOrderWrite;
  assign validSink_9_bits_decodeResult_unOrderWrite = shifterReg_9_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_9_0_bits_decodeResult_compress;
  assign validSink_9_bits_decodeResult_compress = shifterReg_9_0_bits_decodeResult_compress;
  reg          shifterReg_9_0_bits_decodeResult_gather16;
  assign validSink_9_bits_decodeResult_gather16 = shifterReg_9_0_bits_decodeResult_gather16;
  reg          shifterReg_9_0_bits_decodeResult_gather;
  assign validSink_9_bits_decodeResult_gather = shifterReg_9_0_bits_decodeResult_gather;
  reg          shifterReg_9_0_bits_decodeResult_slid;
  assign validSink_9_bits_decodeResult_slid = shifterReg_9_0_bits_decodeResult_slid;
  reg          shifterReg_9_0_bits_decodeResult_targetRd;
  assign validSink_9_bits_decodeResult_targetRd = shifterReg_9_0_bits_decodeResult_targetRd;
  reg          shifterReg_9_0_bits_decodeResult_widenReduce;
  assign validSink_9_bits_decodeResult_widenReduce = shifterReg_9_0_bits_decodeResult_widenReduce;
  reg          shifterReg_9_0_bits_decodeResult_red;
  assign validSink_9_bits_decodeResult_red = shifterReg_9_0_bits_decodeResult_red;
  reg          shifterReg_9_0_bits_decodeResult_nr;
  assign validSink_9_bits_decodeResult_nr = shifterReg_9_0_bits_decodeResult_nr;
  reg          shifterReg_9_0_bits_decodeResult_itype;
  assign validSink_9_bits_decodeResult_itype = shifterReg_9_0_bits_decodeResult_itype;
  reg          shifterReg_9_0_bits_decodeResult_unsigned1;
  assign validSink_9_bits_decodeResult_unsigned1 = shifterReg_9_0_bits_decodeResult_unsigned1;
  reg          shifterReg_9_0_bits_decodeResult_unsigned0;
  assign validSink_9_bits_decodeResult_unsigned0 = shifterReg_9_0_bits_decodeResult_unsigned0;
  reg          shifterReg_9_0_bits_decodeResult_other;
  assign validSink_9_bits_decodeResult_other = shifterReg_9_0_bits_decodeResult_other;
  reg          shifterReg_9_0_bits_decodeResult_multiCycle;
  assign validSink_9_bits_decodeResult_multiCycle = shifterReg_9_0_bits_decodeResult_multiCycle;
  reg          shifterReg_9_0_bits_decodeResult_divider;
  assign validSink_9_bits_decodeResult_divider = shifterReg_9_0_bits_decodeResult_divider;
  reg          shifterReg_9_0_bits_decodeResult_multiplier;
  assign validSink_9_bits_decodeResult_multiplier = shifterReg_9_0_bits_decodeResult_multiplier;
  reg          shifterReg_9_0_bits_decodeResult_shift;
  assign validSink_9_bits_decodeResult_shift = shifterReg_9_0_bits_decodeResult_shift;
  reg          shifterReg_9_0_bits_decodeResult_adder;
  assign validSink_9_bits_decodeResult_adder = shifterReg_9_0_bits_decodeResult_adder;
  reg          shifterReg_9_0_bits_decodeResult_logic;
  assign validSink_9_bits_decodeResult_logic = shifterReg_9_0_bits_decodeResult_logic;
  reg          shifterReg_9_0_bits_loadStore;
  assign validSink_9_bits_loadStore = shifterReg_9_0_bits_loadStore;
  reg          shifterReg_9_0_bits_issueInst;
  assign validSink_9_bits_issueInst = shifterReg_9_0_bits_issueInst;
  reg          shifterReg_9_0_bits_store;
  assign validSink_9_bits_store = shifterReg_9_0_bits_store;
  reg          shifterReg_9_0_bits_special;
  assign validSink_9_bits_special = shifterReg_9_0_bits_special;
  reg          shifterReg_9_0_bits_lsWholeReg;
  assign validSink_9_bits_lsWholeReg = shifterReg_9_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_9_0_bits_vs1;
  assign validSink_9_bits_vs1 = shifterReg_9_0_bits_vs1;
  reg  [4:0]   shifterReg_9_0_bits_vs2;
  assign validSink_9_bits_vs2 = shifterReg_9_0_bits_vs2;
  reg  [4:0]   shifterReg_9_0_bits_vd;
  assign validSink_9_bits_vd = shifterReg_9_0_bits_vd;
  reg  [1:0]   shifterReg_9_0_bits_loadStoreEEW;
  assign validSink_9_bits_loadStoreEEW = shifterReg_9_0_bits_loadStoreEEW;
  reg          shifterReg_9_0_bits_mask;
  assign validSink_9_bits_mask = shifterReg_9_0_bits_mask;
  reg  [2:0]   shifterReg_9_0_bits_segment;
  assign validSink_9_bits_segment = shifterReg_9_0_bits_segment;
  reg  [31:0]  shifterReg_9_0_bits_readFromScalar;
  assign validSink_9_bits_readFromScalar = shifterReg_9_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_9_0_bits_csrInterface_vl;
  assign validSink_9_bits_csrInterface_vl = shifterReg_9_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_9_0_bits_csrInterface_vStart;
  assign validSink_9_bits_csrInterface_vStart = shifterReg_9_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_9_0_bits_csrInterface_vlmul;
  assign validSink_9_bits_csrInterface_vlmul = shifterReg_9_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_9_0_bits_csrInterface_vSew;
  assign validSink_9_bits_csrInterface_vSew = shifterReg_9_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_9_0_bits_csrInterface_vxrm;
  assign validSink_9_bits_csrInterface_vxrm = shifterReg_9_0_bits_csrInterface_vxrm;
  reg          shifterReg_9_0_bits_csrInterface_vta;
  assign validSink_9_bits_csrInterface_vta = shifterReg_9_0_bits_csrInterface_vta;
  reg          shifterReg_9_0_bits_csrInterface_vma;
  assign validSink_9_bits_csrInterface_vma = shifterReg_9_0_bits_csrInterface_vma;
  wire         shifterValid_9 = shifterReg_9_0_valid | validSource_9_valid;
  wire         validSink_10_valid;
  wire [2:0]   validSink_10_bits_instructionIndex;
  wire         validSink_10_bits_decodeResult_orderReduce;
  wire         validSink_10_bits_decodeResult_floatMul;
  wire [1:0]   validSink_10_bits_decodeResult_fpExecutionType;
  wire         validSink_10_bits_decodeResult_float;
  wire         validSink_10_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_10_bits_decodeResult_topUop;
  wire         validSink_10_bits_decodeResult_popCount;
  wire         validSink_10_bits_decodeResult_ffo;
  wire         validSink_10_bits_decodeResult_average;
  wire         validSink_10_bits_decodeResult_reverse;
  wire         validSink_10_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_10_bits_decodeResult_scheduler;
  wire         validSink_10_bits_decodeResult_sReadVD;
  wire         validSink_10_bits_decodeResult_vtype;
  wire         validSink_10_bits_decodeResult_sWrite;
  wire         validSink_10_bits_decodeResult_crossRead;
  wire         validSink_10_bits_decodeResult_crossWrite;
  wire         validSink_10_bits_decodeResult_maskUnit;
  wire         validSink_10_bits_decodeResult_special;
  wire         validSink_10_bits_decodeResult_saturate;
  wire         validSink_10_bits_decodeResult_vwmacc;
  wire         validSink_10_bits_decodeResult_readOnly;
  wire         validSink_10_bits_decodeResult_maskSource;
  wire         validSink_10_bits_decodeResult_maskDestination;
  wire         validSink_10_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_10_bits_decodeResult_uop;
  wire         validSink_10_bits_decodeResult_iota;
  wire         validSink_10_bits_decodeResult_mv;
  wire         validSink_10_bits_decodeResult_extend;
  wire         validSink_10_bits_decodeResult_unOrderWrite;
  wire         validSink_10_bits_decodeResult_compress;
  wire         validSink_10_bits_decodeResult_gather16;
  wire         validSink_10_bits_decodeResult_gather;
  wire         validSink_10_bits_decodeResult_slid;
  wire         validSink_10_bits_decodeResult_targetRd;
  wire         validSink_10_bits_decodeResult_widenReduce;
  wire         validSink_10_bits_decodeResult_red;
  wire         validSink_10_bits_decodeResult_nr;
  wire         validSink_10_bits_decodeResult_itype;
  wire         validSink_10_bits_decodeResult_unsigned1;
  wire         validSink_10_bits_decodeResult_unsigned0;
  wire         validSink_10_bits_decodeResult_other;
  wire         validSink_10_bits_decodeResult_multiCycle;
  wire         validSink_10_bits_decodeResult_divider;
  wire         validSink_10_bits_decodeResult_multiplier;
  wire         validSink_10_bits_decodeResult_shift;
  wire         validSink_10_bits_decodeResult_adder;
  wire         validSink_10_bits_decodeResult_logic;
  wire         validSink_10_bits_loadStore;
  wire         validSink_10_bits_issueInst;
  wire         validSink_10_bits_store;
  wire         validSink_10_bits_special;
  wire         validSink_10_bits_lsWholeReg;
  wire [4:0]   validSink_10_bits_vs1;
  wire [4:0]   validSink_10_bits_vs2;
  wire [4:0]   validSink_10_bits_vd;
  wire [1:0]   validSink_10_bits_loadStoreEEW;
  wire         validSink_10_bits_mask;
  wire [2:0]   validSink_10_bits_segment;
  wire [31:0]  validSink_10_bits_readFromScalar;
  wire [11:0]  validSink_10_bits_csrInterface_vl;
  wire [11:0]  validSink_10_bits_csrInterface_vStart;
  wire [2:0]   validSink_10_bits_csrInterface_vlmul;
  wire [1:0]   validSink_10_bits_csrInterface_vSew;
  wire [1:0]   validSink_10_bits_csrInterface_vxrm;
  wire         validSink_10_bits_csrInterface_vta;
  wire         validSink_10_bits_csrInterface_vma;
  wire         laneRequestSinkWire_10_valid = queue_10_deq_valid;
  wire [2:0]   laneRequestSinkWire_10_bits_instructionIndex = queue_10_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_10_bits_decodeResult_orderReduce = queue_10_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_10_bits_decodeResult_floatMul = queue_10_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_10_bits_decodeResult_fpExecutionType = queue_10_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_10_bits_decodeResult_float = queue_10_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_10_bits_decodeResult_specialSlot = queue_10_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_10_bits_decodeResult_topUop = queue_10_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_10_bits_decodeResult_popCount = queue_10_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_10_bits_decodeResult_ffo = queue_10_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_10_bits_decodeResult_average = queue_10_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_10_bits_decodeResult_reverse = queue_10_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_10_bits_decodeResult_dontNeedExecuteInLane = queue_10_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_10_bits_decodeResult_scheduler = queue_10_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_10_bits_decodeResult_sReadVD = queue_10_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_10_bits_decodeResult_vtype = queue_10_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_10_bits_decodeResult_sWrite = queue_10_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_10_bits_decodeResult_crossRead = queue_10_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_10_bits_decodeResult_crossWrite = queue_10_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_10_bits_decodeResult_maskUnit = queue_10_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_10_bits_decodeResult_special = queue_10_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_10_bits_decodeResult_saturate = queue_10_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_10_bits_decodeResult_vwmacc = queue_10_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_10_bits_decodeResult_readOnly = queue_10_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_10_bits_decodeResult_maskSource = queue_10_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_10_bits_decodeResult_maskDestination = queue_10_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_10_bits_decodeResult_maskLogic = queue_10_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_10_bits_decodeResult_uop = queue_10_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_10_bits_decodeResult_iota = queue_10_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_10_bits_decodeResult_mv = queue_10_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_10_bits_decodeResult_extend = queue_10_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_10_bits_decodeResult_unOrderWrite = queue_10_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_10_bits_decodeResult_compress = queue_10_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_10_bits_decodeResult_gather16 = queue_10_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_10_bits_decodeResult_gather = queue_10_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_10_bits_decodeResult_slid = queue_10_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_10_bits_decodeResult_targetRd = queue_10_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_10_bits_decodeResult_widenReduce = queue_10_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_10_bits_decodeResult_red = queue_10_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_10_bits_decodeResult_nr = queue_10_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_10_bits_decodeResult_itype = queue_10_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_10_bits_decodeResult_unsigned1 = queue_10_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_10_bits_decodeResult_unsigned0 = queue_10_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_10_bits_decodeResult_other = queue_10_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_10_bits_decodeResult_multiCycle = queue_10_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_10_bits_decodeResult_divider = queue_10_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_10_bits_decodeResult_multiplier = queue_10_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_10_bits_decodeResult_shift = queue_10_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_10_bits_decodeResult_adder = queue_10_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_10_bits_decodeResult_logic = queue_10_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_10_bits_loadStore = queue_10_deq_bits_loadStore;
  wire         laneRequestSinkWire_10_bits_issueInst = queue_10_deq_bits_issueInst;
  wire         laneRequestSinkWire_10_bits_store = queue_10_deq_bits_store;
  wire         laneRequestSinkWire_10_bits_special = queue_10_deq_bits_special;
  wire         laneRequestSinkWire_10_bits_lsWholeReg = queue_10_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_10_bits_vs1 = queue_10_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_10_bits_vs2 = queue_10_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_10_bits_vd = queue_10_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_10_bits_loadStoreEEW = queue_10_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_10_bits_mask = queue_10_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_10_bits_segment = queue_10_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_10_bits_readFromScalar = queue_10_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_10_bits_csrInterface_vl = queue_10_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_10_bits_csrInterface_vStart = queue_10_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_10_bits_csrInterface_vlmul = queue_10_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_10_bits_csrInterface_vSew = queue_10_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_10_bits_csrInterface_vxrm = queue_10_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_10_bits_csrInterface_vta = queue_10_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_10_bits_csrInterface_vma = queue_10_deq_bits_csrInterface_vma;
  wire [1:0]   queue_10_enq_bits_csrInterface_vxrm;
  wire         queue_10_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_30 = {queue_10_enq_bits_csrInterface_vxrm, queue_10_enq_bits_csrInterface_vta};
  wire         queue_10_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_30 = {queue_dataIn_lo_hi_30, queue_10_enq_bits_csrInterface_vma};
  wire [2:0]   queue_10_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_10_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_30 = {queue_10_enq_bits_csrInterface_vlmul, queue_10_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_10_enq_bits_csrInterface_vl;
  wire [11:0]  queue_10_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_30 = {queue_10_enq_bits_csrInterface_vl, queue_10_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_30 = {queue_dataIn_hi_hi_30, queue_dataIn_hi_lo_30};
  wire         queue_10_enq_bits_decodeResult_shift;
  wire         queue_10_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_10 = {queue_10_enq_bits_decodeResult_shift, queue_10_enq_bits_decodeResult_adder};
  wire         queue_10_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_10 = {queue_dataIn_lo_lo_lo_lo_hi_10, queue_10_enq_bits_decodeResult_logic};
  wire         queue_10_enq_bits_decodeResult_multiCycle;
  wire         queue_10_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_10 = {queue_10_enq_bits_decodeResult_multiCycle, queue_10_enq_bits_decodeResult_divider};
  wire         queue_10_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_10 = {queue_dataIn_lo_lo_lo_hi_hi_10, queue_10_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_10 = {queue_dataIn_lo_lo_lo_hi_10, queue_dataIn_lo_lo_lo_lo_10};
  wire         queue_10_enq_bits_decodeResult_unsigned1;
  wire         queue_10_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_10 = {queue_10_enq_bits_decodeResult_unsigned1, queue_10_enq_bits_decodeResult_unsigned0};
  wire         queue_10_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_10 = {queue_dataIn_lo_lo_hi_lo_hi_10, queue_10_enq_bits_decodeResult_other};
  wire         queue_10_enq_bits_decodeResult_red;
  wire         queue_10_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_10 = {queue_10_enq_bits_decodeResult_red, queue_10_enq_bits_decodeResult_nr};
  wire         queue_10_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_10 = {queue_dataIn_lo_lo_hi_hi_hi_10, queue_10_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_20 = {queue_dataIn_lo_lo_hi_hi_10, queue_dataIn_lo_lo_hi_lo_10};
  wire [11:0]  queue_dataIn_lo_lo_20 = {queue_dataIn_lo_lo_hi_20, queue_dataIn_lo_lo_lo_10};
  wire         queue_10_enq_bits_decodeResult_slid;
  wire         queue_10_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_10 = {queue_10_enq_bits_decodeResult_slid, queue_10_enq_bits_decodeResult_targetRd};
  wire         queue_10_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_10 = {queue_dataIn_lo_hi_lo_lo_hi_10, queue_10_enq_bits_decodeResult_widenReduce};
  wire         queue_10_enq_bits_decodeResult_compress;
  wire         queue_10_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_10 = {queue_10_enq_bits_decodeResult_compress, queue_10_enq_bits_decodeResult_gather16};
  wire         queue_10_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_10 = {queue_dataIn_lo_hi_lo_hi_hi_10, queue_10_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_20 = {queue_dataIn_lo_hi_lo_hi_10, queue_dataIn_lo_hi_lo_lo_10};
  wire         queue_10_enq_bits_decodeResult_mv;
  wire         queue_10_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_10 = {queue_10_enq_bits_decodeResult_mv, queue_10_enq_bits_decodeResult_extend};
  wire         queue_10_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_10 = {queue_dataIn_lo_hi_hi_lo_hi_10, queue_10_enq_bits_decodeResult_unOrderWrite};
  wire         queue_10_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_10_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_10 = {queue_10_enq_bits_decodeResult_maskLogic, queue_10_enq_bits_decodeResult_uop};
  wire         queue_10_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_10 = {queue_dataIn_lo_hi_hi_hi_hi_10, queue_10_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_20 = {queue_dataIn_lo_hi_hi_hi_10, queue_dataIn_lo_hi_hi_lo_10};
  wire [14:0]  queue_dataIn_lo_hi_31 = {queue_dataIn_lo_hi_hi_20, queue_dataIn_lo_hi_lo_20};
  wire [26:0]  queue_dataIn_lo_31 = {queue_dataIn_lo_hi_31, queue_dataIn_lo_lo_20};
  wire         queue_10_enq_bits_decodeResult_readOnly;
  wire         queue_10_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_10 = {queue_10_enq_bits_decodeResult_readOnly, queue_10_enq_bits_decodeResult_maskSource};
  wire         queue_10_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_10 = {queue_dataIn_hi_lo_lo_lo_hi_10, queue_10_enq_bits_decodeResult_maskDestination};
  wire         queue_10_enq_bits_decodeResult_special;
  wire         queue_10_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_10 = {queue_10_enq_bits_decodeResult_special, queue_10_enq_bits_decodeResult_saturate};
  wire         queue_10_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_10 = {queue_dataIn_hi_lo_lo_hi_hi_10, queue_10_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_20 = {queue_dataIn_hi_lo_lo_hi_10, queue_dataIn_hi_lo_lo_lo_10};
  wire         queue_10_enq_bits_decodeResult_crossRead;
  wire         queue_10_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_10 = {queue_10_enq_bits_decodeResult_crossRead, queue_10_enq_bits_decodeResult_crossWrite};
  wire         queue_10_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_10 = {queue_dataIn_hi_lo_hi_lo_hi_10, queue_10_enq_bits_decodeResult_maskUnit};
  wire         queue_10_enq_bits_decodeResult_sReadVD;
  wire         queue_10_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_10 = {queue_10_enq_bits_decodeResult_sReadVD, queue_10_enq_bits_decodeResult_vtype};
  wire         queue_10_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_10 = {queue_dataIn_hi_lo_hi_hi_hi_10, queue_10_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_20 = {queue_dataIn_hi_lo_hi_hi_10, queue_dataIn_hi_lo_hi_lo_10};
  wire [11:0]  queue_dataIn_hi_lo_31 = {queue_dataIn_hi_lo_hi_20, queue_dataIn_hi_lo_lo_20};
  wire         queue_10_enq_bits_decodeResult_reverse;
  wire         queue_10_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_10 = {queue_10_enq_bits_decodeResult_reverse, queue_10_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_10_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_10 = {queue_dataIn_hi_hi_lo_lo_hi_10, queue_10_enq_bits_decodeResult_scheduler};
  wire         queue_10_enq_bits_decodeResult_popCount;
  wire         queue_10_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_10 = {queue_10_enq_bits_decodeResult_popCount, queue_10_enq_bits_decodeResult_ffo};
  wire         queue_10_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_10 = {queue_dataIn_hi_hi_lo_hi_hi_10, queue_10_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_20 = {queue_dataIn_hi_hi_lo_hi_10, queue_dataIn_hi_hi_lo_lo_10};
  wire         queue_10_enq_bits_decodeResult_float;
  wire         queue_10_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_10 = {queue_10_enq_bits_decodeResult_float, queue_10_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_10_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_10 = {queue_dataIn_hi_hi_hi_lo_hi_10, queue_10_enq_bits_decodeResult_topUop};
  wire         queue_10_enq_bits_decodeResult_orderReduce;
  wire         queue_10_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_10 = {queue_10_enq_bits_decodeResult_orderReduce, queue_10_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_10_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_10 = {queue_dataIn_hi_hi_hi_hi_hi_10, queue_10_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_20 = {queue_dataIn_hi_hi_hi_hi_10, queue_dataIn_hi_hi_hi_lo_10};
  wire [16:0]  queue_dataIn_hi_hi_31 = {queue_dataIn_hi_hi_hi_20, queue_dataIn_hi_hi_lo_20};
  wire [28:0]  queue_dataIn_hi_31 = {queue_dataIn_hi_hi_31, queue_dataIn_hi_lo_31};
  wire [2:0]   queue_10_enq_bits_segment;
  wire [31:0]  queue_10_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_21 = {queue_10_enq_bits_segment, queue_10_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_21 = {queue_dataIn_lo_lo_hi_21, queue_dataIn_hi_30, queue_dataIn_lo_30};
  wire [1:0]   queue_10_enq_bits_loadStoreEEW;
  wire         queue_10_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_21 = {queue_10_enq_bits_loadStoreEEW, queue_10_enq_bits_mask};
  wire [4:0]   queue_10_enq_bits_vs2;
  wire [4:0]   queue_10_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_21 = {queue_10_enq_bits_vs2, queue_10_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_32 = {queue_dataIn_lo_hi_hi_21, queue_dataIn_lo_hi_lo_21};
  wire [80:0]  queue_dataIn_lo_32 = {queue_dataIn_lo_hi_32, queue_dataIn_lo_lo_21};
  wire         queue_10_enq_bits_lsWholeReg;
  wire [4:0]   queue_10_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_21 = {queue_10_enq_bits_lsWholeReg, queue_10_enq_bits_vs1};
  wire         queue_10_enq_bits_store;
  wire         queue_10_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_21 = {queue_10_enq_bits_store, queue_10_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_32 = {queue_dataIn_hi_lo_hi_21, queue_dataIn_hi_lo_lo_21};
  wire         queue_10_enq_bits_loadStore;
  wire         queue_10_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_21 = {queue_10_enq_bits_loadStore, queue_10_enq_bits_issueInst};
  wire [2:0]   queue_10_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_21 = {queue_10_enq_bits_instructionIndex, queue_dataIn_hi_31, queue_dataIn_lo_31};
  wire [60:0]  queue_dataIn_hi_hi_32 = {queue_dataIn_hi_hi_hi_21, queue_dataIn_hi_hi_lo_21};
  wire [68:0]  queue_dataIn_hi_32 = {queue_dataIn_hi_hi_32, queue_dataIn_hi_lo_32};
  wire [149:0] queue_dataIn_10 = {queue_dataIn_hi_32, queue_dataIn_lo_32};
  wire         queue_dataOut_10_csrInterface_vma = _queue_fifo_10_data_out[0];
  wire         queue_dataOut_10_csrInterface_vta = _queue_fifo_10_data_out[1];
  wire [1:0]   queue_dataOut_10_csrInterface_vxrm = _queue_fifo_10_data_out[3:2];
  wire [1:0]   queue_dataOut_10_csrInterface_vSew = _queue_fifo_10_data_out[5:4];
  wire [2:0]   queue_dataOut_10_csrInterface_vlmul = _queue_fifo_10_data_out[8:6];
  wire [11:0]  queue_dataOut_10_csrInterface_vStart = _queue_fifo_10_data_out[20:9];
  wire [11:0]  queue_dataOut_10_csrInterface_vl = _queue_fifo_10_data_out[32:21];
  wire [31:0]  queue_dataOut_10_readFromScalar = _queue_fifo_10_data_out[64:33];
  wire [2:0]   queue_dataOut_10_segment = _queue_fifo_10_data_out[67:65];
  wire         queue_dataOut_10_mask = _queue_fifo_10_data_out[68];
  wire [1:0]   queue_dataOut_10_loadStoreEEW = _queue_fifo_10_data_out[70:69];
  wire [4:0]   queue_dataOut_10_vd = _queue_fifo_10_data_out[75:71];
  wire [4:0]   queue_dataOut_10_vs2 = _queue_fifo_10_data_out[80:76];
  wire [4:0]   queue_dataOut_10_vs1 = _queue_fifo_10_data_out[85:81];
  wire         queue_dataOut_10_lsWholeReg = _queue_fifo_10_data_out[86];
  wire         queue_dataOut_10_special = _queue_fifo_10_data_out[87];
  wire         queue_dataOut_10_store = _queue_fifo_10_data_out[88];
  wire         queue_dataOut_10_issueInst = _queue_fifo_10_data_out[89];
  wire         queue_dataOut_10_loadStore = _queue_fifo_10_data_out[90];
  wire         queue_dataOut_10_decodeResult_logic = _queue_fifo_10_data_out[91];
  wire         queue_dataOut_10_decodeResult_adder = _queue_fifo_10_data_out[92];
  wire         queue_dataOut_10_decodeResult_shift = _queue_fifo_10_data_out[93];
  wire         queue_dataOut_10_decodeResult_multiplier = _queue_fifo_10_data_out[94];
  wire         queue_dataOut_10_decodeResult_divider = _queue_fifo_10_data_out[95];
  wire         queue_dataOut_10_decodeResult_multiCycle = _queue_fifo_10_data_out[96];
  wire         queue_dataOut_10_decodeResult_other = _queue_fifo_10_data_out[97];
  wire         queue_dataOut_10_decodeResult_unsigned0 = _queue_fifo_10_data_out[98];
  wire         queue_dataOut_10_decodeResult_unsigned1 = _queue_fifo_10_data_out[99];
  wire         queue_dataOut_10_decodeResult_itype = _queue_fifo_10_data_out[100];
  wire         queue_dataOut_10_decodeResult_nr = _queue_fifo_10_data_out[101];
  wire         queue_dataOut_10_decodeResult_red = _queue_fifo_10_data_out[102];
  wire         queue_dataOut_10_decodeResult_widenReduce = _queue_fifo_10_data_out[103];
  wire         queue_dataOut_10_decodeResult_targetRd = _queue_fifo_10_data_out[104];
  wire         queue_dataOut_10_decodeResult_slid = _queue_fifo_10_data_out[105];
  wire         queue_dataOut_10_decodeResult_gather = _queue_fifo_10_data_out[106];
  wire         queue_dataOut_10_decodeResult_gather16 = _queue_fifo_10_data_out[107];
  wire         queue_dataOut_10_decodeResult_compress = _queue_fifo_10_data_out[108];
  wire         queue_dataOut_10_decodeResult_unOrderWrite = _queue_fifo_10_data_out[109];
  wire         queue_dataOut_10_decodeResult_extend = _queue_fifo_10_data_out[110];
  wire         queue_dataOut_10_decodeResult_mv = _queue_fifo_10_data_out[111];
  wire         queue_dataOut_10_decodeResult_iota = _queue_fifo_10_data_out[112];
  wire [3:0]   queue_dataOut_10_decodeResult_uop = _queue_fifo_10_data_out[116:113];
  wire         queue_dataOut_10_decodeResult_maskLogic = _queue_fifo_10_data_out[117];
  wire         queue_dataOut_10_decodeResult_maskDestination = _queue_fifo_10_data_out[118];
  wire         queue_dataOut_10_decodeResult_maskSource = _queue_fifo_10_data_out[119];
  wire         queue_dataOut_10_decodeResult_readOnly = _queue_fifo_10_data_out[120];
  wire         queue_dataOut_10_decodeResult_vwmacc = _queue_fifo_10_data_out[121];
  wire         queue_dataOut_10_decodeResult_saturate = _queue_fifo_10_data_out[122];
  wire         queue_dataOut_10_decodeResult_special = _queue_fifo_10_data_out[123];
  wire         queue_dataOut_10_decodeResult_maskUnit = _queue_fifo_10_data_out[124];
  wire         queue_dataOut_10_decodeResult_crossWrite = _queue_fifo_10_data_out[125];
  wire         queue_dataOut_10_decodeResult_crossRead = _queue_fifo_10_data_out[126];
  wire         queue_dataOut_10_decodeResult_sWrite = _queue_fifo_10_data_out[127];
  wire         queue_dataOut_10_decodeResult_vtype = _queue_fifo_10_data_out[128];
  wire         queue_dataOut_10_decodeResult_sReadVD = _queue_fifo_10_data_out[129];
  wire         queue_dataOut_10_decodeResult_scheduler = _queue_fifo_10_data_out[130];
  wire         queue_dataOut_10_decodeResult_dontNeedExecuteInLane = _queue_fifo_10_data_out[131];
  wire         queue_dataOut_10_decodeResult_reverse = _queue_fifo_10_data_out[132];
  wire         queue_dataOut_10_decodeResult_average = _queue_fifo_10_data_out[133];
  wire         queue_dataOut_10_decodeResult_ffo = _queue_fifo_10_data_out[134];
  wire         queue_dataOut_10_decodeResult_popCount = _queue_fifo_10_data_out[135];
  wire [4:0]   queue_dataOut_10_decodeResult_topUop = _queue_fifo_10_data_out[140:136];
  wire         queue_dataOut_10_decodeResult_specialSlot = _queue_fifo_10_data_out[141];
  wire         queue_dataOut_10_decodeResult_float = _queue_fifo_10_data_out[142];
  wire [1:0]   queue_dataOut_10_decodeResult_fpExecutionType = _queue_fifo_10_data_out[144:143];
  wire         queue_dataOut_10_decodeResult_floatMul = _queue_fifo_10_data_out[145];
  wire         queue_dataOut_10_decodeResult_orderReduce = _queue_fifo_10_data_out[146];
  wire [2:0]   queue_dataOut_10_instructionIndex = _queue_fifo_10_data_out[149:147];
  wire         queue_10_enq_ready = ~_queue_fifo_10_full;
  wire         queue_10_enq_valid;
  assign queue_10_deq_valid = ~_queue_fifo_10_empty | queue_10_enq_valid;
  assign queue_10_deq_bits_instructionIndex = _queue_fifo_10_empty ? queue_10_enq_bits_instructionIndex : queue_dataOut_10_instructionIndex;
  assign queue_10_deq_bits_decodeResult_orderReduce = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_orderReduce : queue_dataOut_10_decodeResult_orderReduce;
  assign queue_10_deq_bits_decodeResult_floatMul = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_floatMul : queue_dataOut_10_decodeResult_floatMul;
  assign queue_10_deq_bits_decodeResult_fpExecutionType = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_fpExecutionType : queue_dataOut_10_decodeResult_fpExecutionType;
  assign queue_10_deq_bits_decodeResult_float = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_float : queue_dataOut_10_decodeResult_float;
  assign queue_10_deq_bits_decodeResult_specialSlot = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_specialSlot : queue_dataOut_10_decodeResult_specialSlot;
  assign queue_10_deq_bits_decodeResult_topUop = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_topUop : queue_dataOut_10_decodeResult_topUop;
  assign queue_10_deq_bits_decodeResult_popCount = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_popCount : queue_dataOut_10_decodeResult_popCount;
  assign queue_10_deq_bits_decodeResult_ffo = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_ffo : queue_dataOut_10_decodeResult_ffo;
  assign queue_10_deq_bits_decodeResult_average = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_average : queue_dataOut_10_decodeResult_average;
  assign queue_10_deq_bits_decodeResult_reverse = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_reverse : queue_dataOut_10_decodeResult_reverse;
  assign queue_10_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_10_decodeResult_dontNeedExecuteInLane;
  assign queue_10_deq_bits_decodeResult_scheduler = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_scheduler : queue_dataOut_10_decodeResult_scheduler;
  assign queue_10_deq_bits_decodeResult_sReadVD = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_sReadVD : queue_dataOut_10_decodeResult_sReadVD;
  assign queue_10_deq_bits_decodeResult_vtype = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_vtype : queue_dataOut_10_decodeResult_vtype;
  assign queue_10_deq_bits_decodeResult_sWrite = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_sWrite : queue_dataOut_10_decodeResult_sWrite;
  assign queue_10_deq_bits_decodeResult_crossRead = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_crossRead : queue_dataOut_10_decodeResult_crossRead;
  assign queue_10_deq_bits_decodeResult_crossWrite = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_crossWrite : queue_dataOut_10_decodeResult_crossWrite;
  assign queue_10_deq_bits_decodeResult_maskUnit = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_maskUnit : queue_dataOut_10_decodeResult_maskUnit;
  assign queue_10_deq_bits_decodeResult_special = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_special : queue_dataOut_10_decodeResult_special;
  assign queue_10_deq_bits_decodeResult_saturate = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_saturate : queue_dataOut_10_decodeResult_saturate;
  assign queue_10_deq_bits_decodeResult_vwmacc = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_vwmacc : queue_dataOut_10_decodeResult_vwmacc;
  assign queue_10_deq_bits_decodeResult_readOnly = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_readOnly : queue_dataOut_10_decodeResult_readOnly;
  assign queue_10_deq_bits_decodeResult_maskSource = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_maskSource : queue_dataOut_10_decodeResult_maskSource;
  assign queue_10_deq_bits_decodeResult_maskDestination = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_maskDestination : queue_dataOut_10_decodeResult_maskDestination;
  assign queue_10_deq_bits_decodeResult_maskLogic = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_maskLogic : queue_dataOut_10_decodeResult_maskLogic;
  assign queue_10_deq_bits_decodeResult_uop = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_uop : queue_dataOut_10_decodeResult_uop;
  assign queue_10_deq_bits_decodeResult_iota = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_iota : queue_dataOut_10_decodeResult_iota;
  assign queue_10_deq_bits_decodeResult_mv = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_mv : queue_dataOut_10_decodeResult_mv;
  assign queue_10_deq_bits_decodeResult_extend = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_extend : queue_dataOut_10_decodeResult_extend;
  assign queue_10_deq_bits_decodeResult_unOrderWrite = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_unOrderWrite : queue_dataOut_10_decodeResult_unOrderWrite;
  assign queue_10_deq_bits_decodeResult_compress = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_compress : queue_dataOut_10_decodeResult_compress;
  assign queue_10_deq_bits_decodeResult_gather16 = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_gather16 : queue_dataOut_10_decodeResult_gather16;
  assign queue_10_deq_bits_decodeResult_gather = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_gather : queue_dataOut_10_decodeResult_gather;
  assign queue_10_deq_bits_decodeResult_slid = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_slid : queue_dataOut_10_decodeResult_slid;
  assign queue_10_deq_bits_decodeResult_targetRd = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_targetRd : queue_dataOut_10_decodeResult_targetRd;
  assign queue_10_deq_bits_decodeResult_widenReduce = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_widenReduce : queue_dataOut_10_decodeResult_widenReduce;
  assign queue_10_deq_bits_decodeResult_red = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_red : queue_dataOut_10_decodeResult_red;
  assign queue_10_deq_bits_decodeResult_nr = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_nr : queue_dataOut_10_decodeResult_nr;
  assign queue_10_deq_bits_decodeResult_itype = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_itype : queue_dataOut_10_decodeResult_itype;
  assign queue_10_deq_bits_decodeResult_unsigned1 = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_unsigned1 : queue_dataOut_10_decodeResult_unsigned1;
  assign queue_10_deq_bits_decodeResult_unsigned0 = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_unsigned0 : queue_dataOut_10_decodeResult_unsigned0;
  assign queue_10_deq_bits_decodeResult_other = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_other : queue_dataOut_10_decodeResult_other;
  assign queue_10_deq_bits_decodeResult_multiCycle = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_multiCycle : queue_dataOut_10_decodeResult_multiCycle;
  assign queue_10_deq_bits_decodeResult_divider = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_divider : queue_dataOut_10_decodeResult_divider;
  assign queue_10_deq_bits_decodeResult_multiplier = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_multiplier : queue_dataOut_10_decodeResult_multiplier;
  assign queue_10_deq_bits_decodeResult_shift = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_shift : queue_dataOut_10_decodeResult_shift;
  assign queue_10_deq_bits_decodeResult_adder = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_adder : queue_dataOut_10_decodeResult_adder;
  assign queue_10_deq_bits_decodeResult_logic = _queue_fifo_10_empty ? queue_10_enq_bits_decodeResult_logic : queue_dataOut_10_decodeResult_logic;
  assign queue_10_deq_bits_loadStore = _queue_fifo_10_empty ? queue_10_enq_bits_loadStore : queue_dataOut_10_loadStore;
  assign queue_10_deq_bits_issueInst = _queue_fifo_10_empty ? queue_10_enq_bits_issueInst : queue_dataOut_10_issueInst;
  assign queue_10_deq_bits_store = _queue_fifo_10_empty ? queue_10_enq_bits_store : queue_dataOut_10_store;
  assign queue_10_deq_bits_special = _queue_fifo_10_empty ? queue_10_enq_bits_special : queue_dataOut_10_special;
  assign queue_10_deq_bits_lsWholeReg = _queue_fifo_10_empty ? queue_10_enq_bits_lsWholeReg : queue_dataOut_10_lsWholeReg;
  assign queue_10_deq_bits_vs1 = _queue_fifo_10_empty ? queue_10_enq_bits_vs1 : queue_dataOut_10_vs1;
  assign queue_10_deq_bits_vs2 = _queue_fifo_10_empty ? queue_10_enq_bits_vs2 : queue_dataOut_10_vs2;
  assign queue_10_deq_bits_vd = _queue_fifo_10_empty ? queue_10_enq_bits_vd : queue_dataOut_10_vd;
  assign queue_10_deq_bits_loadStoreEEW = _queue_fifo_10_empty ? queue_10_enq_bits_loadStoreEEW : queue_dataOut_10_loadStoreEEW;
  assign queue_10_deq_bits_mask = _queue_fifo_10_empty ? queue_10_enq_bits_mask : queue_dataOut_10_mask;
  assign queue_10_deq_bits_segment = _queue_fifo_10_empty ? queue_10_enq_bits_segment : queue_dataOut_10_segment;
  assign queue_10_deq_bits_readFromScalar = _queue_fifo_10_empty ? queue_10_enq_bits_readFromScalar : queue_dataOut_10_readFromScalar;
  assign queue_10_deq_bits_csrInterface_vl = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vl : queue_dataOut_10_csrInterface_vl;
  assign queue_10_deq_bits_csrInterface_vStart = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vStart : queue_dataOut_10_csrInterface_vStart;
  assign queue_10_deq_bits_csrInterface_vlmul = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vlmul : queue_dataOut_10_csrInterface_vlmul;
  assign queue_10_deq_bits_csrInterface_vSew = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vSew : queue_dataOut_10_csrInterface_vSew;
  assign queue_10_deq_bits_csrInterface_vxrm = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vxrm : queue_dataOut_10_csrInterface_vxrm;
  assign queue_10_deq_bits_csrInterface_vta = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vta : queue_dataOut_10_csrInterface_vta;
  assign queue_10_deq_bits_csrInterface_vma = _queue_fifo_10_empty ? queue_10_enq_bits_csrInterface_vma : queue_dataOut_10_csrInterface_vma;
  wire         laneVec_10_laneRequest_bits_issueInst = laneRequestSinkWire_10_ready & laneRequestSinkWire_10_valid;
  reg          releasePipe_pipe_v_10;
  wire         releasePipe_pipe_out_10_valid = releasePipe_pipe_v_10;
  wire         laneRequestSourceWire_10_ready;
  wire         validSource_10_valid = laneRequestSourceWire_10_ready & laneRequestSourceWire_10_valid;
  reg  [2:0]   tokenCheck_counter_10;
  wire [2:0]   tokenCheck_counterChange_10 = validSource_10_valid ? 3'h1 : 3'h7;
  assign tokenCheck_10 = ~(tokenCheck_counter_10[2]);
  assign laneRequestSourceWire_10_ready = tokenCheck_10;
  assign queue_10_enq_valid = validSink_10_valid;
  assign queue_10_enq_bits_instructionIndex = validSink_10_bits_instructionIndex;
  assign queue_10_enq_bits_decodeResult_orderReduce = validSink_10_bits_decodeResult_orderReduce;
  assign queue_10_enq_bits_decodeResult_floatMul = validSink_10_bits_decodeResult_floatMul;
  assign queue_10_enq_bits_decodeResult_fpExecutionType = validSink_10_bits_decodeResult_fpExecutionType;
  assign queue_10_enq_bits_decodeResult_float = validSink_10_bits_decodeResult_float;
  assign queue_10_enq_bits_decodeResult_specialSlot = validSink_10_bits_decodeResult_specialSlot;
  assign queue_10_enq_bits_decodeResult_topUop = validSink_10_bits_decodeResult_topUop;
  assign queue_10_enq_bits_decodeResult_popCount = validSink_10_bits_decodeResult_popCount;
  assign queue_10_enq_bits_decodeResult_ffo = validSink_10_bits_decodeResult_ffo;
  assign queue_10_enq_bits_decodeResult_average = validSink_10_bits_decodeResult_average;
  assign queue_10_enq_bits_decodeResult_reverse = validSink_10_bits_decodeResult_reverse;
  assign queue_10_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_10_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_10_enq_bits_decodeResult_scheduler = validSink_10_bits_decodeResult_scheduler;
  assign queue_10_enq_bits_decodeResult_sReadVD = validSink_10_bits_decodeResult_sReadVD;
  assign queue_10_enq_bits_decodeResult_vtype = validSink_10_bits_decodeResult_vtype;
  assign queue_10_enq_bits_decodeResult_sWrite = validSink_10_bits_decodeResult_sWrite;
  assign queue_10_enq_bits_decodeResult_crossRead = validSink_10_bits_decodeResult_crossRead;
  assign queue_10_enq_bits_decodeResult_crossWrite = validSink_10_bits_decodeResult_crossWrite;
  assign queue_10_enq_bits_decodeResult_maskUnit = validSink_10_bits_decodeResult_maskUnit;
  assign queue_10_enq_bits_decodeResult_special = validSink_10_bits_decodeResult_special;
  assign queue_10_enq_bits_decodeResult_saturate = validSink_10_bits_decodeResult_saturate;
  assign queue_10_enq_bits_decodeResult_vwmacc = validSink_10_bits_decodeResult_vwmacc;
  assign queue_10_enq_bits_decodeResult_readOnly = validSink_10_bits_decodeResult_readOnly;
  assign queue_10_enq_bits_decodeResult_maskSource = validSink_10_bits_decodeResult_maskSource;
  assign queue_10_enq_bits_decodeResult_maskDestination = validSink_10_bits_decodeResult_maskDestination;
  assign queue_10_enq_bits_decodeResult_maskLogic = validSink_10_bits_decodeResult_maskLogic;
  assign queue_10_enq_bits_decodeResult_uop = validSink_10_bits_decodeResult_uop;
  assign queue_10_enq_bits_decodeResult_iota = validSink_10_bits_decodeResult_iota;
  assign queue_10_enq_bits_decodeResult_mv = validSink_10_bits_decodeResult_mv;
  assign queue_10_enq_bits_decodeResult_extend = validSink_10_bits_decodeResult_extend;
  assign queue_10_enq_bits_decodeResult_unOrderWrite = validSink_10_bits_decodeResult_unOrderWrite;
  assign queue_10_enq_bits_decodeResult_compress = validSink_10_bits_decodeResult_compress;
  assign queue_10_enq_bits_decodeResult_gather16 = validSink_10_bits_decodeResult_gather16;
  assign queue_10_enq_bits_decodeResult_gather = validSink_10_bits_decodeResult_gather;
  assign queue_10_enq_bits_decodeResult_slid = validSink_10_bits_decodeResult_slid;
  assign queue_10_enq_bits_decodeResult_targetRd = validSink_10_bits_decodeResult_targetRd;
  assign queue_10_enq_bits_decodeResult_widenReduce = validSink_10_bits_decodeResult_widenReduce;
  assign queue_10_enq_bits_decodeResult_red = validSink_10_bits_decodeResult_red;
  assign queue_10_enq_bits_decodeResult_nr = validSink_10_bits_decodeResult_nr;
  assign queue_10_enq_bits_decodeResult_itype = validSink_10_bits_decodeResult_itype;
  assign queue_10_enq_bits_decodeResult_unsigned1 = validSink_10_bits_decodeResult_unsigned1;
  assign queue_10_enq_bits_decodeResult_unsigned0 = validSink_10_bits_decodeResult_unsigned0;
  assign queue_10_enq_bits_decodeResult_other = validSink_10_bits_decodeResult_other;
  assign queue_10_enq_bits_decodeResult_multiCycle = validSink_10_bits_decodeResult_multiCycle;
  assign queue_10_enq_bits_decodeResult_divider = validSink_10_bits_decodeResult_divider;
  assign queue_10_enq_bits_decodeResult_multiplier = validSink_10_bits_decodeResult_multiplier;
  assign queue_10_enq_bits_decodeResult_shift = validSink_10_bits_decodeResult_shift;
  assign queue_10_enq_bits_decodeResult_adder = validSink_10_bits_decodeResult_adder;
  assign queue_10_enq_bits_decodeResult_logic = validSink_10_bits_decodeResult_logic;
  assign queue_10_enq_bits_loadStore = validSink_10_bits_loadStore;
  assign queue_10_enq_bits_issueInst = validSink_10_bits_issueInst;
  assign queue_10_enq_bits_store = validSink_10_bits_store;
  assign queue_10_enq_bits_special = validSink_10_bits_special;
  assign queue_10_enq_bits_lsWholeReg = validSink_10_bits_lsWholeReg;
  assign queue_10_enq_bits_vs1 = validSink_10_bits_vs1;
  assign queue_10_enq_bits_vs2 = validSink_10_bits_vs2;
  assign queue_10_enq_bits_vd = validSink_10_bits_vd;
  assign queue_10_enq_bits_loadStoreEEW = validSink_10_bits_loadStoreEEW;
  assign queue_10_enq_bits_mask = validSink_10_bits_mask;
  assign queue_10_enq_bits_segment = validSink_10_bits_segment;
  assign queue_10_enq_bits_readFromScalar = validSink_10_bits_readFromScalar;
  assign queue_10_enq_bits_csrInterface_vl = validSink_10_bits_csrInterface_vl;
  assign queue_10_enq_bits_csrInterface_vStart = validSink_10_bits_csrInterface_vStart;
  assign queue_10_enq_bits_csrInterface_vlmul = validSink_10_bits_csrInterface_vlmul;
  assign queue_10_enq_bits_csrInterface_vSew = validSink_10_bits_csrInterface_vSew;
  assign queue_10_enq_bits_csrInterface_vxrm = validSink_10_bits_csrInterface_vxrm;
  assign queue_10_enq_bits_csrInterface_vta = validSink_10_bits_csrInterface_vta;
  assign queue_10_enq_bits_csrInterface_vma = validSink_10_bits_csrInterface_vma;
  reg          shifterReg_10_0_valid;
  assign validSink_10_valid = shifterReg_10_0_valid;
  reg  [2:0]   shifterReg_10_0_bits_instructionIndex;
  assign validSink_10_bits_instructionIndex = shifterReg_10_0_bits_instructionIndex;
  reg          shifterReg_10_0_bits_decodeResult_orderReduce;
  assign validSink_10_bits_decodeResult_orderReduce = shifterReg_10_0_bits_decodeResult_orderReduce;
  reg          shifterReg_10_0_bits_decodeResult_floatMul;
  assign validSink_10_bits_decodeResult_floatMul = shifterReg_10_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_10_0_bits_decodeResult_fpExecutionType;
  assign validSink_10_bits_decodeResult_fpExecutionType = shifterReg_10_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_10_0_bits_decodeResult_float;
  assign validSink_10_bits_decodeResult_float = shifterReg_10_0_bits_decodeResult_float;
  reg          shifterReg_10_0_bits_decodeResult_specialSlot;
  assign validSink_10_bits_decodeResult_specialSlot = shifterReg_10_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_10_0_bits_decodeResult_topUop;
  assign validSink_10_bits_decodeResult_topUop = shifterReg_10_0_bits_decodeResult_topUop;
  reg          shifterReg_10_0_bits_decodeResult_popCount;
  assign validSink_10_bits_decodeResult_popCount = shifterReg_10_0_bits_decodeResult_popCount;
  reg          shifterReg_10_0_bits_decodeResult_ffo;
  assign validSink_10_bits_decodeResult_ffo = shifterReg_10_0_bits_decodeResult_ffo;
  reg          shifterReg_10_0_bits_decodeResult_average;
  assign validSink_10_bits_decodeResult_average = shifterReg_10_0_bits_decodeResult_average;
  reg          shifterReg_10_0_bits_decodeResult_reverse;
  assign validSink_10_bits_decodeResult_reverse = shifterReg_10_0_bits_decodeResult_reverse;
  reg          shifterReg_10_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_10_bits_decodeResult_dontNeedExecuteInLane = shifterReg_10_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_10_0_bits_decodeResult_scheduler;
  assign validSink_10_bits_decodeResult_scheduler = shifterReg_10_0_bits_decodeResult_scheduler;
  reg          shifterReg_10_0_bits_decodeResult_sReadVD;
  assign validSink_10_bits_decodeResult_sReadVD = shifterReg_10_0_bits_decodeResult_sReadVD;
  reg          shifterReg_10_0_bits_decodeResult_vtype;
  assign validSink_10_bits_decodeResult_vtype = shifterReg_10_0_bits_decodeResult_vtype;
  reg          shifterReg_10_0_bits_decodeResult_sWrite;
  assign validSink_10_bits_decodeResult_sWrite = shifterReg_10_0_bits_decodeResult_sWrite;
  reg          shifterReg_10_0_bits_decodeResult_crossRead;
  assign validSink_10_bits_decodeResult_crossRead = shifterReg_10_0_bits_decodeResult_crossRead;
  reg          shifterReg_10_0_bits_decodeResult_crossWrite;
  assign validSink_10_bits_decodeResult_crossWrite = shifterReg_10_0_bits_decodeResult_crossWrite;
  reg          shifterReg_10_0_bits_decodeResult_maskUnit;
  assign validSink_10_bits_decodeResult_maskUnit = shifterReg_10_0_bits_decodeResult_maskUnit;
  reg          shifterReg_10_0_bits_decodeResult_special;
  assign validSink_10_bits_decodeResult_special = shifterReg_10_0_bits_decodeResult_special;
  reg          shifterReg_10_0_bits_decodeResult_saturate;
  assign validSink_10_bits_decodeResult_saturate = shifterReg_10_0_bits_decodeResult_saturate;
  reg          shifterReg_10_0_bits_decodeResult_vwmacc;
  assign validSink_10_bits_decodeResult_vwmacc = shifterReg_10_0_bits_decodeResult_vwmacc;
  reg          shifterReg_10_0_bits_decodeResult_readOnly;
  assign validSink_10_bits_decodeResult_readOnly = shifterReg_10_0_bits_decodeResult_readOnly;
  reg          shifterReg_10_0_bits_decodeResult_maskSource;
  assign validSink_10_bits_decodeResult_maskSource = shifterReg_10_0_bits_decodeResult_maskSource;
  reg          shifterReg_10_0_bits_decodeResult_maskDestination;
  assign validSink_10_bits_decodeResult_maskDestination = shifterReg_10_0_bits_decodeResult_maskDestination;
  reg          shifterReg_10_0_bits_decodeResult_maskLogic;
  assign validSink_10_bits_decodeResult_maskLogic = shifterReg_10_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_10_0_bits_decodeResult_uop;
  assign validSink_10_bits_decodeResult_uop = shifterReg_10_0_bits_decodeResult_uop;
  reg          shifterReg_10_0_bits_decodeResult_iota;
  assign validSink_10_bits_decodeResult_iota = shifterReg_10_0_bits_decodeResult_iota;
  reg          shifterReg_10_0_bits_decodeResult_mv;
  assign validSink_10_bits_decodeResult_mv = shifterReg_10_0_bits_decodeResult_mv;
  reg          shifterReg_10_0_bits_decodeResult_extend;
  assign validSink_10_bits_decodeResult_extend = shifterReg_10_0_bits_decodeResult_extend;
  reg          shifterReg_10_0_bits_decodeResult_unOrderWrite;
  assign validSink_10_bits_decodeResult_unOrderWrite = shifterReg_10_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_10_0_bits_decodeResult_compress;
  assign validSink_10_bits_decodeResult_compress = shifterReg_10_0_bits_decodeResult_compress;
  reg          shifterReg_10_0_bits_decodeResult_gather16;
  assign validSink_10_bits_decodeResult_gather16 = shifterReg_10_0_bits_decodeResult_gather16;
  reg          shifterReg_10_0_bits_decodeResult_gather;
  assign validSink_10_bits_decodeResult_gather = shifterReg_10_0_bits_decodeResult_gather;
  reg          shifterReg_10_0_bits_decodeResult_slid;
  assign validSink_10_bits_decodeResult_slid = shifterReg_10_0_bits_decodeResult_slid;
  reg          shifterReg_10_0_bits_decodeResult_targetRd;
  assign validSink_10_bits_decodeResult_targetRd = shifterReg_10_0_bits_decodeResult_targetRd;
  reg          shifterReg_10_0_bits_decodeResult_widenReduce;
  assign validSink_10_bits_decodeResult_widenReduce = shifterReg_10_0_bits_decodeResult_widenReduce;
  reg          shifterReg_10_0_bits_decodeResult_red;
  assign validSink_10_bits_decodeResult_red = shifterReg_10_0_bits_decodeResult_red;
  reg          shifterReg_10_0_bits_decodeResult_nr;
  assign validSink_10_bits_decodeResult_nr = shifterReg_10_0_bits_decodeResult_nr;
  reg          shifterReg_10_0_bits_decodeResult_itype;
  assign validSink_10_bits_decodeResult_itype = shifterReg_10_0_bits_decodeResult_itype;
  reg          shifterReg_10_0_bits_decodeResult_unsigned1;
  assign validSink_10_bits_decodeResult_unsigned1 = shifterReg_10_0_bits_decodeResult_unsigned1;
  reg          shifterReg_10_0_bits_decodeResult_unsigned0;
  assign validSink_10_bits_decodeResult_unsigned0 = shifterReg_10_0_bits_decodeResult_unsigned0;
  reg          shifterReg_10_0_bits_decodeResult_other;
  assign validSink_10_bits_decodeResult_other = shifterReg_10_0_bits_decodeResult_other;
  reg          shifterReg_10_0_bits_decodeResult_multiCycle;
  assign validSink_10_bits_decodeResult_multiCycle = shifterReg_10_0_bits_decodeResult_multiCycle;
  reg          shifterReg_10_0_bits_decodeResult_divider;
  assign validSink_10_bits_decodeResult_divider = shifterReg_10_0_bits_decodeResult_divider;
  reg          shifterReg_10_0_bits_decodeResult_multiplier;
  assign validSink_10_bits_decodeResult_multiplier = shifterReg_10_0_bits_decodeResult_multiplier;
  reg          shifterReg_10_0_bits_decodeResult_shift;
  assign validSink_10_bits_decodeResult_shift = shifterReg_10_0_bits_decodeResult_shift;
  reg          shifterReg_10_0_bits_decodeResult_adder;
  assign validSink_10_bits_decodeResult_adder = shifterReg_10_0_bits_decodeResult_adder;
  reg          shifterReg_10_0_bits_decodeResult_logic;
  assign validSink_10_bits_decodeResult_logic = shifterReg_10_0_bits_decodeResult_logic;
  reg          shifterReg_10_0_bits_loadStore;
  assign validSink_10_bits_loadStore = shifterReg_10_0_bits_loadStore;
  reg          shifterReg_10_0_bits_issueInst;
  assign validSink_10_bits_issueInst = shifterReg_10_0_bits_issueInst;
  reg          shifterReg_10_0_bits_store;
  assign validSink_10_bits_store = shifterReg_10_0_bits_store;
  reg          shifterReg_10_0_bits_special;
  assign validSink_10_bits_special = shifterReg_10_0_bits_special;
  reg          shifterReg_10_0_bits_lsWholeReg;
  assign validSink_10_bits_lsWholeReg = shifterReg_10_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_10_0_bits_vs1;
  assign validSink_10_bits_vs1 = shifterReg_10_0_bits_vs1;
  reg  [4:0]   shifterReg_10_0_bits_vs2;
  assign validSink_10_bits_vs2 = shifterReg_10_0_bits_vs2;
  reg  [4:0]   shifterReg_10_0_bits_vd;
  assign validSink_10_bits_vd = shifterReg_10_0_bits_vd;
  reg  [1:0]   shifterReg_10_0_bits_loadStoreEEW;
  assign validSink_10_bits_loadStoreEEW = shifterReg_10_0_bits_loadStoreEEW;
  reg          shifterReg_10_0_bits_mask;
  assign validSink_10_bits_mask = shifterReg_10_0_bits_mask;
  reg  [2:0]   shifterReg_10_0_bits_segment;
  assign validSink_10_bits_segment = shifterReg_10_0_bits_segment;
  reg  [31:0]  shifterReg_10_0_bits_readFromScalar;
  assign validSink_10_bits_readFromScalar = shifterReg_10_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_10_0_bits_csrInterface_vl;
  assign validSink_10_bits_csrInterface_vl = shifterReg_10_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_10_0_bits_csrInterface_vStart;
  assign validSink_10_bits_csrInterface_vStart = shifterReg_10_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_10_0_bits_csrInterface_vlmul;
  assign validSink_10_bits_csrInterface_vlmul = shifterReg_10_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_10_0_bits_csrInterface_vSew;
  assign validSink_10_bits_csrInterface_vSew = shifterReg_10_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_10_0_bits_csrInterface_vxrm;
  assign validSink_10_bits_csrInterface_vxrm = shifterReg_10_0_bits_csrInterface_vxrm;
  reg          shifterReg_10_0_bits_csrInterface_vta;
  assign validSink_10_bits_csrInterface_vta = shifterReg_10_0_bits_csrInterface_vta;
  reg          shifterReg_10_0_bits_csrInterface_vma;
  assign validSink_10_bits_csrInterface_vma = shifterReg_10_0_bits_csrInterface_vma;
  wire         shifterValid_10 = shifterReg_10_0_valid | validSource_10_valid;
  wire         validSink_11_valid;
  wire [2:0]   validSink_11_bits_instructionIndex;
  wire         validSink_11_bits_decodeResult_orderReduce;
  wire         validSink_11_bits_decodeResult_floatMul;
  wire [1:0]   validSink_11_bits_decodeResult_fpExecutionType;
  wire         validSink_11_bits_decodeResult_float;
  wire         validSink_11_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_11_bits_decodeResult_topUop;
  wire         validSink_11_bits_decodeResult_popCount;
  wire         validSink_11_bits_decodeResult_ffo;
  wire         validSink_11_bits_decodeResult_average;
  wire         validSink_11_bits_decodeResult_reverse;
  wire         validSink_11_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_11_bits_decodeResult_scheduler;
  wire         validSink_11_bits_decodeResult_sReadVD;
  wire         validSink_11_bits_decodeResult_vtype;
  wire         validSink_11_bits_decodeResult_sWrite;
  wire         validSink_11_bits_decodeResult_crossRead;
  wire         validSink_11_bits_decodeResult_crossWrite;
  wire         validSink_11_bits_decodeResult_maskUnit;
  wire         validSink_11_bits_decodeResult_special;
  wire         validSink_11_bits_decodeResult_saturate;
  wire         validSink_11_bits_decodeResult_vwmacc;
  wire         validSink_11_bits_decodeResult_readOnly;
  wire         validSink_11_bits_decodeResult_maskSource;
  wire         validSink_11_bits_decodeResult_maskDestination;
  wire         validSink_11_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_11_bits_decodeResult_uop;
  wire         validSink_11_bits_decodeResult_iota;
  wire         validSink_11_bits_decodeResult_mv;
  wire         validSink_11_bits_decodeResult_extend;
  wire         validSink_11_bits_decodeResult_unOrderWrite;
  wire         validSink_11_bits_decodeResult_compress;
  wire         validSink_11_bits_decodeResult_gather16;
  wire         validSink_11_bits_decodeResult_gather;
  wire         validSink_11_bits_decodeResult_slid;
  wire         validSink_11_bits_decodeResult_targetRd;
  wire         validSink_11_bits_decodeResult_widenReduce;
  wire         validSink_11_bits_decodeResult_red;
  wire         validSink_11_bits_decodeResult_nr;
  wire         validSink_11_bits_decodeResult_itype;
  wire         validSink_11_bits_decodeResult_unsigned1;
  wire         validSink_11_bits_decodeResult_unsigned0;
  wire         validSink_11_bits_decodeResult_other;
  wire         validSink_11_bits_decodeResult_multiCycle;
  wire         validSink_11_bits_decodeResult_divider;
  wire         validSink_11_bits_decodeResult_multiplier;
  wire         validSink_11_bits_decodeResult_shift;
  wire         validSink_11_bits_decodeResult_adder;
  wire         validSink_11_bits_decodeResult_logic;
  wire         validSink_11_bits_loadStore;
  wire         validSink_11_bits_issueInst;
  wire         validSink_11_bits_store;
  wire         validSink_11_bits_special;
  wire         validSink_11_bits_lsWholeReg;
  wire [4:0]   validSink_11_bits_vs1;
  wire [4:0]   validSink_11_bits_vs2;
  wire [4:0]   validSink_11_bits_vd;
  wire [1:0]   validSink_11_bits_loadStoreEEW;
  wire         validSink_11_bits_mask;
  wire [2:0]   validSink_11_bits_segment;
  wire [31:0]  validSink_11_bits_readFromScalar;
  wire [11:0]  validSink_11_bits_csrInterface_vl;
  wire [11:0]  validSink_11_bits_csrInterface_vStart;
  wire [2:0]   validSink_11_bits_csrInterface_vlmul;
  wire [1:0]   validSink_11_bits_csrInterface_vSew;
  wire [1:0]   validSink_11_bits_csrInterface_vxrm;
  wire         validSink_11_bits_csrInterface_vta;
  wire         validSink_11_bits_csrInterface_vma;
  wire         laneRequestSinkWire_11_valid = queue_11_deq_valid;
  wire [2:0]   laneRequestSinkWire_11_bits_instructionIndex = queue_11_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_11_bits_decodeResult_orderReduce = queue_11_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_11_bits_decodeResult_floatMul = queue_11_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_11_bits_decodeResult_fpExecutionType = queue_11_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_11_bits_decodeResult_float = queue_11_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_11_bits_decodeResult_specialSlot = queue_11_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_11_bits_decodeResult_topUop = queue_11_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_11_bits_decodeResult_popCount = queue_11_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_11_bits_decodeResult_ffo = queue_11_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_11_bits_decodeResult_average = queue_11_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_11_bits_decodeResult_reverse = queue_11_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_11_bits_decodeResult_dontNeedExecuteInLane = queue_11_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_11_bits_decodeResult_scheduler = queue_11_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_11_bits_decodeResult_sReadVD = queue_11_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_11_bits_decodeResult_vtype = queue_11_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_11_bits_decodeResult_sWrite = queue_11_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_11_bits_decodeResult_crossRead = queue_11_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_11_bits_decodeResult_crossWrite = queue_11_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_11_bits_decodeResult_maskUnit = queue_11_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_11_bits_decodeResult_special = queue_11_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_11_bits_decodeResult_saturate = queue_11_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_11_bits_decodeResult_vwmacc = queue_11_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_11_bits_decodeResult_readOnly = queue_11_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_11_bits_decodeResult_maskSource = queue_11_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_11_bits_decodeResult_maskDestination = queue_11_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_11_bits_decodeResult_maskLogic = queue_11_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_11_bits_decodeResult_uop = queue_11_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_11_bits_decodeResult_iota = queue_11_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_11_bits_decodeResult_mv = queue_11_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_11_bits_decodeResult_extend = queue_11_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_11_bits_decodeResult_unOrderWrite = queue_11_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_11_bits_decodeResult_compress = queue_11_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_11_bits_decodeResult_gather16 = queue_11_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_11_bits_decodeResult_gather = queue_11_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_11_bits_decodeResult_slid = queue_11_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_11_bits_decodeResult_targetRd = queue_11_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_11_bits_decodeResult_widenReduce = queue_11_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_11_bits_decodeResult_red = queue_11_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_11_bits_decodeResult_nr = queue_11_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_11_bits_decodeResult_itype = queue_11_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_11_bits_decodeResult_unsigned1 = queue_11_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_11_bits_decodeResult_unsigned0 = queue_11_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_11_bits_decodeResult_other = queue_11_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_11_bits_decodeResult_multiCycle = queue_11_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_11_bits_decodeResult_divider = queue_11_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_11_bits_decodeResult_multiplier = queue_11_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_11_bits_decodeResult_shift = queue_11_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_11_bits_decodeResult_adder = queue_11_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_11_bits_decodeResult_logic = queue_11_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_11_bits_loadStore = queue_11_deq_bits_loadStore;
  wire         laneRequestSinkWire_11_bits_issueInst = queue_11_deq_bits_issueInst;
  wire         laneRequestSinkWire_11_bits_store = queue_11_deq_bits_store;
  wire         laneRequestSinkWire_11_bits_special = queue_11_deq_bits_special;
  wire         laneRequestSinkWire_11_bits_lsWholeReg = queue_11_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_11_bits_vs1 = queue_11_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_11_bits_vs2 = queue_11_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_11_bits_vd = queue_11_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_11_bits_loadStoreEEW = queue_11_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_11_bits_mask = queue_11_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_11_bits_segment = queue_11_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_11_bits_readFromScalar = queue_11_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_11_bits_csrInterface_vl = queue_11_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_11_bits_csrInterface_vStart = queue_11_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_11_bits_csrInterface_vlmul = queue_11_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_11_bits_csrInterface_vSew = queue_11_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_11_bits_csrInterface_vxrm = queue_11_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_11_bits_csrInterface_vta = queue_11_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_11_bits_csrInterface_vma = queue_11_deq_bits_csrInterface_vma;
  wire [1:0]   queue_11_enq_bits_csrInterface_vxrm;
  wire         queue_11_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_33 = {queue_11_enq_bits_csrInterface_vxrm, queue_11_enq_bits_csrInterface_vta};
  wire         queue_11_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_33 = {queue_dataIn_lo_hi_33, queue_11_enq_bits_csrInterface_vma};
  wire [2:0]   queue_11_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_11_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_33 = {queue_11_enq_bits_csrInterface_vlmul, queue_11_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_11_enq_bits_csrInterface_vl;
  wire [11:0]  queue_11_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_33 = {queue_11_enq_bits_csrInterface_vl, queue_11_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_33 = {queue_dataIn_hi_hi_33, queue_dataIn_hi_lo_33};
  wire         queue_11_enq_bits_decodeResult_shift;
  wire         queue_11_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_11 = {queue_11_enq_bits_decodeResult_shift, queue_11_enq_bits_decodeResult_adder};
  wire         queue_11_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_11 = {queue_dataIn_lo_lo_lo_lo_hi_11, queue_11_enq_bits_decodeResult_logic};
  wire         queue_11_enq_bits_decodeResult_multiCycle;
  wire         queue_11_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_11 = {queue_11_enq_bits_decodeResult_multiCycle, queue_11_enq_bits_decodeResult_divider};
  wire         queue_11_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_11 = {queue_dataIn_lo_lo_lo_hi_hi_11, queue_11_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_11 = {queue_dataIn_lo_lo_lo_hi_11, queue_dataIn_lo_lo_lo_lo_11};
  wire         queue_11_enq_bits_decodeResult_unsigned1;
  wire         queue_11_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_11 = {queue_11_enq_bits_decodeResult_unsigned1, queue_11_enq_bits_decodeResult_unsigned0};
  wire         queue_11_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_11 = {queue_dataIn_lo_lo_hi_lo_hi_11, queue_11_enq_bits_decodeResult_other};
  wire         queue_11_enq_bits_decodeResult_red;
  wire         queue_11_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_11 = {queue_11_enq_bits_decodeResult_red, queue_11_enq_bits_decodeResult_nr};
  wire         queue_11_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_11 = {queue_dataIn_lo_lo_hi_hi_hi_11, queue_11_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_22 = {queue_dataIn_lo_lo_hi_hi_11, queue_dataIn_lo_lo_hi_lo_11};
  wire [11:0]  queue_dataIn_lo_lo_22 = {queue_dataIn_lo_lo_hi_22, queue_dataIn_lo_lo_lo_11};
  wire         queue_11_enq_bits_decodeResult_slid;
  wire         queue_11_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_11 = {queue_11_enq_bits_decodeResult_slid, queue_11_enq_bits_decodeResult_targetRd};
  wire         queue_11_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_11 = {queue_dataIn_lo_hi_lo_lo_hi_11, queue_11_enq_bits_decodeResult_widenReduce};
  wire         queue_11_enq_bits_decodeResult_compress;
  wire         queue_11_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_11 = {queue_11_enq_bits_decodeResult_compress, queue_11_enq_bits_decodeResult_gather16};
  wire         queue_11_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_11 = {queue_dataIn_lo_hi_lo_hi_hi_11, queue_11_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_22 = {queue_dataIn_lo_hi_lo_hi_11, queue_dataIn_lo_hi_lo_lo_11};
  wire         queue_11_enq_bits_decodeResult_mv;
  wire         queue_11_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_11 = {queue_11_enq_bits_decodeResult_mv, queue_11_enq_bits_decodeResult_extend};
  wire         queue_11_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_11 = {queue_dataIn_lo_hi_hi_lo_hi_11, queue_11_enq_bits_decodeResult_unOrderWrite};
  wire         queue_11_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_11_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_11 = {queue_11_enq_bits_decodeResult_maskLogic, queue_11_enq_bits_decodeResult_uop};
  wire         queue_11_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_11 = {queue_dataIn_lo_hi_hi_hi_hi_11, queue_11_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_22 = {queue_dataIn_lo_hi_hi_hi_11, queue_dataIn_lo_hi_hi_lo_11};
  wire [14:0]  queue_dataIn_lo_hi_34 = {queue_dataIn_lo_hi_hi_22, queue_dataIn_lo_hi_lo_22};
  wire [26:0]  queue_dataIn_lo_34 = {queue_dataIn_lo_hi_34, queue_dataIn_lo_lo_22};
  wire         queue_11_enq_bits_decodeResult_readOnly;
  wire         queue_11_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_11 = {queue_11_enq_bits_decodeResult_readOnly, queue_11_enq_bits_decodeResult_maskSource};
  wire         queue_11_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_11 = {queue_dataIn_hi_lo_lo_lo_hi_11, queue_11_enq_bits_decodeResult_maskDestination};
  wire         queue_11_enq_bits_decodeResult_special;
  wire         queue_11_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_11 = {queue_11_enq_bits_decodeResult_special, queue_11_enq_bits_decodeResult_saturate};
  wire         queue_11_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_11 = {queue_dataIn_hi_lo_lo_hi_hi_11, queue_11_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_22 = {queue_dataIn_hi_lo_lo_hi_11, queue_dataIn_hi_lo_lo_lo_11};
  wire         queue_11_enq_bits_decodeResult_crossRead;
  wire         queue_11_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_11 = {queue_11_enq_bits_decodeResult_crossRead, queue_11_enq_bits_decodeResult_crossWrite};
  wire         queue_11_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_11 = {queue_dataIn_hi_lo_hi_lo_hi_11, queue_11_enq_bits_decodeResult_maskUnit};
  wire         queue_11_enq_bits_decodeResult_sReadVD;
  wire         queue_11_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_11 = {queue_11_enq_bits_decodeResult_sReadVD, queue_11_enq_bits_decodeResult_vtype};
  wire         queue_11_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_11 = {queue_dataIn_hi_lo_hi_hi_hi_11, queue_11_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_22 = {queue_dataIn_hi_lo_hi_hi_11, queue_dataIn_hi_lo_hi_lo_11};
  wire [11:0]  queue_dataIn_hi_lo_34 = {queue_dataIn_hi_lo_hi_22, queue_dataIn_hi_lo_lo_22};
  wire         queue_11_enq_bits_decodeResult_reverse;
  wire         queue_11_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_11 = {queue_11_enq_bits_decodeResult_reverse, queue_11_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_11_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_11 = {queue_dataIn_hi_hi_lo_lo_hi_11, queue_11_enq_bits_decodeResult_scheduler};
  wire         queue_11_enq_bits_decodeResult_popCount;
  wire         queue_11_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_11 = {queue_11_enq_bits_decodeResult_popCount, queue_11_enq_bits_decodeResult_ffo};
  wire         queue_11_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_11 = {queue_dataIn_hi_hi_lo_hi_hi_11, queue_11_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_22 = {queue_dataIn_hi_hi_lo_hi_11, queue_dataIn_hi_hi_lo_lo_11};
  wire         queue_11_enq_bits_decodeResult_float;
  wire         queue_11_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_11 = {queue_11_enq_bits_decodeResult_float, queue_11_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_11_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_11 = {queue_dataIn_hi_hi_hi_lo_hi_11, queue_11_enq_bits_decodeResult_topUop};
  wire         queue_11_enq_bits_decodeResult_orderReduce;
  wire         queue_11_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_11 = {queue_11_enq_bits_decodeResult_orderReduce, queue_11_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_11_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_11 = {queue_dataIn_hi_hi_hi_hi_hi_11, queue_11_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_22 = {queue_dataIn_hi_hi_hi_hi_11, queue_dataIn_hi_hi_hi_lo_11};
  wire [16:0]  queue_dataIn_hi_hi_34 = {queue_dataIn_hi_hi_hi_22, queue_dataIn_hi_hi_lo_22};
  wire [28:0]  queue_dataIn_hi_34 = {queue_dataIn_hi_hi_34, queue_dataIn_hi_lo_34};
  wire [2:0]   queue_11_enq_bits_segment;
  wire [31:0]  queue_11_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_23 = {queue_11_enq_bits_segment, queue_11_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_23 = {queue_dataIn_lo_lo_hi_23, queue_dataIn_hi_33, queue_dataIn_lo_33};
  wire [1:0]   queue_11_enq_bits_loadStoreEEW;
  wire         queue_11_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_23 = {queue_11_enq_bits_loadStoreEEW, queue_11_enq_bits_mask};
  wire [4:0]   queue_11_enq_bits_vs2;
  wire [4:0]   queue_11_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_23 = {queue_11_enq_bits_vs2, queue_11_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_35 = {queue_dataIn_lo_hi_hi_23, queue_dataIn_lo_hi_lo_23};
  wire [80:0]  queue_dataIn_lo_35 = {queue_dataIn_lo_hi_35, queue_dataIn_lo_lo_23};
  wire         queue_11_enq_bits_lsWholeReg;
  wire [4:0]   queue_11_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_23 = {queue_11_enq_bits_lsWholeReg, queue_11_enq_bits_vs1};
  wire         queue_11_enq_bits_store;
  wire         queue_11_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_23 = {queue_11_enq_bits_store, queue_11_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_35 = {queue_dataIn_hi_lo_hi_23, queue_dataIn_hi_lo_lo_23};
  wire         queue_11_enq_bits_loadStore;
  wire         queue_11_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_23 = {queue_11_enq_bits_loadStore, queue_11_enq_bits_issueInst};
  wire [2:0]   queue_11_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_23 = {queue_11_enq_bits_instructionIndex, queue_dataIn_hi_34, queue_dataIn_lo_34};
  wire [60:0]  queue_dataIn_hi_hi_35 = {queue_dataIn_hi_hi_hi_23, queue_dataIn_hi_hi_lo_23};
  wire [68:0]  queue_dataIn_hi_35 = {queue_dataIn_hi_hi_35, queue_dataIn_hi_lo_35};
  wire [149:0] queue_dataIn_11 = {queue_dataIn_hi_35, queue_dataIn_lo_35};
  wire         queue_dataOut_11_csrInterface_vma = _queue_fifo_11_data_out[0];
  wire         queue_dataOut_11_csrInterface_vta = _queue_fifo_11_data_out[1];
  wire [1:0]   queue_dataOut_11_csrInterface_vxrm = _queue_fifo_11_data_out[3:2];
  wire [1:0]   queue_dataOut_11_csrInterface_vSew = _queue_fifo_11_data_out[5:4];
  wire [2:0]   queue_dataOut_11_csrInterface_vlmul = _queue_fifo_11_data_out[8:6];
  wire [11:0]  queue_dataOut_11_csrInterface_vStart = _queue_fifo_11_data_out[20:9];
  wire [11:0]  queue_dataOut_11_csrInterface_vl = _queue_fifo_11_data_out[32:21];
  wire [31:0]  queue_dataOut_11_readFromScalar = _queue_fifo_11_data_out[64:33];
  wire [2:0]   queue_dataOut_11_segment = _queue_fifo_11_data_out[67:65];
  wire         queue_dataOut_11_mask = _queue_fifo_11_data_out[68];
  wire [1:0]   queue_dataOut_11_loadStoreEEW = _queue_fifo_11_data_out[70:69];
  wire [4:0]   queue_dataOut_11_vd = _queue_fifo_11_data_out[75:71];
  wire [4:0]   queue_dataOut_11_vs2 = _queue_fifo_11_data_out[80:76];
  wire [4:0]   queue_dataOut_11_vs1 = _queue_fifo_11_data_out[85:81];
  wire         queue_dataOut_11_lsWholeReg = _queue_fifo_11_data_out[86];
  wire         queue_dataOut_11_special = _queue_fifo_11_data_out[87];
  wire         queue_dataOut_11_store = _queue_fifo_11_data_out[88];
  wire         queue_dataOut_11_issueInst = _queue_fifo_11_data_out[89];
  wire         queue_dataOut_11_loadStore = _queue_fifo_11_data_out[90];
  wire         queue_dataOut_11_decodeResult_logic = _queue_fifo_11_data_out[91];
  wire         queue_dataOut_11_decodeResult_adder = _queue_fifo_11_data_out[92];
  wire         queue_dataOut_11_decodeResult_shift = _queue_fifo_11_data_out[93];
  wire         queue_dataOut_11_decodeResult_multiplier = _queue_fifo_11_data_out[94];
  wire         queue_dataOut_11_decodeResult_divider = _queue_fifo_11_data_out[95];
  wire         queue_dataOut_11_decodeResult_multiCycle = _queue_fifo_11_data_out[96];
  wire         queue_dataOut_11_decodeResult_other = _queue_fifo_11_data_out[97];
  wire         queue_dataOut_11_decodeResult_unsigned0 = _queue_fifo_11_data_out[98];
  wire         queue_dataOut_11_decodeResult_unsigned1 = _queue_fifo_11_data_out[99];
  wire         queue_dataOut_11_decodeResult_itype = _queue_fifo_11_data_out[100];
  wire         queue_dataOut_11_decodeResult_nr = _queue_fifo_11_data_out[101];
  wire         queue_dataOut_11_decodeResult_red = _queue_fifo_11_data_out[102];
  wire         queue_dataOut_11_decodeResult_widenReduce = _queue_fifo_11_data_out[103];
  wire         queue_dataOut_11_decodeResult_targetRd = _queue_fifo_11_data_out[104];
  wire         queue_dataOut_11_decodeResult_slid = _queue_fifo_11_data_out[105];
  wire         queue_dataOut_11_decodeResult_gather = _queue_fifo_11_data_out[106];
  wire         queue_dataOut_11_decodeResult_gather16 = _queue_fifo_11_data_out[107];
  wire         queue_dataOut_11_decodeResult_compress = _queue_fifo_11_data_out[108];
  wire         queue_dataOut_11_decodeResult_unOrderWrite = _queue_fifo_11_data_out[109];
  wire         queue_dataOut_11_decodeResult_extend = _queue_fifo_11_data_out[110];
  wire         queue_dataOut_11_decodeResult_mv = _queue_fifo_11_data_out[111];
  wire         queue_dataOut_11_decodeResult_iota = _queue_fifo_11_data_out[112];
  wire [3:0]   queue_dataOut_11_decodeResult_uop = _queue_fifo_11_data_out[116:113];
  wire         queue_dataOut_11_decodeResult_maskLogic = _queue_fifo_11_data_out[117];
  wire         queue_dataOut_11_decodeResult_maskDestination = _queue_fifo_11_data_out[118];
  wire         queue_dataOut_11_decodeResult_maskSource = _queue_fifo_11_data_out[119];
  wire         queue_dataOut_11_decodeResult_readOnly = _queue_fifo_11_data_out[120];
  wire         queue_dataOut_11_decodeResult_vwmacc = _queue_fifo_11_data_out[121];
  wire         queue_dataOut_11_decodeResult_saturate = _queue_fifo_11_data_out[122];
  wire         queue_dataOut_11_decodeResult_special = _queue_fifo_11_data_out[123];
  wire         queue_dataOut_11_decodeResult_maskUnit = _queue_fifo_11_data_out[124];
  wire         queue_dataOut_11_decodeResult_crossWrite = _queue_fifo_11_data_out[125];
  wire         queue_dataOut_11_decodeResult_crossRead = _queue_fifo_11_data_out[126];
  wire         queue_dataOut_11_decodeResult_sWrite = _queue_fifo_11_data_out[127];
  wire         queue_dataOut_11_decodeResult_vtype = _queue_fifo_11_data_out[128];
  wire         queue_dataOut_11_decodeResult_sReadVD = _queue_fifo_11_data_out[129];
  wire         queue_dataOut_11_decodeResult_scheduler = _queue_fifo_11_data_out[130];
  wire         queue_dataOut_11_decodeResult_dontNeedExecuteInLane = _queue_fifo_11_data_out[131];
  wire         queue_dataOut_11_decodeResult_reverse = _queue_fifo_11_data_out[132];
  wire         queue_dataOut_11_decodeResult_average = _queue_fifo_11_data_out[133];
  wire         queue_dataOut_11_decodeResult_ffo = _queue_fifo_11_data_out[134];
  wire         queue_dataOut_11_decodeResult_popCount = _queue_fifo_11_data_out[135];
  wire [4:0]   queue_dataOut_11_decodeResult_topUop = _queue_fifo_11_data_out[140:136];
  wire         queue_dataOut_11_decodeResult_specialSlot = _queue_fifo_11_data_out[141];
  wire         queue_dataOut_11_decodeResult_float = _queue_fifo_11_data_out[142];
  wire [1:0]   queue_dataOut_11_decodeResult_fpExecutionType = _queue_fifo_11_data_out[144:143];
  wire         queue_dataOut_11_decodeResult_floatMul = _queue_fifo_11_data_out[145];
  wire         queue_dataOut_11_decodeResult_orderReduce = _queue_fifo_11_data_out[146];
  wire [2:0]   queue_dataOut_11_instructionIndex = _queue_fifo_11_data_out[149:147];
  wire         queue_11_enq_ready = ~_queue_fifo_11_full;
  wire         queue_11_enq_valid;
  assign queue_11_deq_valid = ~_queue_fifo_11_empty | queue_11_enq_valid;
  assign queue_11_deq_bits_instructionIndex = _queue_fifo_11_empty ? queue_11_enq_bits_instructionIndex : queue_dataOut_11_instructionIndex;
  assign queue_11_deq_bits_decodeResult_orderReduce = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_orderReduce : queue_dataOut_11_decodeResult_orderReduce;
  assign queue_11_deq_bits_decodeResult_floatMul = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_floatMul : queue_dataOut_11_decodeResult_floatMul;
  assign queue_11_deq_bits_decodeResult_fpExecutionType = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_fpExecutionType : queue_dataOut_11_decodeResult_fpExecutionType;
  assign queue_11_deq_bits_decodeResult_float = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_float : queue_dataOut_11_decodeResult_float;
  assign queue_11_deq_bits_decodeResult_specialSlot = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_specialSlot : queue_dataOut_11_decodeResult_specialSlot;
  assign queue_11_deq_bits_decodeResult_topUop = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_topUop : queue_dataOut_11_decodeResult_topUop;
  assign queue_11_deq_bits_decodeResult_popCount = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_popCount : queue_dataOut_11_decodeResult_popCount;
  assign queue_11_deq_bits_decodeResult_ffo = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_ffo : queue_dataOut_11_decodeResult_ffo;
  assign queue_11_deq_bits_decodeResult_average = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_average : queue_dataOut_11_decodeResult_average;
  assign queue_11_deq_bits_decodeResult_reverse = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_reverse : queue_dataOut_11_decodeResult_reverse;
  assign queue_11_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_11_decodeResult_dontNeedExecuteInLane;
  assign queue_11_deq_bits_decodeResult_scheduler = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_scheduler : queue_dataOut_11_decodeResult_scheduler;
  assign queue_11_deq_bits_decodeResult_sReadVD = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_sReadVD : queue_dataOut_11_decodeResult_sReadVD;
  assign queue_11_deq_bits_decodeResult_vtype = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_vtype : queue_dataOut_11_decodeResult_vtype;
  assign queue_11_deq_bits_decodeResult_sWrite = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_sWrite : queue_dataOut_11_decodeResult_sWrite;
  assign queue_11_deq_bits_decodeResult_crossRead = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_crossRead : queue_dataOut_11_decodeResult_crossRead;
  assign queue_11_deq_bits_decodeResult_crossWrite = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_crossWrite : queue_dataOut_11_decodeResult_crossWrite;
  assign queue_11_deq_bits_decodeResult_maskUnit = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_maskUnit : queue_dataOut_11_decodeResult_maskUnit;
  assign queue_11_deq_bits_decodeResult_special = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_special : queue_dataOut_11_decodeResult_special;
  assign queue_11_deq_bits_decodeResult_saturate = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_saturate : queue_dataOut_11_decodeResult_saturate;
  assign queue_11_deq_bits_decodeResult_vwmacc = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_vwmacc : queue_dataOut_11_decodeResult_vwmacc;
  assign queue_11_deq_bits_decodeResult_readOnly = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_readOnly : queue_dataOut_11_decodeResult_readOnly;
  assign queue_11_deq_bits_decodeResult_maskSource = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_maskSource : queue_dataOut_11_decodeResult_maskSource;
  assign queue_11_deq_bits_decodeResult_maskDestination = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_maskDestination : queue_dataOut_11_decodeResult_maskDestination;
  assign queue_11_deq_bits_decodeResult_maskLogic = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_maskLogic : queue_dataOut_11_decodeResult_maskLogic;
  assign queue_11_deq_bits_decodeResult_uop = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_uop : queue_dataOut_11_decodeResult_uop;
  assign queue_11_deq_bits_decodeResult_iota = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_iota : queue_dataOut_11_decodeResult_iota;
  assign queue_11_deq_bits_decodeResult_mv = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_mv : queue_dataOut_11_decodeResult_mv;
  assign queue_11_deq_bits_decodeResult_extend = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_extend : queue_dataOut_11_decodeResult_extend;
  assign queue_11_deq_bits_decodeResult_unOrderWrite = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_unOrderWrite : queue_dataOut_11_decodeResult_unOrderWrite;
  assign queue_11_deq_bits_decodeResult_compress = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_compress : queue_dataOut_11_decodeResult_compress;
  assign queue_11_deq_bits_decodeResult_gather16 = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_gather16 : queue_dataOut_11_decodeResult_gather16;
  assign queue_11_deq_bits_decodeResult_gather = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_gather : queue_dataOut_11_decodeResult_gather;
  assign queue_11_deq_bits_decodeResult_slid = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_slid : queue_dataOut_11_decodeResult_slid;
  assign queue_11_deq_bits_decodeResult_targetRd = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_targetRd : queue_dataOut_11_decodeResult_targetRd;
  assign queue_11_deq_bits_decodeResult_widenReduce = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_widenReduce : queue_dataOut_11_decodeResult_widenReduce;
  assign queue_11_deq_bits_decodeResult_red = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_red : queue_dataOut_11_decodeResult_red;
  assign queue_11_deq_bits_decodeResult_nr = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_nr : queue_dataOut_11_decodeResult_nr;
  assign queue_11_deq_bits_decodeResult_itype = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_itype : queue_dataOut_11_decodeResult_itype;
  assign queue_11_deq_bits_decodeResult_unsigned1 = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_unsigned1 : queue_dataOut_11_decodeResult_unsigned1;
  assign queue_11_deq_bits_decodeResult_unsigned0 = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_unsigned0 : queue_dataOut_11_decodeResult_unsigned0;
  assign queue_11_deq_bits_decodeResult_other = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_other : queue_dataOut_11_decodeResult_other;
  assign queue_11_deq_bits_decodeResult_multiCycle = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_multiCycle : queue_dataOut_11_decodeResult_multiCycle;
  assign queue_11_deq_bits_decodeResult_divider = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_divider : queue_dataOut_11_decodeResult_divider;
  assign queue_11_deq_bits_decodeResult_multiplier = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_multiplier : queue_dataOut_11_decodeResult_multiplier;
  assign queue_11_deq_bits_decodeResult_shift = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_shift : queue_dataOut_11_decodeResult_shift;
  assign queue_11_deq_bits_decodeResult_adder = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_adder : queue_dataOut_11_decodeResult_adder;
  assign queue_11_deq_bits_decodeResult_logic = _queue_fifo_11_empty ? queue_11_enq_bits_decodeResult_logic : queue_dataOut_11_decodeResult_logic;
  assign queue_11_deq_bits_loadStore = _queue_fifo_11_empty ? queue_11_enq_bits_loadStore : queue_dataOut_11_loadStore;
  assign queue_11_deq_bits_issueInst = _queue_fifo_11_empty ? queue_11_enq_bits_issueInst : queue_dataOut_11_issueInst;
  assign queue_11_deq_bits_store = _queue_fifo_11_empty ? queue_11_enq_bits_store : queue_dataOut_11_store;
  assign queue_11_deq_bits_special = _queue_fifo_11_empty ? queue_11_enq_bits_special : queue_dataOut_11_special;
  assign queue_11_deq_bits_lsWholeReg = _queue_fifo_11_empty ? queue_11_enq_bits_lsWholeReg : queue_dataOut_11_lsWholeReg;
  assign queue_11_deq_bits_vs1 = _queue_fifo_11_empty ? queue_11_enq_bits_vs1 : queue_dataOut_11_vs1;
  assign queue_11_deq_bits_vs2 = _queue_fifo_11_empty ? queue_11_enq_bits_vs2 : queue_dataOut_11_vs2;
  assign queue_11_deq_bits_vd = _queue_fifo_11_empty ? queue_11_enq_bits_vd : queue_dataOut_11_vd;
  assign queue_11_deq_bits_loadStoreEEW = _queue_fifo_11_empty ? queue_11_enq_bits_loadStoreEEW : queue_dataOut_11_loadStoreEEW;
  assign queue_11_deq_bits_mask = _queue_fifo_11_empty ? queue_11_enq_bits_mask : queue_dataOut_11_mask;
  assign queue_11_deq_bits_segment = _queue_fifo_11_empty ? queue_11_enq_bits_segment : queue_dataOut_11_segment;
  assign queue_11_deq_bits_readFromScalar = _queue_fifo_11_empty ? queue_11_enq_bits_readFromScalar : queue_dataOut_11_readFromScalar;
  assign queue_11_deq_bits_csrInterface_vl = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vl : queue_dataOut_11_csrInterface_vl;
  assign queue_11_deq_bits_csrInterface_vStart = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vStart : queue_dataOut_11_csrInterface_vStart;
  assign queue_11_deq_bits_csrInterface_vlmul = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vlmul : queue_dataOut_11_csrInterface_vlmul;
  assign queue_11_deq_bits_csrInterface_vSew = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vSew : queue_dataOut_11_csrInterface_vSew;
  assign queue_11_deq_bits_csrInterface_vxrm = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vxrm : queue_dataOut_11_csrInterface_vxrm;
  assign queue_11_deq_bits_csrInterface_vta = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vta : queue_dataOut_11_csrInterface_vta;
  assign queue_11_deq_bits_csrInterface_vma = _queue_fifo_11_empty ? queue_11_enq_bits_csrInterface_vma : queue_dataOut_11_csrInterface_vma;
  wire         laneVec_11_laneRequest_bits_issueInst = laneRequestSinkWire_11_ready & laneRequestSinkWire_11_valid;
  reg          releasePipe_pipe_v_11;
  wire         releasePipe_pipe_out_11_valid = releasePipe_pipe_v_11;
  wire         laneRequestSourceWire_11_ready;
  wire         validSource_11_valid = laneRequestSourceWire_11_ready & laneRequestSourceWire_11_valid;
  reg  [2:0]   tokenCheck_counter_11;
  wire [2:0]   tokenCheck_counterChange_11 = validSource_11_valid ? 3'h1 : 3'h7;
  assign tokenCheck_11 = ~(tokenCheck_counter_11[2]);
  assign laneRequestSourceWire_11_ready = tokenCheck_11;
  assign queue_11_enq_valid = validSink_11_valid;
  assign queue_11_enq_bits_instructionIndex = validSink_11_bits_instructionIndex;
  assign queue_11_enq_bits_decodeResult_orderReduce = validSink_11_bits_decodeResult_orderReduce;
  assign queue_11_enq_bits_decodeResult_floatMul = validSink_11_bits_decodeResult_floatMul;
  assign queue_11_enq_bits_decodeResult_fpExecutionType = validSink_11_bits_decodeResult_fpExecutionType;
  assign queue_11_enq_bits_decodeResult_float = validSink_11_bits_decodeResult_float;
  assign queue_11_enq_bits_decodeResult_specialSlot = validSink_11_bits_decodeResult_specialSlot;
  assign queue_11_enq_bits_decodeResult_topUop = validSink_11_bits_decodeResult_topUop;
  assign queue_11_enq_bits_decodeResult_popCount = validSink_11_bits_decodeResult_popCount;
  assign queue_11_enq_bits_decodeResult_ffo = validSink_11_bits_decodeResult_ffo;
  assign queue_11_enq_bits_decodeResult_average = validSink_11_bits_decodeResult_average;
  assign queue_11_enq_bits_decodeResult_reverse = validSink_11_bits_decodeResult_reverse;
  assign queue_11_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_11_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_11_enq_bits_decodeResult_scheduler = validSink_11_bits_decodeResult_scheduler;
  assign queue_11_enq_bits_decodeResult_sReadVD = validSink_11_bits_decodeResult_sReadVD;
  assign queue_11_enq_bits_decodeResult_vtype = validSink_11_bits_decodeResult_vtype;
  assign queue_11_enq_bits_decodeResult_sWrite = validSink_11_bits_decodeResult_sWrite;
  assign queue_11_enq_bits_decodeResult_crossRead = validSink_11_bits_decodeResult_crossRead;
  assign queue_11_enq_bits_decodeResult_crossWrite = validSink_11_bits_decodeResult_crossWrite;
  assign queue_11_enq_bits_decodeResult_maskUnit = validSink_11_bits_decodeResult_maskUnit;
  assign queue_11_enq_bits_decodeResult_special = validSink_11_bits_decodeResult_special;
  assign queue_11_enq_bits_decodeResult_saturate = validSink_11_bits_decodeResult_saturate;
  assign queue_11_enq_bits_decodeResult_vwmacc = validSink_11_bits_decodeResult_vwmacc;
  assign queue_11_enq_bits_decodeResult_readOnly = validSink_11_bits_decodeResult_readOnly;
  assign queue_11_enq_bits_decodeResult_maskSource = validSink_11_bits_decodeResult_maskSource;
  assign queue_11_enq_bits_decodeResult_maskDestination = validSink_11_bits_decodeResult_maskDestination;
  assign queue_11_enq_bits_decodeResult_maskLogic = validSink_11_bits_decodeResult_maskLogic;
  assign queue_11_enq_bits_decodeResult_uop = validSink_11_bits_decodeResult_uop;
  assign queue_11_enq_bits_decodeResult_iota = validSink_11_bits_decodeResult_iota;
  assign queue_11_enq_bits_decodeResult_mv = validSink_11_bits_decodeResult_mv;
  assign queue_11_enq_bits_decodeResult_extend = validSink_11_bits_decodeResult_extend;
  assign queue_11_enq_bits_decodeResult_unOrderWrite = validSink_11_bits_decodeResult_unOrderWrite;
  assign queue_11_enq_bits_decodeResult_compress = validSink_11_bits_decodeResult_compress;
  assign queue_11_enq_bits_decodeResult_gather16 = validSink_11_bits_decodeResult_gather16;
  assign queue_11_enq_bits_decodeResult_gather = validSink_11_bits_decodeResult_gather;
  assign queue_11_enq_bits_decodeResult_slid = validSink_11_bits_decodeResult_slid;
  assign queue_11_enq_bits_decodeResult_targetRd = validSink_11_bits_decodeResult_targetRd;
  assign queue_11_enq_bits_decodeResult_widenReduce = validSink_11_bits_decodeResult_widenReduce;
  assign queue_11_enq_bits_decodeResult_red = validSink_11_bits_decodeResult_red;
  assign queue_11_enq_bits_decodeResult_nr = validSink_11_bits_decodeResult_nr;
  assign queue_11_enq_bits_decodeResult_itype = validSink_11_bits_decodeResult_itype;
  assign queue_11_enq_bits_decodeResult_unsigned1 = validSink_11_bits_decodeResult_unsigned1;
  assign queue_11_enq_bits_decodeResult_unsigned0 = validSink_11_bits_decodeResult_unsigned0;
  assign queue_11_enq_bits_decodeResult_other = validSink_11_bits_decodeResult_other;
  assign queue_11_enq_bits_decodeResult_multiCycle = validSink_11_bits_decodeResult_multiCycle;
  assign queue_11_enq_bits_decodeResult_divider = validSink_11_bits_decodeResult_divider;
  assign queue_11_enq_bits_decodeResult_multiplier = validSink_11_bits_decodeResult_multiplier;
  assign queue_11_enq_bits_decodeResult_shift = validSink_11_bits_decodeResult_shift;
  assign queue_11_enq_bits_decodeResult_adder = validSink_11_bits_decodeResult_adder;
  assign queue_11_enq_bits_decodeResult_logic = validSink_11_bits_decodeResult_logic;
  assign queue_11_enq_bits_loadStore = validSink_11_bits_loadStore;
  assign queue_11_enq_bits_issueInst = validSink_11_bits_issueInst;
  assign queue_11_enq_bits_store = validSink_11_bits_store;
  assign queue_11_enq_bits_special = validSink_11_bits_special;
  assign queue_11_enq_bits_lsWholeReg = validSink_11_bits_lsWholeReg;
  assign queue_11_enq_bits_vs1 = validSink_11_bits_vs1;
  assign queue_11_enq_bits_vs2 = validSink_11_bits_vs2;
  assign queue_11_enq_bits_vd = validSink_11_bits_vd;
  assign queue_11_enq_bits_loadStoreEEW = validSink_11_bits_loadStoreEEW;
  assign queue_11_enq_bits_mask = validSink_11_bits_mask;
  assign queue_11_enq_bits_segment = validSink_11_bits_segment;
  assign queue_11_enq_bits_readFromScalar = validSink_11_bits_readFromScalar;
  assign queue_11_enq_bits_csrInterface_vl = validSink_11_bits_csrInterface_vl;
  assign queue_11_enq_bits_csrInterface_vStart = validSink_11_bits_csrInterface_vStart;
  assign queue_11_enq_bits_csrInterface_vlmul = validSink_11_bits_csrInterface_vlmul;
  assign queue_11_enq_bits_csrInterface_vSew = validSink_11_bits_csrInterface_vSew;
  assign queue_11_enq_bits_csrInterface_vxrm = validSink_11_bits_csrInterface_vxrm;
  assign queue_11_enq_bits_csrInterface_vta = validSink_11_bits_csrInterface_vta;
  assign queue_11_enq_bits_csrInterface_vma = validSink_11_bits_csrInterface_vma;
  reg          shifterReg_11_0_valid;
  assign validSink_11_valid = shifterReg_11_0_valid;
  reg  [2:0]   shifterReg_11_0_bits_instructionIndex;
  assign validSink_11_bits_instructionIndex = shifterReg_11_0_bits_instructionIndex;
  reg          shifterReg_11_0_bits_decodeResult_orderReduce;
  assign validSink_11_bits_decodeResult_orderReduce = shifterReg_11_0_bits_decodeResult_orderReduce;
  reg          shifterReg_11_0_bits_decodeResult_floatMul;
  assign validSink_11_bits_decodeResult_floatMul = shifterReg_11_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_11_0_bits_decodeResult_fpExecutionType;
  assign validSink_11_bits_decodeResult_fpExecutionType = shifterReg_11_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_11_0_bits_decodeResult_float;
  assign validSink_11_bits_decodeResult_float = shifterReg_11_0_bits_decodeResult_float;
  reg          shifterReg_11_0_bits_decodeResult_specialSlot;
  assign validSink_11_bits_decodeResult_specialSlot = shifterReg_11_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_11_0_bits_decodeResult_topUop;
  assign validSink_11_bits_decodeResult_topUop = shifterReg_11_0_bits_decodeResult_topUop;
  reg          shifterReg_11_0_bits_decodeResult_popCount;
  assign validSink_11_bits_decodeResult_popCount = shifterReg_11_0_bits_decodeResult_popCount;
  reg          shifterReg_11_0_bits_decodeResult_ffo;
  assign validSink_11_bits_decodeResult_ffo = shifterReg_11_0_bits_decodeResult_ffo;
  reg          shifterReg_11_0_bits_decodeResult_average;
  assign validSink_11_bits_decodeResult_average = shifterReg_11_0_bits_decodeResult_average;
  reg          shifterReg_11_0_bits_decodeResult_reverse;
  assign validSink_11_bits_decodeResult_reverse = shifterReg_11_0_bits_decodeResult_reverse;
  reg          shifterReg_11_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_11_bits_decodeResult_dontNeedExecuteInLane = shifterReg_11_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_11_0_bits_decodeResult_scheduler;
  assign validSink_11_bits_decodeResult_scheduler = shifterReg_11_0_bits_decodeResult_scheduler;
  reg          shifterReg_11_0_bits_decodeResult_sReadVD;
  assign validSink_11_bits_decodeResult_sReadVD = shifterReg_11_0_bits_decodeResult_sReadVD;
  reg          shifterReg_11_0_bits_decodeResult_vtype;
  assign validSink_11_bits_decodeResult_vtype = shifterReg_11_0_bits_decodeResult_vtype;
  reg          shifterReg_11_0_bits_decodeResult_sWrite;
  assign validSink_11_bits_decodeResult_sWrite = shifterReg_11_0_bits_decodeResult_sWrite;
  reg          shifterReg_11_0_bits_decodeResult_crossRead;
  assign validSink_11_bits_decodeResult_crossRead = shifterReg_11_0_bits_decodeResult_crossRead;
  reg          shifterReg_11_0_bits_decodeResult_crossWrite;
  assign validSink_11_bits_decodeResult_crossWrite = shifterReg_11_0_bits_decodeResult_crossWrite;
  reg          shifterReg_11_0_bits_decodeResult_maskUnit;
  assign validSink_11_bits_decodeResult_maskUnit = shifterReg_11_0_bits_decodeResult_maskUnit;
  reg          shifterReg_11_0_bits_decodeResult_special;
  assign validSink_11_bits_decodeResult_special = shifterReg_11_0_bits_decodeResult_special;
  reg          shifterReg_11_0_bits_decodeResult_saturate;
  assign validSink_11_bits_decodeResult_saturate = shifterReg_11_0_bits_decodeResult_saturate;
  reg          shifterReg_11_0_bits_decodeResult_vwmacc;
  assign validSink_11_bits_decodeResult_vwmacc = shifterReg_11_0_bits_decodeResult_vwmacc;
  reg          shifterReg_11_0_bits_decodeResult_readOnly;
  assign validSink_11_bits_decodeResult_readOnly = shifterReg_11_0_bits_decodeResult_readOnly;
  reg          shifterReg_11_0_bits_decodeResult_maskSource;
  assign validSink_11_bits_decodeResult_maskSource = shifterReg_11_0_bits_decodeResult_maskSource;
  reg          shifterReg_11_0_bits_decodeResult_maskDestination;
  assign validSink_11_bits_decodeResult_maskDestination = shifterReg_11_0_bits_decodeResult_maskDestination;
  reg          shifterReg_11_0_bits_decodeResult_maskLogic;
  assign validSink_11_bits_decodeResult_maskLogic = shifterReg_11_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_11_0_bits_decodeResult_uop;
  assign validSink_11_bits_decodeResult_uop = shifterReg_11_0_bits_decodeResult_uop;
  reg          shifterReg_11_0_bits_decodeResult_iota;
  assign validSink_11_bits_decodeResult_iota = shifterReg_11_0_bits_decodeResult_iota;
  reg          shifterReg_11_0_bits_decodeResult_mv;
  assign validSink_11_bits_decodeResult_mv = shifterReg_11_0_bits_decodeResult_mv;
  reg          shifterReg_11_0_bits_decodeResult_extend;
  assign validSink_11_bits_decodeResult_extend = shifterReg_11_0_bits_decodeResult_extend;
  reg          shifterReg_11_0_bits_decodeResult_unOrderWrite;
  assign validSink_11_bits_decodeResult_unOrderWrite = shifterReg_11_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_11_0_bits_decodeResult_compress;
  assign validSink_11_bits_decodeResult_compress = shifterReg_11_0_bits_decodeResult_compress;
  reg          shifterReg_11_0_bits_decodeResult_gather16;
  assign validSink_11_bits_decodeResult_gather16 = shifterReg_11_0_bits_decodeResult_gather16;
  reg          shifterReg_11_0_bits_decodeResult_gather;
  assign validSink_11_bits_decodeResult_gather = shifterReg_11_0_bits_decodeResult_gather;
  reg          shifterReg_11_0_bits_decodeResult_slid;
  assign validSink_11_bits_decodeResult_slid = shifterReg_11_0_bits_decodeResult_slid;
  reg          shifterReg_11_0_bits_decodeResult_targetRd;
  assign validSink_11_bits_decodeResult_targetRd = shifterReg_11_0_bits_decodeResult_targetRd;
  reg          shifterReg_11_0_bits_decodeResult_widenReduce;
  assign validSink_11_bits_decodeResult_widenReduce = shifterReg_11_0_bits_decodeResult_widenReduce;
  reg          shifterReg_11_0_bits_decodeResult_red;
  assign validSink_11_bits_decodeResult_red = shifterReg_11_0_bits_decodeResult_red;
  reg          shifterReg_11_0_bits_decodeResult_nr;
  assign validSink_11_bits_decodeResult_nr = shifterReg_11_0_bits_decodeResult_nr;
  reg          shifterReg_11_0_bits_decodeResult_itype;
  assign validSink_11_bits_decodeResult_itype = shifterReg_11_0_bits_decodeResult_itype;
  reg          shifterReg_11_0_bits_decodeResult_unsigned1;
  assign validSink_11_bits_decodeResult_unsigned1 = shifterReg_11_0_bits_decodeResult_unsigned1;
  reg          shifterReg_11_0_bits_decodeResult_unsigned0;
  assign validSink_11_bits_decodeResult_unsigned0 = shifterReg_11_0_bits_decodeResult_unsigned0;
  reg          shifterReg_11_0_bits_decodeResult_other;
  assign validSink_11_bits_decodeResult_other = shifterReg_11_0_bits_decodeResult_other;
  reg          shifterReg_11_0_bits_decodeResult_multiCycle;
  assign validSink_11_bits_decodeResult_multiCycle = shifterReg_11_0_bits_decodeResult_multiCycle;
  reg          shifterReg_11_0_bits_decodeResult_divider;
  assign validSink_11_bits_decodeResult_divider = shifterReg_11_0_bits_decodeResult_divider;
  reg          shifterReg_11_0_bits_decodeResult_multiplier;
  assign validSink_11_bits_decodeResult_multiplier = shifterReg_11_0_bits_decodeResult_multiplier;
  reg          shifterReg_11_0_bits_decodeResult_shift;
  assign validSink_11_bits_decodeResult_shift = shifterReg_11_0_bits_decodeResult_shift;
  reg          shifterReg_11_0_bits_decodeResult_adder;
  assign validSink_11_bits_decodeResult_adder = shifterReg_11_0_bits_decodeResult_adder;
  reg          shifterReg_11_0_bits_decodeResult_logic;
  assign validSink_11_bits_decodeResult_logic = shifterReg_11_0_bits_decodeResult_logic;
  reg          shifterReg_11_0_bits_loadStore;
  assign validSink_11_bits_loadStore = shifterReg_11_0_bits_loadStore;
  reg          shifterReg_11_0_bits_issueInst;
  assign validSink_11_bits_issueInst = shifterReg_11_0_bits_issueInst;
  reg          shifterReg_11_0_bits_store;
  assign validSink_11_bits_store = shifterReg_11_0_bits_store;
  reg          shifterReg_11_0_bits_special;
  assign validSink_11_bits_special = shifterReg_11_0_bits_special;
  reg          shifterReg_11_0_bits_lsWholeReg;
  assign validSink_11_bits_lsWholeReg = shifterReg_11_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_11_0_bits_vs1;
  assign validSink_11_bits_vs1 = shifterReg_11_0_bits_vs1;
  reg  [4:0]   shifterReg_11_0_bits_vs2;
  assign validSink_11_bits_vs2 = shifterReg_11_0_bits_vs2;
  reg  [4:0]   shifterReg_11_0_bits_vd;
  assign validSink_11_bits_vd = shifterReg_11_0_bits_vd;
  reg  [1:0]   shifterReg_11_0_bits_loadStoreEEW;
  assign validSink_11_bits_loadStoreEEW = shifterReg_11_0_bits_loadStoreEEW;
  reg          shifterReg_11_0_bits_mask;
  assign validSink_11_bits_mask = shifterReg_11_0_bits_mask;
  reg  [2:0]   shifterReg_11_0_bits_segment;
  assign validSink_11_bits_segment = shifterReg_11_0_bits_segment;
  reg  [31:0]  shifterReg_11_0_bits_readFromScalar;
  assign validSink_11_bits_readFromScalar = shifterReg_11_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_11_0_bits_csrInterface_vl;
  assign validSink_11_bits_csrInterface_vl = shifterReg_11_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_11_0_bits_csrInterface_vStart;
  assign validSink_11_bits_csrInterface_vStart = shifterReg_11_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_11_0_bits_csrInterface_vlmul;
  assign validSink_11_bits_csrInterface_vlmul = shifterReg_11_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_11_0_bits_csrInterface_vSew;
  assign validSink_11_bits_csrInterface_vSew = shifterReg_11_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_11_0_bits_csrInterface_vxrm;
  assign validSink_11_bits_csrInterface_vxrm = shifterReg_11_0_bits_csrInterface_vxrm;
  reg          shifterReg_11_0_bits_csrInterface_vta;
  assign validSink_11_bits_csrInterface_vta = shifterReg_11_0_bits_csrInterface_vta;
  reg          shifterReg_11_0_bits_csrInterface_vma;
  assign validSink_11_bits_csrInterface_vma = shifterReg_11_0_bits_csrInterface_vma;
  wire         shifterValid_11 = shifterReg_11_0_valid | validSource_11_valid;
  wire         validSink_12_valid;
  wire [2:0]   validSink_12_bits_instructionIndex;
  wire         validSink_12_bits_decodeResult_orderReduce;
  wire         validSink_12_bits_decodeResult_floatMul;
  wire [1:0]   validSink_12_bits_decodeResult_fpExecutionType;
  wire         validSink_12_bits_decodeResult_float;
  wire         validSink_12_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_12_bits_decodeResult_topUop;
  wire         validSink_12_bits_decodeResult_popCount;
  wire         validSink_12_bits_decodeResult_ffo;
  wire         validSink_12_bits_decodeResult_average;
  wire         validSink_12_bits_decodeResult_reverse;
  wire         validSink_12_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_12_bits_decodeResult_scheduler;
  wire         validSink_12_bits_decodeResult_sReadVD;
  wire         validSink_12_bits_decodeResult_vtype;
  wire         validSink_12_bits_decodeResult_sWrite;
  wire         validSink_12_bits_decodeResult_crossRead;
  wire         validSink_12_bits_decodeResult_crossWrite;
  wire         validSink_12_bits_decodeResult_maskUnit;
  wire         validSink_12_bits_decodeResult_special;
  wire         validSink_12_bits_decodeResult_saturate;
  wire         validSink_12_bits_decodeResult_vwmacc;
  wire         validSink_12_bits_decodeResult_readOnly;
  wire         validSink_12_bits_decodeResult_maskSource;
  wire         validSink_12_bits_decodeResult_maskDestination;
  wire         validSink_12_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_12_bits_decodeResult_uop;
  wire         validSink_12_bits_decodeResult_iota;
  wire         validSink_12_bits_decodeResult_mv;
  wire         validSink_12_bits_decodeResult_extend;
  wire         validSink_12_bits_decodeResult_unOrderWrite;
  wire         validSink_12_bits_decodeResult_compress;
  wire         validSink_12_bits_decodeResult_gather16;
  wire         validSink_12_bits_decodeResult_gather;
  wire         validSink_12_bits_decodeResult_slid;
  wire         validSink_12_bits_decodeResult_targetRd;
  wire         validSink_12_bits_decodeResult_widenReduce;
  wire         validSink_12_bits_decodeResult_red;
  wire         validSink_12_bits_decodeResult_nr;
  wire         validSink_12_bits_decodeResult_itype;
  wire         validSink_12_bits_decodeResult_unsigned1;
  wire         validSink_12_bits_decodeResult_unsigned0;
  wire         validSink_12_bits_decodeResult_other;
  wire         validSink_12_bits_decodeResult_multiCycle;
  wire         validSink_12_bits_decodeResult_divider;
  wire         validSink_12_bits_decodeResult_multiplier;
  wire         validSink_12_bits_decodeResult_shift;
  wire         validSink_12_bits_decodeResult_adder;
  wire         validSink_12_bits_decodeResult_logic;
  wire         validSink_12_bits_loadStore;
  wire         validSink_12_bits_issueInst;
  wire         validSink_12_bits_store;
  wire         validSink_12_bits_special;
  wire         validSink_12_bits_lsWholeReg;
  wire [4:0]   validSink_12_bits_vs1;
  wire [4:0]   validSink_12_bits_vs2;
  wire [4:0]   validSink_12_bits_vd;
  wire [1:0]   validSink_12_bits_loadStoreEEW;
  wire         validSink_12_bits_mask;
  wire [2:0]   validSink_12_bits_segment;
  wire [31:0]  validSink_12_bits_readFromScalar;
  wire [11:0]  validSink_12_bits_csrInterface_vl;
  wire [11:0]  validSink_12_bits_csrInterface_vStart;
  wire [2:0]   validSink_12_bits_csrInterface_vlmul;
  wire [1:0]   validSink_12_bits_csrInterface_vSew;
  wire [1:0]   validSink_12_bits_csrInterface_vxrm;
  wire         validSink_12_bits_csrInterface_vta;
  wire         validSink_12_bits_csrInterface_vma;
  wire         laneRequestSinkWire_12_valid = queue_12_deq_valid;
  wire [2:0]   laneRequestSinkWire_12_bits_instructionIndex = queue_12_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_12_bits_decodeResult_orderReduce = queue_12_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_12_bits_decodeResult_floatMul = queue_12_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_12_bits_decodeResult_fpExecutionType = queue_12_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_12_bits_decodeResult_float = queue_12_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_12_bits_decodeResult_specialSlot = queue_12_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_12_bits_decodeResult_topUop = queue_12_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_12_bits_decodeResult_popCount = queue_12_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_12_bits_decodeResult_ffo = queue_12_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_12_bits_decodeResult_average = queue_12_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_12_bits_decodeResult_reverse = queue_12_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_12_bits_decodeResult_dontNeedExecuteInLane = queue_12_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_12_bits_decodeResult_scheduler = queue_12_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_12_bits_decodeResult_sReadVD = queue_12_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_12_bits_decodeResult_vtype = queue_12_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_12_bits_decodeResult_sWrite = queue_12_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_12_bits_decodeResult_crossRead = queue_12_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_12_bits_decodeResult_crossWrite = queue_12_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_12_bits_decodeResult_maskUnit = queue_12_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_12_bits_decodeResult_special = queue_12_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_12_bits_decodeResult_saturate = queue_12_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_12_bits_decodeResult_vwmacc = queue_12_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_12_bits_decodeResult_readOnly = queue_12_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_12_bits_decodeResult_maskSource = queue_12_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_12_bits_decodeResult_maskDestination = queue_12_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_12_bits_decodeResult_maskLogic = queue_12_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_12_bits_decodeResult_uop = queue_12_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_12_bits_decodeResult_iota = queue_12_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_12_bits_decodeResult_mv = queue_12_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_12_bits_decodeResult_extend = queue_12_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_12_bits_decodeResult_unOrderWrite = queue_12_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_12_bits_decodeResult_compress = queue_12_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_12_bits_decodeResult_gather16 = queue_12_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_12_bits_decodeResult_gather = queue_12_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_12_bits_decodeResult_slid = queue_12_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_12_bits_decodeResult_targetRd = queue_12_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_12_bits_decodeResult_widenReduce = queue_12_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_12_bits_decodeResult_red = queue_12_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_12_bits_decodeResult_nr = queue_12_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_12_bits_decodeResult_itype = queue_12_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_12_bits_decodeResult_unsigned1 = queue_12_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_12_bits_decodeResult_unsigned0 = queue_12_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_12_bits_decodeResult_other = queue_12_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_12_bits_decodeResult_multiCycle = queue_12_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_12_bits_decodeResult_divider = queue_12_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_12_bits_decodeResult_multiplier = queue_12_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_12_bits_decodeResult_shift = queue_12_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_12_bits_decodeResult_adder = queue_12_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_12_bits_decodeResult_logic = queue_12_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_12_bits_loadStore = queue_12_deq_bits_loadStore;
  wire         laneRequestSinkWire_12_bits_issueInst = queue_12_deq_bits_issueInst;
  wire         laneRequestSinkWire_12_bits_store = queue_12_deq_bits_store;
  wire         laneRequestSinkWire_12_bits_special = queue_12_deq_bits_special;
  wire         laneRequestSinkWire_12_bits_lsWholeReg = queue_12_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_12_bits_vs1 = queue_12_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_12_bits_vs2 = queue_12_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_12_bits_vd = queue_12_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_12_bits_loadStoreEEW = queue_12_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_12_bits_mask = queue_12_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_12_bits_segment = queue_12_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_12_bits_readFromScalar = queue_12_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_12_bits_csrInterface_vl = queue_12_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_12_bits_csrInterface_vStart = queue_12_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_12_bits_csrInterface_vlmul = queue_12_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_12_bits_csrInterface_vSew = queue_12_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_12_bits_csrInterface_vxrm = queue_12_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_12_bits_csrInterface_vta = queue_12_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_12_bits_csrInterface_vma = queue_12_deq_bits_csrInterface_vma;
  wire [1:0]   queue_12_enq_bits_csrInterface_vxrm;
  wire         queue_12_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_36 = {queue_12_enq_bits_csrInterface_vxrm, queue_12_enq_bits_csrInterface_vta};
  wire         queue_12_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_36 = {queue_dataIn_lo_hi_36, queue_12_enq_bits_csrInterface_vma};
  wire [2:0]   queue_12_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_12_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_36 = {queue_12_enq_bits_csrInterface_vlmul, queue_12_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_12_enq_bits_csrInterface_vl;
  wire [11:0]  queue_12_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_36 = {queue_12_enq_bits_csrInterface_vl, queue_12_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_36 = {queue_dataIn_hi_hi_36, queue_dataIn_hi_lo_36};
  wire         queue_12_enq_bits_decodeResult_shift;
  wire         queue_12_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_12 = {queue_12_enq_bits_decodeResult_shift, queue_12_enq_bits_decodeResult_adder};
  wire         queue_12_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_12 = {queue_dataIn_lo_lo_lo_lo_hi_12, queue_12_enq_bits_decodeResult_logic};
  wire         queue_12_enq_bits_decodeResult_multiCycle;
  wire         queue_12_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_12 = {queue_12_enq_bits_decodeResult_multiCycle, queue_12_enq_bits_decodeResult_divider};
  wire         queue_12_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_12 = {queue_dataIn_lo_lo_lo_hi_hi_12, queue_12_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_12 = {queue_dataIn_lo_lo_lo_hi_12, queue_dataIn_lo_lo_lo_lo_12};
  wire         queue_12_enq_bits_decodeResult_unsigned1;
  wire         queue_12_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_12 = {queue_12_enq_bits_decodeResult_unsigned1, queue_12_enq_bits_decodeResult_unsigned0};
  wire         queue_12_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_12 = {queue_dataIn_lo_lo_hi_lo_hi_12, queue_12_enq_bits_decodeResult_other};
  wire         queue_12_enq_bits_decodeResult_red;
  wire         queue_12_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_12 = {queue_12_enq_bits_decodeResult_red, queue_12_enq_bits_decodeResult_nr};
  wire         queue_12_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_12 = {queue_dataIn_lo_lo_hi_hi_hi_12, queue_12_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_24 = {queue_dataIn_lo_lo_hi_hi_12, queue_dataIn_lo_lo_hi_lo_12};
  wire [11:0]  queue_dataIn_lo_lo_24 = {queue_dataIn_lo_lo_hi_24, queue_dataIn_lo_lo_lo_12};
  wire         queue_12_enq_bits_decodeResult_slid;
  wire         queue_12_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_12 = {queue_12_enq_bits_decodeResult_slid, queue_12_enq_bits_decodeResult_targetRd};
  wire         queue_12_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_12 = {queue_dataIn_lo_hi_lo_lo_hi_12, queue_12_enq_bits_decodeResult_widenReduce};
  wire         queue_12_enq_bits_decodeResult_compress;
  wire         queue_12_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_12 = {queue_12_enq_bits_decodeResult_compress, queue_12_enq_bits_decodeResult_gather16};
  wire         queue_12_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_12 = {queue_dataIn_lo_hi_lo_hi_hi_12, queue_12_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_24 = {queue_dataIn_lo_hi_lo_hi_12, queue_dataIn_lo_hi_lo_lo_12};
  wire         queue_12_enq_bits_decodeResult_mv;
  wire         queue_12_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_12 = {queue_12_enq_bits_decodeResult_mv, queue_12_enq_bits_decodeResult_extend};
  wire         queue_12_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_12 = {queue_dataIn_lo_hi_hi_lo_hi_12, queue_12_enq_bits_decodeResult_unOrderWrite};
  wire         queue_12_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_12_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_12 = {queue_12_enq_bits_decodeResult_maskLogic, queue_12_enq_bits_decodeResult_uop};
  wire         queue_12_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_12 = {queue_dataIn_lo_hi_hi_hi_hi_12, queue_12_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_24 = {queue_dataIn_lo_hi_hi_hi_12, queue_dataIn_lo_hi_hi_lo_12};
  wire [14:0]  queue_dataIn_lo_hi_37 = {queue_dataIn_lo_hi_hi_24, queue_dataIn_lo_hi_lo_24};
  wire [26:0]  queue_dataIn_lo_37 = {queue_dataIn_lo_hi_37, queue_dataIn_lo_lo_24};
  wire         queue_12_enq_bits_decodeResult_readOnly;
  wire         queue_12_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_12 = {queue_12_enq_bits_decodeResult_readOnly, queue_12_enq_bits_decodeResult_maskSource};
  wire         queue_12_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_12 = {queue_dataIn_hi_lo_lo_lo_hi_12, queue_12_enq_bits_decodeResult_maskDestination};
  wire         queue_12_enq_bits_decodeResult_special;
  wire         queue_12_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_12 = {queue_12_enq_bits_decodeResult_special, queue_12_enq_bits_decodeResult_saturate};
  wire         queue_12_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_12 = {queue_dataIn_hi_lo_lo_hi_hi_12, queue_12_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_24 = {queue_dataIn_hi_lo_lo_hi_12, queue_dataIn_hi_lo_lo_lo_12};
  wire         queue_12_enq_bits_decodeResult_crossRead;
  wire         queue_12_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_12 = {queue_12_enq_bits_decodeResult_crossRead, queue_12_enq_bits_decodeResult_crossWrite};
  wire         queue_12_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_12 = {queue_dataIn_hi_lo_hi_lo_hi_12, queue_12_enq_bits_decodeResult_maskUnit};
  wire         queue_12_enq_bits_decodeResult_sReadVD;
  wire         queue_12_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_12 = {queue_12_enq_bits_decodeResult_sReadVD, queue_12_enq_bits_decodeResult_vtype};
  wire         queue_12_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_12 = {queue_dataIn_hi_lo_hi_hi_hi_12, queue_12_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_24 = {queue_dataIn_hi_lo_hi_hi_12, queue_dataIn_hi_lo_hi_lo_12};
  wire [11:0]  queue_dataIn_hi_lo_37 = {queue_dataIn_hi_lo_hi_24, queue_dataIn_hi_lo_lo_24};
  wire         queue_12_enq_bits_decodeResult_reverse;
  wire         queue_12_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_12 = {queue_12_enq_bits_decodeResult_reverse, queue_12_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_12_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_12 = {queue_dataIn_hi_hi_lo_lo_hi_12, queue_12_enq_bits_decodeResult_scheduler};
  wire         queue_12_enq_bits_decodeResult_popCount;
  wire         queue_12_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_12 = {queue_12_enq_bits_decodeResult_popCount, queue_12_enq_bits_decodeResult_ffo};
  wire         queue_12_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_12 = {queue_dataIn_hi_hi_lo_hi_hi_12, queue_12_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_24 = {queue_dataIn_hi_hi_lo_hi_12, queue_dataIn_hi_hi_lo_lo_12};
  wire         queue_12_enq_bits_decodeResult_float;
  wire         queue_12_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_12 = {queue_12_enq_bits_decodeResult_float, queue_12_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_12_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_12 = {queue_dataIn_hi_hi_hi_lo_hi_12, queue_12_enq_bits_decodeResult_topUop};
  wire         queue_12_enq_bits_decodeResult_orderReduce;
  wire         queue_12_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_12 = {queue_12_enq_bits_decodeResult_orderReduce, queue_12_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_12_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_12 = {queue_dataIn_hi_hi_hi_hi_hi_12, queue_12_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_24 = {queue_dataIn_hi_hi_hi_hi_12, queue_dataIn_hi_hi_hi_lo_12};
  wire [16:0]  queue_dataIn_hi_hi_37 = {queue_dataIn_hi_hi_hi_24, queue_dataIn_hi_hi_lo_24};
  wire [28:0]  queue_dataIn_hi_37 = {queue_dataIn_hi_hi_37, queue_dataIn_hi_lo_37};
  wire [2:0]   queue_12_enq_bits_segment;
  wire [31:0]  queue_12_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_25 = {queue_12_enq_bits_segment, queue_12_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_25 = {queue_dataIn_lo_lo_hi_25, queue_dataIn_hi_36, queue_dataIn_lo_36};
  wire [1:0]   queue_12_enq_bits_loadStoreEEW;
  wire         queue_12_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_25 = {queue_12_enq_bits_loadStoreEEW, queue_12_enq_bits_mask};
  wire [4:0]   queue_12_enq_bits_vs2;
  wire [4:0]   queue_12_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_25 = {queue_12_enq_bits_vs2, queue_12_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_38 = {queue_dataIn_lo_hi_hi_25, queue_dataIn_lo_hi_lo_25};
  wire [80:0]  queue_dataIn_lo_38 = {queue_dataIn_lo_hi_38, queue_dataIn_lo_lo_25};
  wire         queue_12_enq_bits_lsWholeReg;
  wire [4:0]   queue_12_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_25 = {queue_12_enq_bits_lsWholeReg, queue_12_enq_bits_vs1};
  wire         queue_12_enq_bits_store;
  wire         queue_12_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_25 = {queue_12_enq_bits_store, queue_12_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_38 = {queue_dataIn_hi_lo_hi_25, queue_dataIn_hi_lo_lo_25};
  wire         queue_12_enq_bits_loadStore;
  wire         queue_12_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_25 = {queue_12_enq_bits_loadStore, queue_12_enq_bits_issueInst};
  wire [2:0]   queue_12_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_25 = {queue_12_enq_bits_instructionIndex, queue_dataIn_hi_37, queue_dataIn_lo_37};
  wire [60:0]  queue_dataIn_hi_hi_38 = {queue_dataIn_hi_hi_hi_25, queue_dataIn_hi_hi_lo_25};
  wire [68:0]  queue_dataIn_hi_38 = {queue_dataIn_hi_hi_38, queue_dataIn_hi_lo_38};
  wire [149:0] queue_dataIn_12 = {queue_dataIn_hi_38, queue_dataIn_lo_38};
  wire         queue_dataOut_12_csrInterface_vma = _queue_fifo_12_data_out[0];
  wire         queue_dataOut_12_csrInterface_vta = _queue_fifo_12_data_out[1];
  wire [1:0]   queue_dataOut_12_csrInterface_vxrm = _queue_fifo_12_data_out[3:2];
  wire [1:0]   queue_dataOut_12_csrInterface_vSew = _queue_fifo_12_data_out[5:4];
  wire [2:0]   queue_dataOut_12_csrInterface_vlmul = _queue_fifo_12_data_out[8:6];
  wire [11:0]  queue_dataOut_12_csrInterface_vStart = _queue_fifo_12_data_out[20:9];
  wire [11:0]  queue_dataOut_12_csrInterface_vl = _queue_fifo_12_data_out[32:21];
  wire [31:0]  queue_dataOut_12_readFromScalar = _queue_fifo_12_data_out[64:33];
  wire [2:0]   queue_dataOut_12_segment = _queue_fifo_12_data_out[67:65];
  wire         queue_dataOut_12_mask = _queue_fifo_12_data_out[68];
  wire [1:0]   queue_dataOut_12_loadStoreEEW = _queue_fifo_12_data_out[70:69];
  wire [4:0]   queue_dataOut_12_vd = _queue_fifo_12_data_out[75:71];
  wire [4:0]   queue_dataOut_12_vs2 = _queue_fifo_12_data_out[80:76];
  wire [4:0]   queue_dataOut_12_vs1 = _queue_fifo_12_data_out[85:81];
  wire         queue_dataOut_12_lsWholeReg = _queue_fifo_12_data_out[86];
  wire         queue_dataOut_12_special = _queue_fifo_12_data_out[87];
  wire         queue_dataOut_12_store = _queue_fifo_12_data_out[88];
  wire         queue_dataOut_12_issueInst = _queue_fifo_12_data_out[89];
  wire         queue_dataOut_12_loadStore = _queue_fifo_12_data_out[90];
  wire         queue_dataOut_12_decodeResult_logic = _queue_fifo_12_data_out[91];
  wire         queue_dataOut_12_decodeResult_adder = _queue_fifo_12_data_out[92];
  wire         queue_dataOut_12_decodeResult_shift = _queue_fifo_12_data_out[93];
  wire         queue_dataOut_12_decodeResult_multiplier = _queue_fifo_12_data_out[94];
  wire         queue_dataOut_12_decodeResult_divider = _queue_fifo_12_data_out[95];
  wire         queue_dataOut_12_decodeResult_multiCycle = _queue_fifo_12_data_out[96];
  wire         queue_dataOut_12_decodeResult_other = _queue_fifo_12_data_out[97];
  wire         queue_dataOut_12_decodeResult_unsigned0 = _queue_fifo_12_data_out[98];
  wire         queue_dataOut_12_decodeResult_unsigned1 = _queue_fifo_12_data_out[99];
  wire         queue_dataOut_12_decodeResult_itype = _queue_fifo_12_data_out[100];
  wire         queue_dataOut_12_decodeResult_nr = _queue_fifo_12_data_out[101];
  wire         queue_dataOut_12_decodeResult_red = _queue_fifo_12_data_out[102];
  wire         queue_dataOut_12_decodeResult_widenReduce = _queue_fifo_12_data_out[103];
  wire         queue_dataOut_12_decodeResult_targetRd = _queue_fifo_12_data_out[104];
  wire         queue_dataOut_12_decodeResult_slid = _queue_fifo_12_data_out[105];
  wire         queue_dataOut_12_decodeResult_gather = _queue_fifo_12_data_out[106];
  wire         queue_dataOut_12_decodeResult_gather16 = _queue_fifo_12_data_out[107];
  wire         queue_dataOut_12_decodeResult_compress = _queue_fifo_12_data_out[108];
  wire         queue_dataOut_12_decodeResult_unOrderWrite = _queue_fifo_12_data_out[109];
  wire         queue_dataOut_12_decodeResult_extend = _queue_fifo_12_data_out[110];
  wire         queue_dataOut_12_decodeResult_mv = _queue_fifo_12_data_out[111];
  wire         queue_dataOut_12_decodeResult_iota = _queue_fifo_12_data_out[112];
  wire [3:0]   queue_dataOut_12_decodeResult_uop = _queue_fifo_12_data_out[116:113];
  wire         queue_dataOut_12_decodeResult_maskLogic = _queue_fifo_12_data_out[117];
  wire         queue_dataOut_12_decodeResult_maskDestination = _queue_fifo_12_data_out[118];
  wire         queue_dataOut_12_decodeResult_maskSource = _queue_fifo_12_data_out[119];
  wire         queue_dataOut_12_decodeResult_readOnly = _queue_fifo_12_data_out[120];
  wire         queue_dataOut_12_decodeResult_vwmacc = _queue_fifo_12_data_out[121];
  wire         queue_dataOut_12_decodeResult_saturate = _queue_fifo_12_data_out[122];
  wire         queue_dataOut_12_decodeResult_special = _queue_fifo_12_data_out[123];
  wire         queue_dataOut_12_decodeResult_maskUnit = _queue_fifo_12_data_out[124];
  wire         queue_dataOut_12_decodeResult_crossWrite = _queue_fifo_12_data_out[125];
  wire         queue_dataOut_12_decodeResult_crossRead = _queue_fifo_12_data_out[126];
  wire         queue_dataOut_12_decodeResult_sWrite = _queue_fifo_12_data_out[127];
  wire         queue_dataOut_12_decodeResult_vtype = _queue_fifo_12_data_out[128];
  wire         queue_dataOut_12_decodeResult_sReadVD = _queue_fifo_12_data_out[129];
  wire         queue_dataOut_12_decodeResult_scheduler = _queue_fifo_12_data_out[130];
  wire         queue_dataOut_12_decodeResult_dontNeedExecuteInLane = _queue_fifo_12_data_out[131];
  wire         queue_dataOut_12_decodeResult_reverse = _queue_fifo_12_data_out[132];
  wire         queue_dataOut_12_decodeResult_average = _queue_fifo_12_data_out[133];
  wire         queue_dataOut_12_decodeResult_ffo = _queue_fifo_12_data_out[134];
  wire         queue_dataOut_12_decodeResult_popCount = _queue_fifo_12_data_out[135];
  wire [4:0]   queue_dataOut_12_decodeResult_topUop = _queue_fifo_12_data_out[140:136];
  wire         queue_dataOut_12_decodeResult_specialSlot = _queue_fifo_12_data_out[141];
  wire         queue_dataOut_12_decodeResult_float = _queue_fifo_12_data_out[142];
  wire [1:0]   queue_dataOut_12_decodeResult_fpExecutionType = _queue_fifo_12_data_out[144:143];
  wire         queue_dataOut_12_decodeResult_floatMul = _queue_fifo_12_data_out[145];
  wire         queue_dataOut_12_decodeResult_orderReduce = _queue_fifo_12_data_out[146];
  wire [2:0]   queue_dataOut_12_instructionIndex = _queue_fifo_12_data_out[149:147];
  wire         queue_12_enq_ready = ~_queue_fifo_12_full;
  wire         queue_12_enq_valid;
  assign queue_12_deq_valid = ~_queue_fifo_12_empty | queue_12_enq_valid;
  assign queue_12_deq_bits_instructionIndex = _queue_fifo_12_empty ? queue_12_enq_bits_instructionIndex : queue_dataOut_12_instructionIndex;
  assign queue_12_deq_bits_decodeResult_orderReduce = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_orderReduce : queue_dataOut_12_decodeResult_orderReduce;
  assign queue_12_deq_bits_decodeResult_floatMul = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_floatMul : queue_dataOut_12_decodeResult_floatMul;
  assign queue_12_deq_bits_decodeResult_fpExecutionType = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_fpExecutionType : queue_dataOut_12_decodeResult_fpExecutionType;
  assign queue_12_deq_bits_decodeResult_float = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_float : queue_dataOut_12_decodeResult_float;
  assign queue_12_deq_bits_decodeResult_specialSlot = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_specialSlot : queue_dataOut_12_decodeResult_specialSlot;
  assign queue_12_deq_bits_decodeResult_topUop = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_topUop : queue_dataOut_12_decodeResult_topUop;
  assign queue_12_deq_bits_decodeResult_popCount = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_popCount : queue_dataOut_12_decodeResult_popCount;
  assign queue_12_deq_bits_decodeResult_ffo = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_ffo : queue_dataOut_12_decodeResult_ffo;
  assign queue_12_deq_bits_decodeResult_average = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_average : queue_dataOut_12_decodeResult_average;
  assign queue_12_deq_bits_decodeResult_reverse = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_reverse : queue_dataOut_12_decodeResult_reverse;
  assign queue_12_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_12_decodeResult_dontNeedExecuteInLane;
  assign queue_12_deq_bits_decodeResult_scheduler = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_scheduler : queue_dataOut_12_decodeResult_scheduler;
  assign queue_12_deq_bits_decodeResult_sReadVD = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_sReadVD : queue_dataOut_12_decodeResult_sReadVD;
  assign queue_12_deq_bits_decodeResult_vtype = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_vtype : queue_dataOut_12_decodeResult_vtype;
  assign queue_12_deq_bits_decodeResult_sWrite = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_sWrite : queue_dataOut_12_decodeResult_sWrite;
  assign queue_12_deq_bits_decodeResult_crossRead = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_crossRead : queue_dataOut_12_decodeResult_crossRead;
  assign queue_12_deq_bits_decodeResult_crossWrite = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_crossWrite : queue_dataOut_12_decodeResult_crossWrite;
  assign queue_12_deq_bits_decodeResult_maskUnit = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_maskUnit : queue_dataOut_12_decodeResult_maskUnit;
  assign queue_12_deq_bits_decodeResult_special = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_special : queue_dataOut_12_decodeResult_special;
  assign queue_12_deq_bits_decodeResult_saturate = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_saturate : queue_dataOut_12_decodeResult_saturate;
  assign queue_12_deq_bits_decodeResult_vwmacc = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_vwmacc : queue_dataOut_12_decodeResult_vwmacc;
  assign queue_12_deq_bits_decodeResult_readOnly = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_readOnly : queue_dataOut_12_decodeResult_readOnly;
  assign queue_12_deq_bits_decodeResult_maskSource = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_maskSource : queue_dataOut_12_decodeResult_maskSource;
  assign queue_12_deq_bits_decodeResult_maskDestination = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_maskDestination : queue_dataOut_12_decodeResult_maskDestination;
  assign queue_12_deq_bits_decodeResult_maskLogic = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_maskLogic : queue_dataOut_12_decodeResult_maskLogic;
  assign queue_12_deq_bits_decodeResult_uop = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_uop : queue_dataOut_12_decodeResult_uop;
  assign queue_12_deq_bits_decodeResult_iota = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_iota : queue_dataOut_12_decodeResult_iota;
  assign queue_12_deq_bits_decodeResult_mv = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_mv : queue_dataOut_12_decodeResult_mv;
  assign queue_12_deq_bits_decodeResult_extend = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_extend : queue_dataOut_12_decodeResult_extend;
  assign queue_12_deq_bits_decodeResult_unOrderWrite = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_unOrderWrite : queue_dataOut_12_decodeResult_unOrderWrite;
  assign queue_12_deq_bits_decodeResult_compress = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_compress : queue_dataOut_12_decodeResult_compress;
  assign queue_12_deq_bits_decodeResult_gather16 = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_gather16 : queue_dataOut_12_decodeResult_gather16;
  assign queue_12_deq_bits_decodeResult_gather = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_gather : queue_dataOut_12_decodeResult_gather;
  assign queue_12_deq_bits_decodeResult_slid = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_slid : queue_dataOut_12_decodeResult_slid;
  assign queue_12_deq_bits_decodeResult_targetRd = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_targetRd : queue_dataOut_12_decodeResult_targetRd;
  assign queue_12_deq_bits_decodeResult_widenReduce = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_widenReduce : queue_dataOut_12_decodeResult_widenReduce;
  assign queue_12_deq_bits_decodeResult_red = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_red : queue_dataOut_12_decodeResult_red;
  assign queue_12_deq_bits_decodeResult_nr = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_nr : queue_dataOut_12_decodeResult_nr;
  assign queue_12_deq_bits_decodeResult_itype = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_itype : queue_dataOut_12_decodeResult_itype;
  assign queue_12_deq_bits_decodeResult_unsigned1 = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_unsigned1 : queue_dataOut_12_decodeResult_unsigned1;
  assign queue_12_deq_bits_decodeResult_unsigned0 = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_unsigned0 : queue_dataOut_12_decodeResult_unsigned0;
  assign queue_12_deq_bits_decodeResult_other = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_other : queue_dataOut_12_decodeResult_other;
  assign queue_12_deq_bits_decodeResult_multiCycle = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_multiCycle : queue_dataOut_12_decodeResult_multiCycle;
  assign queue_12_deq_bits_decodeResult_divider = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_divider : queue_dataOut_12_decodeResult_divider;
  assign queue_12_deq_bits_decodeResult_multiplier = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_multiplier : queue_dataOut_12_decodeResult_multiplier;
  assign queue_12_deq_bits_decodeResult_shift = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_shift : queue_dataOut_12_decodeResult_shift;
  assign queue_12_deq_bits_decodeResult_adder = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_adder : queue_dataOut_12_decodeResult_adder;
  assign queue_12_deq_bits_decodeResult_logic = _queue_fifo_12_empty ? queue_12_enq_bits_decodeResult_logic : queue_dataOut_12_decodeResult_logic;
  assign queue_12_deq_bits_loadStore = _queue_fifo_12_empty ? queue_12_enq_bits_loadStore : queue_dataOut_12_loadStore;
  assign queue_12_deq_bits_issueInst = _queue_fifo_12_empty ? queue_12_enq_bits_issueInst : queue_dataOut_12_issueInst;
  assign queue_12_deq_bits_store = _queue_fifo_12_empty ? queue_12_enq_bits_store : queue_dataOut_12_store;
  assign queue_12_deq_bits_special = _queue_fifo_12_empty ? queue_12_enq_bits_special : queue_dataOut_12_special;
  assign queue_12_deq_bits_lsWholeReg = _queue_fifo_12_empty ? queue_12_enq_bits_lsWholeReg : queue_dataOut_12_lsWholeReg;
  assign queue_12_deq_bits_vs1 = _queue_fifo_12_empty ? queue_12_enq_bits_vs1 : queue_dataOut_12_vs1;
  assign queue_12_deq_bits_vs2 = _queue_fifo_12_empty ? queue_12_enq_bits_vs2 : queue_dataOut_12_vs2;
  assign queue_12_deq_bits_vd = _queue_fifo_12_empty ? queue_12_enq_bits_vd : queue_dataOut_12_vd;
  assign queue_12_deq_bits_loadStoreEEW = _queue_fifo_12_empty ? queue_12_enq_bits_loadStoreEEW : queue_dataOut_12_loadStoreEEW;
  assign queue_12_deq_bits_mask = _queue_fifo_12_empty ? queue_12_enq_bits_mask : queue_dataOut_12_mask;
  assign queue_12_deq_bits_segment = _queue_fifo_12_empty ? queue_12_enq_bits_segment : queue_dataOut_12_segment;
  assign queue_12_deq_bits_readFromScalar = _queue_fifo_12_empty ? queue_12_enq_bits_readFromScalar : queue_dataOut_12_readFromScalar;
  assign queue_12_deq_bits_csrInterface_vl = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vl : queue_dataOut_12_csrInterface_vl;
  assign queue_12_deq_bits_csrInterface_vStart = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vStart : queue_dataOut_12_csrInterface_vStart;
  assign queue_12_deq_bits_csrInterface_vlmul = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vlmul : queue_dataOut_12_csrInterface_vlmul;
  assign queue_12_deq_bits_csrInterface_vSew = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vSew : queue_dataOut_12_csrInterface_vSew;
  assign queue_12_deq_bits_csrInterface_vxrm = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vxrm : queue_dataOut_12_csrInterface_vxrm;
  assign queue_12_deq_bits_csrInterface_vta = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vta : queue_dataOut_12_csrInterface_vta;
  assign queue_12_deq_bits_csrInterface_vma = _queue_fifo_12_empty ? queue_12_enq_bits_csrInterface_vma : queue_dataOut_12_csrInterface_vma;
  wire         laneVec_12_laneRequest_bits_issueInst = laneRequestSinkWire_12_ready & laneRequestSinkWire_12_valid;
  reg          releasePipe_pipe_v_12;
  wire         releasePipe_pipe_out_12_valid = releasePipe_pipe_v_12;
  wire         laneRequestSourceWire_12_ready;
  wire         validSource_12_valid = laneRequestSourceWire_12_ready & laneRequestSourceWire_12_valid;
  reg  [2:0]   tokenCheck_counter_12;
  wire [2:0]   tokenCheck_counterChange_12 = validSource_12_valid ? 3'h1 : 3'h7;
  assign tokenCheck_12 = ~(tokenCheck_counter_12[2]);
  assign laneRequestSourceWire_12_ready = tokenCheck_12;
  assign queue_12_enq_valid = validSink_12_valid;
  assign queue_12_enq_bits_instructionIndex = validSink_12_bits_instructionIndex;
  assign queue_12_enq_bits_decodeResult_orderReduce = validSink_12_bits_decodeResult_orderReduce;
  assign queue_12_enq_bits_decodeResult_floatMul = validSink_12_bits_decodeResult_floatMul;
  assign queue_12_enq_bits_decodeResult_fpExecutionType = validSink_12_bits_decodeResult_fpExecutionType;
  assign queue_12_enq_bits_decodeResult_float = validSink_12_bits_decodeResult_float;
  assign queue_12_enq_bits_decodeResult_specialSlot = validSink_12_bits_decodeResult_specialSlot;
  assign queue_12_enq_bits_decodeResult_topUop = validSink_12_bits_decodeResult_topUop;
  assign queue_12_enq_bits_decodeResult_popCount = validSink_12_bits_decodeResult_popCount;
  assign queue_12_enq_bits_decodeResult_ffo = validSink_12_bits_decodeResult_ffo;
  assign queue_12_enq_bits_decodeResult_average = validSink_12_bits_decodeResult_average;
  assign queue_12_enq_bits_decodeResult_reverse = validSink_12_bits_decodeResult_reverse;
  assign queue_12_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_12_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_12_enq_bits_decodeResult_scheduler = validSink_12_bits_decodeResult_scheduler;
  assign queue_12_enq_bits_decodeResult_sReadVD = validSink_12_bits_decodeResult_sReadVD;
  assign queue_12_enq_bits_decodeResult_vtype = validSink_12_bits_decodeResult_vtype;
  assign queue_12_enq_bits_decodeResult_sWrite = validSink_12_bits_decodeResult_sWrite;
  assign queue_12_enq_bits_decodeResult_crossRead = validSink_12_bits_decodeResult_crossRead;
  assign queue_12_enq_bits_decodeResult_crossWrite = validSink_12_bits_decodeResult_crossWrite;
  assign queue_12_enq_bits_decodeResult_maskUnit = validSink_12_bits_decodeResult_maskUnit;
  assign queue_12_enq_bits_decodeResult_special = validSink_12_bits_decodeResult_special;
  assign queue_12_enq_bits_decodeResult_saturate = validSink_12_bits_decodeResult_saturate;
  assign queue_12_enq_bits_decodeResult_vwmacc = validSink_12_bits_decodeResult_vwmacc;
  assign queue_12_enq_bits_decodeResult_readOnly = validSink_12_bits_decodeResult_readOnly;
  assign queue_12_enq_bits_decodeResult_maskSource = validSink_12_bits_decodeResult_maskSource;
  assign queue_12_enq_bits_decodeResult_maskDestination = validSink_12_bits_decodeResult_maskDestination;
  assign queue_12_enq_bits_decodeResult_maskLogic = validSink_12_bits_decodeResult_maskLogic;
  assign queue_12_enq_bits_decodeResult_uop = validSink_12_bits_decodeResult_uop;
  assign queue_12_enq_bits_decodeResult_iota = validSink_12_bits_decodeResult_iota;
  assign queue_12_enq_bits_decodeResult_mv = validSink_12_bits_decodeResult_mv;
  assign queue_12_enq_bits_decodeResult_extend = validSink_12_bits_decodeResult_extend;
  assign queue_12_enq_bits_decodeResult_unOrderWrite = validSink_12_bits_decodeResult_unOrderWrite;
  assign queue_12_enq_bits_decodeResult_compress = validSink_12_bits_decodeResult_compress;
  assign queue_12_enq_bits_decodeResult_gather16 = validSink_12_bits_decodeResult_gather16;
  assign queue_12_enq_bits_decodeResult_gather = validSink_12_bits_decodeResult_gather;
  assign queue_12_enq_bits_decodeResult_slid = validSink_12_bits_decodeResult_slid;
  assign queue_12_enq_bits_decodeResult_targetRd = validSink_12_bits_decodeResult_targetRd;
  assign queue_12_enq_bits_decodeResult_widenReduce = validSink_12_bits_decodeResult_widenReduce;
  assign queue_12_enq_bits_decodeResult_red = validSink_12_bits_decodeResult_red;
  assign queue_12_enq_bits_decodeResult_nr = validSink_12_bits_decodeResult_nr;
  assign queue_12_enq_bits_decodeResult_itype = validSink_12_bits_decodeResult_itype;
  assign queue_12_enq_bits_decodeResult_unsigned1 = validSink_12_bits_decodeResult_unsigned1;
  assign queue_12_enq_bits_decodeResult_unsigned0 = validSink_12_bits_decodeResult_unsigned0;
  assign queue_12_enq_bits_decodeResult_other = validSink_12_bits_decodeResult_other;
  assign queue_12_enq_bits_decodeResult_multiCycle = validSink_12_bits_decodeResult_multiCycle;
  assign queue_12_enq_bits_decodeResult_divider = validSink_12_bits_decodeResult_divider;
  assign queue_12_enq_bits_decodeResult_multiplier = validSink_12_bits_decodeResult_multiplier;
  assign queue_12_enq_bits_decodeResult_shift = validSink_12_bits_decodeResult_shift;
  assign queue_12_enq_bits_decodeResult_adder = validSink_12_bits_decodeResult_adder;
  assign queue_12_enq_bits_decodeResult_logic = validSink_12_bits_decodeResult_logic;
  assign queue_12_enq_bits_loadStore = validSink_12_bits_loadStore;
  assign queue_12_enq_bits_issueInst = validSink_12_bits_issueInst;
  assign queue_12_enq_bits_store = validSink_12_bits_store;
  assign queue_12_enq_bits_special = validSink_12_bits_special;
  assign queue_12_enq_bits_lsWholeReg = validSink_12_bits_lsWholeReg;
  assign queue_12_enq_bits_vs1 = validSink_12_bits_vs1;
  assign queue_12_enq_bits_vs2 = validSink_12_bits_vs2;
  assign queue_12_enq_bits_vd = validSink_12_bits_vd;
  assign queue_12_enq_bits_loadStoreEEW = validSink_12_bits_loadStoreEEW;
  assign queue_12_enq_bits_mask = validSink_12_bits_mask;
  assign queue_12_enq_bits_segment = validSink_12_bits_segment;
  assign queue_12_enq_bits_readFromScalar = validSink_12_bits_readFromScalar;
  assign queue_12_enq_bits_csrInterface_vl = validSink_12_bits_csrInterface_vl;
  assign queue_12_enq_bits_csrInterface_vStart = validSink_12_bits_csrInterface_vStart;
  assign queue_12_enq_bits_csrInterface_vlmul = validSink_12_bits_csrInterface_vlmul;
  assign queue_12_enq_bits_csrInterface_vSew = validSink_12_bits_csrInterface_vSew;
  assign queue_12_enq_bits_csrInterface_vxrm = validSink_12_bits_csrInterface_vxrm;
  assign queue_12_enq_bits_csrInterface_vta = validSink_12_bits_csrInterface_vta;
  assign queue_12_enq_bits_csrInterface_vma = validSink_12_bits_csrInterface_vma;
  reg          shifterReg_12_0_valid;
  assign validSink_12_valid = shifterReg_12_0_valid;
  reg  [2:0]   shifterReg_12_0_bits_instructionIndex;
  assign validSink_12_bits_instructionIndex = shifterReg_12_0_bits_instructionIndex;
  reg          shifterReg_12_0_bits_decodeResult_orderReduce;
  assign validSink_12_bits_decodeResult_orderReduce = shifterReg_12_0_bits_decodeResult_orderReduce;
  reg          shifterReg_12_0_bits_decodeResult_floatMul;
  assign validSink_12_bits_decodeResult_floatMul = shifterReg_12_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_12_0_bits_decodeResult_fpExecutionType;
  assign validSink_12_bits_decodeResult_fpExecutionType = shifterReg_12_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_12_0_bits_decodeResult_float;
  assign validSink_12_bits_decodeResult_float = shifterReg_12_0_bits_decodeResult_float;
  reg          shifterReg_12_0_bits_decodeResult_specialSlot;
  assign validSink_12_bits_decodeResult_specialSlot = shifterReg_12_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_12_0_bits_decodeResult_topUop;
  assign validSink_12_bits_decodeResult_topUop = shifterReg_12_0_bits_decodeResult_topUop;
  reg          shifterReg_12_0_bits_decodeResult_popCount;
  assign validSink_12_bits_decodeResult_popCount = shifterReg_12_0_bits_decodeResult_popCount;
  reg          shifterReg_12_0_bits_decodeResult_ffo;
  assign validSink_12_bits_decodeResult_ffo = shifterReg_12_0_bits_decodeResult_ffo;
  reg          shifterReg_12_0_bits_decodeResult_average;
  assign validSink_12_bits_decodeResult_average = shifterReg_12_0_bits_decodeResult_average;
  reg          shifterReg_12_0_bits_decodeResult_reverse;
  assign validSink_12_bits_decodeResult_reverse = shifterReg_12_0_bits_decodeResult_reverse;
  reg          shifterReg_12_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_12_bits_decodeResult_dontNeedExecuteInLane = shifterReg_12_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_12_0_bits_decodeResult_scheduler;
  assign validSink_12_bits_decodeResult_scheduler = shifterReg_12_0_bits_decodeResult_scheduler;
  reg          shifterReg_12_0_bits_decodeResult_sReadVD;
  assign validSink_12_bits_decodeResult_sReadVD = shifterReg_12_0_bits_decodeResult_sReadVD;
  reg          shifterReg_12_0_bits_decodeResult_vtype;
  assign validSink_12_bits_decodeResult_vtype = shifterReg_12_0_bits_decodeResult_vtype;
  reg          shifterReg_12_0_bits_decodeResult_sWrite;
  assign validSink_12_bits_decodeResult_sWrite = shifterReg_12_0_bits_decodeResult_sWrite;
  reg          shifterReg_12_0_bits_decodeResult_crossRead;
  assign validSink_12_bits_decodeResult_crossRead = shifterReg_12_0_bits_decodeResult_crossRead;
  reg          shifterReg_12_0_bits_decodeResult_crossWrite;
  assign validSink_12_bits_decodeResult_crossWrite = shifterReg_12_0_bits_decodeResult_crossWrite;
  reg          shifterReg_12_0_bits_decodeResult_maskUnit;
  assign validSink_12_bits_decodeResult_maskUnit = shifterReg_12_0_bits_decodeResult_maskUnit;
  reg          shifterReg_12_0_bits_decodeResult_special;
  assign validSink_12_bits_decodeResult_special = shifterReg_12_0_bits_decodeResult_special;
  reg          shifterReg_12_0_bits_decodeResult_saturate;
  assign validSink_12_bits_decodeResult_saturate = shifterReg_12_0_bits_decodeResult_saturate;
  reg          shifterReg_12_0_bits_decodeResult_vwmacc;
  assign validSink_12_bits_decodeResult_vwmacc = shifterReg_12_0_bits_decodeResult_vwmacc;
  reg          shifterReg_12_0_bits_decodeResult_readOnly;
  assign validSink_12_bits_decodeResult_readOnly = shifterReg_12_0_bits_decodeResult_readOnly;
  reg          shifterReg_12_0_bits_decodeResult_maskSource;
  assign validSink_12_bits_decodeResult_maskSource = shifterReg_12_0_bits_decodeResult_maskSource;
  reg          shifterReg_12_0_bits_decodeResult_maskDestination;
  assign validSink_12_bits_decodeResult_maskDestination = shifterReg_12_0_bits_decodeResult_maskDestination;
  reg          shifterReg_12_0_bits_decodeResult_maskLogic;
  assign validSink_12_bits_decodeResult_maskLogic = shifterReg_12_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_12_0_bits_decodeResult_uop;
  assign validSink_12_bits_decodeResult_uop = shifterReg_12_0_bits_decodeResult_uop;
  reg          shifterReg_12_0_bits_decodeResult_iota;
  assign validSink_12_bits_decodeResult_iota = shifterReg_12_0_bits_decodeResult_iota;
  reg          shifterReg_12_0_bits_decodeResult_mv;
  assign validSink_12_bits_decodeResult_mv = shifterReg_12_0_bits_decodeResult_mv;
  reg          shifterReg_12_0_bits_decodeResult_extend;
  assign validSink_12_bits_decodeResult_extend = shifterReg_12_0_bits_decodeResult_extend;
  reg          shifterReg_12_0_bits_decodeResult_unOrderWrite;
  assign validSink_12_bits_decodeResult_unOrderWrite = shifterReg_12_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_12_0_bits_decodeResult_compress;
  assign validSink_12_bits_decodeResult_compress = shifterReg_12_0_bits_decodeResult_compress;
  reg          shifterReg_12_0_bits_decodeResult_gather16;
  assign validSink_12_bits_decodeResult_gather16 = shifterReg_12_0_bits_decodeResult_gather16;
  reg          shifterReg_12_0_bits_decodeResult_gather;
  assign validSink_12_bits_decodeResult_gather = shifterReg_12_0_bits_decodeResult_gather;
  reg          shifterReg_12_0_bits_decodeResult_slid;
  assign validSink_12_bits_decodeResult_slid = shifterReg_12_0_bits_decodeResult_slid;
  reg          shifterReg_12_0_bits_decodeResult_targetRd;
  assign validSink_12_bits_decodeResult_targetRd = shifterReg_12_0_bits_decodeResult_targetRd;
  reg          shifterReg_12_0_bits_decodeResult_widenReduce;
  assign validSink_12_bits_decodeResult_widenReduce = shifterReg_12_0_bits_decodeResult_widenReduce;
  reg          shifterReg_12_0_bits_decodeResult_red;
  assign validSink_12_bits_decodeResult_red = shifterReg_12_0_bits_decodeResult_red;
  reg          shifterReg_12_0_bits_decodeResult_nr;
  assign validSink_12_bits_decodeResult_nr = shifterReg_12_0_bits_decodeResult_nr;
  reg          shifterReg_12_0_bits_decodeResult_itype;
  assign validSink_12_bits_decodeResult_itype = shifterReg_12_0_bits_decodeResult_itype;
  reg          shifterReg_12_0_bits_decodeResult_unsigned1;
  assign validSink_12_bits_decodeResult_unsigned1 = shifterReg_12_0_bits_decodeResult_unsigned1;
  reg          shifterReg_12_0_bits_decodeResult_unsigned0;
  assign validSink_12_bits_decodeResult_unsigned0 = shifterReg_12_0_bits_decodeResult_unsigned0;
  reg          shifterReg_12_0_bits_decodeResult_other;
  assign validSink_12_bits_decodeResult_other = shifterReg_12_0_bits_decodeResult_other;
  reg          shifterReg_12_0_bits_decodeResult_multiCycle;
  assign validSink_12_bits_decodeResult_multiCycle = shifterReg_12_0_bits_decodeResult_multiCycle;
  reg          shifterReg_12_0_bits_decodeResult_divider;
  assign validSink_12_bits_decodeResult_divider = shifterReg_12_0_bits_decodeResult_divider;
  reg          shifterReg_12_0_bits_decodeResult_multiplier;
  assign validSink_12_bits_decodeResult_multiplier = shifterReg_12_0_bits_decodeResult_multiplier;
  reg          shifterReg_12_0_bits_decodeResult_shift;
  assign validSink_12_bits_decodeResult_shift = shifterReg_12_0_bits_decodeResult_shift;
  reg          shifterReg_12_0_bits_decodeResult_adder;
  assign validSink_12_bits_decodeResult_adder = shifterReg_12_0_bits_decodeResult_adder;
  reg          shifterReg_12_0_bits_decodeResult_logic;
  assign validSink_12_bits_decodeResult_logic = shifterReg_12_0_bits_decodeResult_logic;
  reg          shifterReg_12_0_bits_loadStore;
  assign validSink_12_bits_loadStore = shifterReg_12_0_bits_loadStore;
  reg          shifterReg_12_0_bits_issueInst;
  assign validSink_12_bits_issueInst = shifterReg_12_0_bits_issueInst;
  reg          shifterReg_12_0_bits_store;
  assign validSink_12_bits_store = shifterReg_12_0_bits_store;
  reg          shifterReg_12_0_bits_special;
  assign validSink_12_bits_special = shifterReg_12_0_bits_special;
  reg          shifterReg_12_0_bits_lsWholeReg;
  assign validSink_12_bits_lsWholeReg = shifterReg_12_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_12_0_bits_vs1;
  assign validSink_12_bits_vs1 = shifterReg_12_0_bits_vs1;
  reg  [4:0]   shifterReg_12_0_bits_vs2;
  assign validSink_12_bits_vs2 = shifterReg_12_0_bits_vs2;
  reg  [4:0]   shifterReg_12_0_bits_vd;
  assign validSink_12_bits_vd = shifterReg_12_0_bits_vd;
  reg  [1:0]   shifterReg_12_0_bits_loadStoreEEW;
  assign validSink_12_bits_loadStoreEEW = shifterReg_12_0_bits_loadStoreEEW;
  reg          shifterReg_12_0_bits_mask;
  assign validSink_12_bits_mask = shifterReg_12_0_bits_mask;
  reg  [2:0]   shifterReg_12_0_bits_segment;
  assign validSink_12_bits_segment = shifterReg_12_0_bits_segment;
  reg  [31:0]  shifterReg_12_0_bits_readFromScalar;
  assign validSink_12_bits_readFromScalar = shifterReg_12_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_12_0_bits_csrInterface_vl;
  assign validSink_12_bits_csrInterface_vl = shifterReg_12_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_12_0_bits_csrInterface_vStart;
  assign validSink_12_bits_csrInterface_vStart = shifterReg_12_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_12_0_bits_csrInterface_vlmul;
  assign validSink_12_bits_csrInterface_vlmul = shifterReg_12_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_12_0_bits_csrInterface_vSew;
  assign validSink_12_bits_csrInterface_vSew = shifterReg_12_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_12_0_bits_csrInterface_vxrm;
  assign validSink_12_bits_csrInterface_vxrm = shifterReg_12_0_bits_csrInterface_vxrm;
  reg          shifterReg_12_0_bits_csrInterface_vta;
  assign validSink_12_bits_csrInterface_vta = shifterReg_12_0_bits_csrInterface_vta;
  reg          shifterReg_12_0_bits_csrInterface_vma;
  assign validSink_12_bits_csrInterface_vma = shifterReg_12_0_bits_csrInterface_vma;
  wire         shifterValid_12 = shifterReg_12_0_valid | validSource_12_valid;
  wire         validSink_13_valid;
  wire [2:0]   validSink_13_bits_instructionIndex;
  wire         validSink_13_bits_decodeResult_orderReduce;
  wire         validSink_13_bits_decodeResult_floatMul;
  wire [1:0]   validSink_13_bits_decodeResult_fpExecutionType;
  wire         validSink_13_bits_decodeResult_float;
  wire         validSink_13_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_13_bits_decodeResult_topUop;
  wire         validSink_13_bits_decodeResult_popCount;
  wire         validSink_13_bits_decodeResult_ffo;
  wire         validSink_13_bits_decodeResult_average;
  wire         validSink_13_bits_decodeResult_reverse;
  wire         validSink_13_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_13_bits_decodeResult_scheduler;
  wire         validSink_13_bits_decodeResult_sReadVD;
  wire         validSink_13_bits_decodeResult_vtype;
  wire         validSink_13_bits_decodeResult_sWrite;
  wire         validSink_13_bits_decodeResult_crossRead;
  wire         validSink_13_bits_decodeResult_crossWrite;
  wire         validSink_13_bits_decodeResult_maskUnit;
  wire         validSink_13_bits_decodeResult_special;
  wire         validSink_13_bits_decodeResult_saturate;
  wire         validSink_13_bits_decodeResult_vwmacc;
  wire         validSink_13_bits_decodeResult_readOnly;
  wire         validSink_13_bits_decodeResult_maskSource;
  wire         validSink_13_bits_decodeResult_maskDestination;
  wire         validSink_13_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_13_bits_decodeResult_uop;
  wire         validSink_13_bits_decodeResult_iota;
  wire         validSink_13_bits_decodeResult_mv;
  wire         validSink_13_bits_decodeResult_extend;
  wire         validSink_13_bits_decodeResult_unOrderWrite;
  wire         validSink_13_bits_decodeResult_compress;
  wire         validSink_13_bits_decodeResult_gather16;
  wire         validSink_13_bits_decodeResult_gather;
  wire         validSink_13_bits_decodeResult_slid;
  wire         validSink_13_bits_decodeResult_targetRd;
  wire         validSink_13_bits_decodeResult_widenReduce;
  wire         validSink_13_bits_decodeResult_red;
  wire         validSink_13_bits_decodeResult_nr;
  wire         validSink_13_bits_decodeResult_itype;
  wire         validSink_13_bits_decodeResult_unsigned1;
  wire         validSink_13_bits_decodeResult_unsigned0;
  wire         validSink_13_bits_decodeResult_other;
  wire         validSink_13_bits_decodeResult_multiCycle;
  wire         validSink_13_bits_decodeResult_divider;
  wire         validSink_13_bits_decodeResult_multiplier;
  wire         validSink_13_bits_decodeResult_shift;
  wire         validSink_13_bits_decodeResult_adder;
  wire         validSink_13_bits_decodeResult_logic;
  wire         validSink_13_bits_loadStore;
  wire         validSink_13_bits_issueInst;
  wire         validSink_13_bits_store;
  wire         validSink_13_bits_special;
  wire         validSink_13_bits_lsWholeReg;
  wire [4:0]   validSink_13_bits_vs1;
  wire [4:0]   validSink_13_bits_vs2;
  wire [4:0]   validSink_13_bits_vd;
  wire [1:0]   validSink_13_bits_loadStoreEEW;
  wire         validSink_13_bits_mask;
  wire [2:0]   validSink_13_bits_segment;
  wire [31:0]  validSink_13_bits_readFromScalar;
  wire [11:0]  validSink_13_bits_csrInterface_vl;
  wire [11:0]  validSink_13_bits_csrInterface_vStart;
  wire [2:0]   validSink_13_bits_csrInterface_vlmul;
  wire [1:0]   validSink_13_bits_csrInterface_vSew;
  wire [1:0]   validSink_13_bits_csrInterface_vxrm;
  wire         validSink_13_bits_csrInterface_vta;
  wire         validSink_13_bits_csrInterface_vma;
  wire         laneRequestSinkWire_13_valid = queue_13_deq_valid;
  wire [2:0]   laneRequestSinkWire_13_bits_instructionIndex = queue_13_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_13_bits_decodeResult_orderReduce = queue_13_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_13_bits_decodeResult_floatMul = queue_13_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_13_bits_decodeResult_fpExecutionType = queue_13_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_13_bits_decodeResult_float = queue_13_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_13_bits_decodeResult_specialSlot = queue_13_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_13_bits_decodeResult_topUop = queue_13_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_13_bits_decodeResult_popCount = queue_13_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_13_bits_decodeResult_ffo = queue_13_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_13_bits_decodeResult_average = queue_13_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_13_bits_decodeResult_reverse = queue_13_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_13_bits_decodeResult_dontNeedExecuteInLane = queue_13_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_13_bits_decodeResult_scheduler = queue_13_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_13_bits_decodeResult_sReadVD = queue_13_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_13_bits_decodeResult_vtype = queue_13_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_13_bits_decodeResult_sWrite = queue_13_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_13_bits_decodeResult_crossRead = queue_13_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_13_bits_decodeResult_crossWrite = queue_13_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_13_bits_decodeResult_maskUnit = queue_13_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_13_bits_decodeResult_special = queue_13_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_13_bits_decodeResult_saturate = queue_13_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_13_bits_decodeResult_vwmacc = queue_13_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_13_bits_decodeResult_readOnly = queue_13_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_13_bits_decodeResult_maskSource = queue_13_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_13_bits_decodeResult_maskDestination = queue_13_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_13_bits_decodeResult_maskLogic = queue_13_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_13_bits_decodeResult_uop = queue_13_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_13_bits_decodeResult_iota = queue_13_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_13_bits_decodeResult_mv = queue_13_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_13_bits_decodeResult_extend = queue_13_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_13_bits_decodeResult_unOrderWrite = queue_13_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_13_bits_decodeResult_compress = queue_13_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_13_bits_decodeResult_gather16 = queue_13_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_13_bits_decodeResult_gather = queue_13_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_13_bits_decodeResult_slid = queue_13_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_13_bits_decodeResult_targetRd = queue_13_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_13_bits_decodeResult_widenReduce = queue_13_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_13_bits_decodeResult_red = queue_13_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_13_bits_decodeResult_nr = queue_13_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_13_bits_decodeResult_itype = queue_13_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_13_bits_decodeResult_unsigned1 = queue_13_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_13_bits_decodeResult_unsigned0 = queue_13_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_13_bits_decodeResult_other = queue_13_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_13_bits_decodeResult_multiCycle = queue_13_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_13_bits_decodeResult_divider = queue_13_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_13_bits_decodeResult_multiplier = queue_13_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_13_bits_decodeResult_shift = queue_13_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_13_bits_decodeResult_adder = queue_13_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_13_bits_decodeResult_logic = queue_13_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_13_bits_loadStore = queue_13_deq_bits_loadStore;
  wire         laneRequestSinkWire_13_bits_issueInst = queue_13_deq_bits_issueInst;
  wire         laneRequestSinkWire_13_bits_store = queue_13_deq_bits_store;
  wire         laneRequestSinkWire_13_bits_special = queue_13_deq_bits_special;
  wire         laneRequestSinkWire_13_bits_lsWholeReg = queue_13_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_13_bits_vs1 = queue_13_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_13_bits_vs2 = queue_13_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_13_bits_vd = queue_13_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_13_bits_loadStoreEEW = queue_13_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_13_bits_mask = queue_13_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_13_bits_segment = queue_13_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_13_bits_readFromScalar = queue_13_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_13_bits_csrInterface_vl = queue_13_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_13_bits_csrInterface_vStart = queue_13_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_13_bits_csrInterface_vlmul = queue_13_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_13_bits_csrInterface_vSew = queue_13_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_13_bits_csrInterface_vxrm = queue_13_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_13_bits_csrInterface_vta = queue_13_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_13_bits_csrInterface_vma = queue_13_deq_bits_csrInterface_vma;
  wire [1:0]   queue_13_enq_bits_csrInterface_vxrm;
  wire         queue_13_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_39 = {queue_13_enq_bits_csrInterface_vxrm, queue_13_enq_bits_csrInterface_vta};
  wire         queue_13_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_39 = {queue_dataIn_lo_hi_39, queue_13_enq_bits_csrInterface_vma};
  wire [2:0]   queue_13_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_13_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_39 = {queue_13_enq_bits_csrInterface_vlmul, queue_13_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_13_enq_bits_csrInterface_vl;
  wire [11:0]  queue_13_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_39 = {queue_13_enq_bits_csrInterface_vl, queue_13_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_39 = {queue_dataIn_hi_hi_39, queue_dataIn_hi_lo_39};
  wire         queue_13_enq_bits_decodeResult_shift;
  wire         queue_13_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_13 = {queue_13_enq_bits_decodeResult_shift, queue_13_enq_bits_decodeResult_adder};
  wire         queue_13_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_13 = {queue_dataIn_lo_lo_lo_lo_hi_13, queue_13_enq_bits_decodeResult_logic};
  wire         queue_13_enq_bits_decodeResult_multiCycle;
  wire         queue_13_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_13 = {queue_13_enq_bits_decodeResult_multiCycle, queue_13_enq_bits_decodeResult_divider};
  wire         queue_13_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_13 = {queue_dataIn_lo_lo_lo_hi_hi_13, queue_13_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_13 = {queue_dataIn_lo_lo_lo_hi_13, queue_dataIn_lo_lo_lo_lo_13};
  wire         queue_13_enq_bits_decodeResult_unsigned1;
  wire         queue_13_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_13 = {queue_13_enq_bits_decodeResult_unsigned1, queue_13_enq_bits_decodeResult_unsigned0};
  wire         queue_13_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_13 = {queue_dataIn_lo_lo_hi_lo_hi_13, queue_13_enq_bits_decodeResult_other};
  wire         queue_13_enq_bits_decodeResult_red;
  wire         queue_13_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_13 = {queue_13_enq_bits_decodeResult_red, queue_13_enq_bits_decodeResult_nr};
  wire         queue_13_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_13 = {queue_dataIn_lo_lo_hi_hi_hi_13, queue_13_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_26 = {queue_dataIn_lo_lo_hi_hi_13, queue_dataIn_lo_lo_hi_lo_13};
  wire [11:0]  queue_dataIn_lo_lo_26 = {queue_dataIn_lo_lo_hi_26, queue_dataIn_lo_lo_lo_13};
  wire         queue_13_enq_bits_decodeResult_slid;
  wire         queue_13_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_13 = {queue_13_enq_bits_decodeResult_slid, queue_13_enq_bits_decodeResult_targetRd};
  wire         queue_13_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_13 = {queue_dataIn_lo_hi_lo_lo_hi_13, queue_13_enq_bits_decodeResult_widenReduce};
  wire         queue_13_enq_bits_decodeResult_compress;
  wire         queue_13_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_13 = {queue_13_enq_bits_decodeResult_compress, queue_13_enq_bits_decodeResult_gather16};
  wire         queue_13_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_13 = {queue_dataIn_lo_hi_lo_hi_hi_13, queue_13_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_26 = {queue_dataIn_lo_hi_lo_hi_13, queue_dataIn_lo_hi_lo_lo_13};
  wire         queue_13_enq_bits_decodeResult_mv;
  wire         queue_13_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_13 = {queue_13_enq_bits_decodeResult_mv, queue_13_enq_bits_decodeResult_extend};
  wire         queue_13_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_13 = {queue_dataIn_lo_hi_hi_lo_hi_13, queue_13_enq_bits_decodeResult_unOrderWrite};
  wire         queue_13_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_13_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_13 = {queue_13_enq_bits_decodeResult_maskLogic, queue_13_enq_bits_decodeResult_uop};
  wire         queue_13_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_13 = {queue_dataIn_lo_hi_hi_hi_hi_13, queue_13_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_26 = {queue_dataIn_lo_hi_hi_hi_13, queue_dataIn_lo_hi_hi_lo_13};
  wire [14:0]  queue_dataIn_lo_hi_40 = {queue_dataIn_lo_hi_hi_26, queue_dataIn_lo_hi_lo_26};
  wire [26:0]  queue_dataIn_lo_40 = {queue_dataIn_lo_hi_40, queue_dataIn_lo_lo_26};
  wire         queue_13_enq_bits_decodeResult_readOnly;
  wire         queue_13_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_13 = {queue_13_enq_bits_decodeResult_readOnly, queue_13_enq_bits_decodeResult_maskSource};
  wire         queue_13_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_13 = {queue_dataIn_hi_lo_lo_lo_hi_13, queue_13_enq_bits_decodeResult_maskDestination};
  wire         queue_13_enq_bits_decodeResult_special;
  wire         queue_13_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_13 = {queue_13_enq_bits_decodeResult_special, queue_13_enq_bits_decodeResult_saturate};
  wire         queue_13_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_13 = {queue_dataIn_hi_lo_lo_hi_hi_13, queue_13_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_26 = {queue_dataIn_hi_lo_lo_hi_13, queue_dataIn_hi_lo_lo_lo_13};
  wire         queue_13_enq_bits_decodeResult_crossRead;
  wire         queue_13_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_13 = {queue_13_enq_bits_decodeResult_crossRead, queue_13_enq_bits_decodeResult_crossWrite};
  wire         queue_13_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_13 = {queue_dataIn_hi_lo_hi_lo_hi_13, queue_13_enq_bits_decodeResult_maskUnit};
  wire         queue_13_enq_bits_decodeResult_sReadVD;
  wire         queue_13_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_13 = {queue_13_enq_bits_decodeResult_sReadVD, queue_13_enq_bits_decodeResult_vtype};
  wire         queue_13_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_13 = {queue_dataIn_hi_lo_hi_hi_hi_13, queue_13_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_26 = {queue_dataIn_hi_lo_hi_hi_13, queue_dataIn_hi_lo_hi_lo_13};
  wire [11:0]  queue_dataIn_hi_lo_40 = {queue_dataIn_hi_lo_hi_26, queue_dataIn_hi_lo_lo_26};
  wire         queue_13_enq_bits_decodeResult_reverse;
  wire         queue_13_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_13 = {queue_13_enq_bits_decodeResult_reverse, queue_13_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_13_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_13 = {queue_dataIn_hi_hi_lo_lo_hi_13, queue_13_enq_bits_decodeResult_scheduler};
  wire         queue_13_enq_bits_decodeResult_popCount;
  wire         queue_13_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_13 = {queue_13_enq_bits_decodeResult_popCount, queue_13_enq_bits_decodeResult_ffo};
  wire         queue_13_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_13 = {queue_dataIn_hi_hi_lo_hi_hi_13, queue_13_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_26 = {queue_dataIn_hi_hi_lo_hi_13, queue_dataIn_hi_hi_lo_lo_13};
  wire         queue_13_enq_bits_decodeResult_float;
  wire         queue_13_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_13 = {queue_13_enq_bits_decodeResult_float, queue_13_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_13_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_13 = {queue_dataIn_hi_hi_hi_lo_hi_13, queue_13_enq_bits_decodeResult_topUop};
  wire         queue_13_enq_bits_decodeResult_orderReduce;
  wire         queue_13_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_13 = {queue_13_enq_bits_decodeResult_orderReduce, queue_13_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_13_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_13 = {queue_dataIn_hi_hi_hi_hi_hi_13, queue_13_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_26 = {queue_dataIn_hi_hi_hi_hi_13, queue_dataIn_hi_hi_hi_lo_13};
  wire [16:0]  queue_dataIn_hi_hi_40 = {queue_dataIn_hi_hi_hi_26, queue_dataIn_hi_hi_lo_26};
  wire [28:0]  queue_dataIn_hi_40 = {queue_dataIn_hi_hi_40, queue_dataIn_hi_lo_40};
  wire [2:0]   queue_13_enq_bits_segment;
  wire [31:0]  queue_13_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_27 = {queue_13_enq_bits_segment, queue_13_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_27 = {queue_dataIn_lo_lo_hi_27, queue_dataIn_hi_39, queue_dataIn_lo_39};
  wire [1:0]   queue_13_enq_bits_loadStoreEEW;
  wire         queue_13_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_27 = {queue_13_enq_bits_loadStoreEEW, queue_13_enq_bits_mask};
  wire [4:0]   queue_13_enq_bits_vs2;
  wire [4:0]   queue_13_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_27 = {queue_13_enq_bits_vs2, queue_13_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_41 = {queue_dataIn_lo_hi_hi_27, queue_dataIn_lo_hi_lo_27};
  wire [80:0]  queue_dataIn_lo_41 = {queue_dataIn_lo_hi_41, queue_dataIn_lo_lo_27};
  wire         queue_13_enq_bits_lsWholeReg;
  wire [4:0]   queue_13_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_27 = {queue_13_enq_bits_lsWholeReg, queue_13_enq_bits_vs1};
  wire         queue_13_enq_bits_store;
  wire         queue_13_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_27 = {queue_13_enq_bits_store, queue_13_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_41 = {queue_dataIn_hi_lo_hi_27, queue_dataIn_hi_lo_lo_27};
  wire         queue_13_enq_bits_loadStore;
  wire         queue_13_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_27 = {queue_13_enq_bits_loadStore, queue_13_enq_bits_issueInst};
  wire [2:0]   queue_13_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_27 = {queue_13_enq_bits_instructionIndex, queue_dataIn_hi_40, queue_dataIn_lo_40};
  wire [60:0]  queue_dataIn_hi_hi_41 = {queue_dataIn_hi_hi_hi_27, queue_dataIn_hi_hi_lo_27};
  wire [68:0]  queue_dataIn_hi_41 = {queue_dataIn_hi_hi_41, queue_dataIn_hi_lo_41};
  wire [149:0] queue_dataIn_13 = {queue_dataIn_hi_41, queue_dataIn_lo_41};
  wire         queue_dataOut_13_csrInterface_vma = _queue_fifo_13_data_out[0];
  wire         queue_dataOut_13_csrInterface_vta = _queue_fifo_13_data_out[1];
  wire [1:0]   queue_dataOut_13_csrInterface_vxrm = _queue_fifo_13_data_out[3:2];
  wire [1:0]   queue_dataOut_13_csrInterface_vSew = _queue_fifo_13_data_out[5:4];
  wire [2:0]   queue_dataOut_13_csrInterface_vlmul = _queue_fifo_13_data_out[8:6];
  wire [11:0]  queue_dataOut_13_csrInterface_vStart = _queue_fifo_13_data_out[20:9];
  wire [11:0]  queue_dataOut_13_csrInterface_vl = _queue_fifo_13_data_out[32:21];
  wire [31:0]  queue_dataOut_13_readFromScalar = _queue_fifo_13_data_out[64:33];
  wire [2:0]   queue_dataOut_13_segment = _queue_fifo_13_data_out[67:65];
  wire         queue_dataOut_13_mask = _queue_fifo_13_data_out[68];
  wire [1:0]   queue_dataOut_13_loadStoreEEW = _queue_fifo_13_data_out[70:69];
  wire [4:0]   queue_dataOut_13_vd = _queue_fifo_13_data_out[75:71];
  wire [4:0]   queue_dataOut_13_vs2 = _queue_fifo_13_data_out[80:76];
  wire [4:0]   queue_dataOut_13_vs1 = _queue_fifo_13_data_out[85:81];
  wire         queue_dataOut_13_lsWholeReg = _queue_fifo_13_data_out[86];
  wire         queue_dataOut_13_special = _queue_fifo_13_data_out[87];
  wire         queue_dataOut_13_store = _queue_fifo_13_data_out[88];
  wire         queue_dataOut_13_issueInst = _queue_fifo_13_data_out[89];
  wire         queue_dataOut_13_loadStore = _queue_fifo_13_data_out[90];
  wire         queue_dataOut_13_decodeResult_logic = _queue_fifo_13_data_out[91];
  wire         queue_dataOut_13_decodeResult_adder = _queue_fifo_13_data_out[92];
  wire         queue_dataOut_13_decodeResult_shift = _queue_fifo_13_data_out[93];
  wire         queue_dataOut_13_decodeResult_multiplier = _queue_fifo_13_data_out[94];
  wire         queue_dataOut_13_decodeResult_divider = _queue_fifo_13_data_out[95];
  wire         queue_dataOut_13_decodeResult_multiCycle = _queue_fifo_13_data_out[96];
  wire         queue_dataOut_13_decodeResult_other = _queue_fifo_13_data_out[97];
  wire         queue_dataOut_13_decodeResult_unsigned0 = _queue_fifo_13_data_out[98];
  wire         queue_dataOut_13_decodeResult_unsigned1 = _queue_fifo_13_data_out[99];
  wire         queue_dataOut_13_decodeResult_itype = _queue_fifo_13_data_out[100];
  wire         queue_dataOut_13_decodeResult_nr = _queue_fifo_13_data_out[101];
  wire         queue_dataOut_13_decodeResult_red = _queue_fifo_13_data_out[102];
  wire         queue_dataOut_13_decodeResult_widenReduce = _queue_fifo_13_data_out[103];
  wire         queue_dataOut_13_decodeResult_targetRd = _queue_fifo_13_data_out[104];
  wire         queue_dataOut_13_decodeResult_slid = _queue_fifo_13_data_out[105];
  wire         queue_dataOut_13_decodeResult_gather = _queue_fifo_13_data_out[106];
  wire         queue_dataOut_13_decodeResult_gather16 = _queue_fifo_13_data_out[107];
  wire         queue_dataOut_13_decodeResult_compress = _queue_fifo_13_data_out[108];
  wire         queue_dataOut_13_decodeResult_unOrderWrite = _queue_fifo_13_data_out[109];
  wire         queue_dataOut_13_decodeResult_extend = _queue_fifo_13_data_out[110];
  wire         queue_dataOut_13_decodeResult_mv = _queue_fifo_13_data_out[111];
  wire         queue_dataOut_13_decodeResult_iota = _queue_fifo_13_data_out[112];
  wire [3:0]   queue_dataOut_13_decodeResult_uop = _queue_fifo_13_data_out[116:113];
  wire         queue_dataOut_13_decodeResult_maskLogic = _queue_fifo_13_data_out[117];
  wire         queue_dataOut_13_decodeResult_maskDestination = _queue_fifo_13_data_out[118];
  wire         queue_dataOut_13_decodeResult_maskSource = _queue_fifo_13_data_out[119];
  wire         queue_dataOut_13_decodeResult_readOnly = _queue_fifo_13_data_out[120];
  wire         queue_dataOut_13_decodeResult_vwmacc = _queue_fifo_13_data_out[121];
  wire         queue_dataOut_13_decodeResult_saturate = _queue_fifo_13_data_out[122];
  wire         queue_dataOut_13_decodeResult_special = _queue_fifo_13_data_out[123];
  wire         queue_dataOut_13_decodeResult_maskUnit = _queue_fifo_13_data_out[124];
  wire         queue_dataOut_13_decodeResult_crossWrite = _queue_fifo_13_data_out[125];
  wire         queue_dataOut_13_decodeResult_crossRead = _queue_fifo_13_data_out[126];
  wire         queue_dataOut_13_decodeResult_sWrite = _queue_fifo_13_data_out[127];
  wire         queue_dataOut_13_decodeResult_vtype = _queue_fifo_13_data_out[128];
  wire         queue_dataOut_13_decodeResult_sReadVD = _queue_fifo_13_data_out[129];
  wire         queue_dataOut_13_decodeResult_scheduler = _queue_fifo_13_data_out[130];
  wire         queue_dataOut_13_decodeResult_dontNeedExecuteInLane = _queue_fifo_13_data_out[131];
  wire         queue_dataOut_13_decodeResult_reverse = _queue_fifo_13_data_out[132];
  wire         queue_dataOut_13_decodeResult_average = _queue_fifo_13_data_out[133];
  wire         queue_dataOut_13_decodeResult_ffo = _queue_fifo_13_data_out[134];
  wire         queue_dataOut_13_decodeResult_popCount = _queue_fifo_13_data_out[135];
  wire [4:0]   queue_dataOut_13_decodeResult_topUop = _queue_fifo_13_data_out[140:136];
  wire         queue_dataOut_13_decodeResult_specialSlot = _queue_fifo_13_data_out[141];
  wire         queue_dataOut_13_decodeResult_float = _queue_fifo_13_data_out[142];
  wire [1:0]   queue_dataOut_13_decodeResult_fpExecutionType = _queue_fifo_13_data_out[144:143];
  wire         queue_dataOut_13_decodeResult_floatMul = _queue_fifo_13_data_out[145];
  wire         queue_dataOut_13_decodeResult_orderReduce = _queue_fifo_13_data_out[146];
  wire [2:0]   queue_dataOut_13_instructionIndex = _queue_fifo_13_data_out[149:147];
  wire         queue_13_enq_ready = ~_queue_fifo_13_full;
  wire         queue_13_enq_valid;
  assign queue_13_deq_valid = ~_queue_fifo_13_empty | queue_13_enq_valid;
  assign queue_13_deq_bits_instructionIndex = _queue_fifo_13_empty ? queue_13_enq_bits_instructionIndex : queue_dataOut_13_instructionIndex;
  assign queue_13_deq_bits_decodeResult_orderReduce = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_orderReduce : queue_dataOut_13_decodeResult_orderReduce;
  assign queue_13_deq_bits_decodeResult_floatMul = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_floatMul : queue_dataOut_13_decodeResult_floatMul;
  assign queue_13_deq_bits_decodeResult_fpExecutionType = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_fpExecutionType : queue_dataOut_13_decodeResult_fpExecutionType;
  assign queue_13_deq_bits_decodeResult_float = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_float : queue_dataOut_13_decodeResult_float;
  assign queue_13_deq_bits_decodeResult_specialSlot = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_specialSlot : queue_dataOut_13_decodeResult_specialSlot;
  assign queue_13_deq_bits_decodeResult_topUop = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_topUop : queue_dataOut_13_decodeResult_topUop;
  assign queue_13_deq_bits_decodeResult_popCount = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_popCount : queue_dataOut_13_decodeResult_popCount;
  assign queue_13_deq_bits_decodeResult_ffo = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_ffo : queue_dataOut_13_decodeResult_ffo;
  assign queue_13_deq_bits_decodeResult_average = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_average : queue_dataOut_13_decodeResult_average;
  assign queue_13_deq_bits_decodeResult_reverse = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_reverse : queue_dataOut_13_decodeResult_reverse;
  assign queue_13_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_13_decodeResult_dontNeedExecuteInLane;
  assign queue_13_deq_bits_decodeResult_scheduler = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_scheduler : queue_dataOut_13_decodeResult_scheduler;
  assign queue_13_deq_bits_decodeResult_sReadVD = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_sReadVD : queue_dataOut_13_decodeResult_sReadVD;
  assign queue_13_deq_bits_decodeResult_vtype = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_vtype : queue_dataOut_13_decodeResult_vtype;
  assign queue_13_deq_bits_decodeResult_sWrite = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_sWrite : queue_dataOut_13_decodeResult_sWrite;
  assign queue_13_deq_bits_decodeResult_crossRead = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_crossRead : queue_dataOut_13_decodeResult_crossRead;
  assign queue_13_deq_bits_decodeResult_crossWrite = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_crossWrite : queue_dataOut_13_decodeResult_crossWrite;
  assign queue_13_deq_bits_decodeResult_maskUnit = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_maskUnit : queue_dataOut_13_decodeResult_maskUnit;
  assign queue_13_deq_bits_decodeResult_special = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_special : queue_dataOut_13_decodeResult_special;
  assign queue_13_deq_bits_decodeResult_saturate = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_saturate : queue_dataOut_13_decodeResult_saturate;
  assign queue_13_deq_bits_decodeResult_vwmacc = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_vwmacc : queue_dataOut_13_decodeResult_vwmacc;
  assign queue_13_deq_bits_decodeResult_readOnly = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_readOnly : queue_dataOut_13_decodeResult_readOnly;
  assign queue_13_deq_bits_decodeResult_maskSource = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_maskSource : queue_dataOut_13_decodeResult_maskSource;
  assign queue_13_deq_bits_decodeResult_maskDestination = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_maskDestination : queue_dataOut_13_decodeResult_maskDestination;
  assign queue_13_deq_bits_decodeResult_maskLogic = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_maskLogic : queue_dataOut_13_decodeResult_maskLogic;
  assign queue_13_deq_bits_decodeResult_uop = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_uop : queue_dataOut_13_decodeResult_uop;
  assign queue_13_deq_bits_decodeResult_iota = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_iota : queue_dataOut_13_decodeResult_iota;
  assign queue_13_deq_bits_decodeResult_mv = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_mv : queue_dataOut_13_decodeResult_mv;
  assign queue_13_deq_bits_decodeResult_extend = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_extend : queue_dataOut_13_decodeResult_extend;
  assign queue_13_deq_bits_decodeResult_unOrderWrite = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_unOrderWrite : queue_dataOut_13_decodeResult_unOrderWrite;
  assign queue_13_deq_bits_decodeResult_compress = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_compress : queue_dataOut_13_decodeResult_compress;
  assign queue_13_deq_bits_decodeResult_gather16 = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_gather16 : queue_dataOut_13_decodeResult_gather16;
  assign queue_13_deq_bits_decodeResult_gather = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_gather : queue_dataOut_13_decodeResult_gather;
  assign queue_13_deq_bits_decodeResult_slid = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_slid : queue_dataOut_13_decodeResult_slid;
  assign queue_13_deq_bits_decodeResult_targetRd = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_targetRd : queue_dataOut_13_decodeResult_targetRd;
  assign queue_13_deq_bits_decodeResult_widenReduce = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_widenReduce : queue_dataOut_13_decodeResult_widenReduce;
  assign queue_13_deq_bits_decodeResult_red = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_red : queue_dataOut_13_decodeResult_red;
  assign queue_13_deq_bits_decodeResult_nr = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_nr : queue_dataOut_13_decodeResult_nr;
  assign queue_13_deq_bits_decodeResult_itype = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_itype : queue_dataOut_13_decodeResult_itype;
  assign queue_13_deq_bits_decodeResult_unsigned1 = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_unsigned1 : queue_dataOut_13_decodeResult_unsigned1;
  assign queue_13_deq_bits_decodeResult_unsigned0 = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_unsigned0 : queue_dataOut_13_decodeResult_unsigned0;
  assign queue_13_deq_bits_decodeResult_other = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_other : queue_dataOut_13_decodeResult_other;
  assign queue_13_deq_bits_decodeResult_multiCycle = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_multiCycle : queue_dataOut_13_decodeResult_multiCycle;
  assign queue_13_deq_bits_decodeResult_divider = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_divider : queue_dataOut_13_decodeResult_divider;
  assign queue_13_deq_bits_decodeResult_multiplier = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_multiplier : queue_dataOut_13_decodeResult_multiplier;
  assign queue_13_deq_bits_decodeResult_shift = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_shift : queue_dataOut_13_decodeResult_shift;
  assign queue_13_deq_bits_decodeResult_adder = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_adder : queue_dataOut_13_decodeResult_adder;
  assign queue_13_deq_bits_decodeResult_logic = _queue_fifo_13_empty ? queue_13_enq_bits_decodeResult_logic : queue_dataOut_13_decodeResult_logic;
  assign queue_13_deq_bits_loadStore = _queue_fifo_13_empty ? queue_13_enq_bits_loadStore : queue_dataOut_13_loadStore;
  assign queue_13_deq_bits_issueInst = _queue_fifo_13_empty ? queue_13_enq_bits_issueInst : queue_dataOut_13_issueInst;
  assign queue_13_deq_bits_store = _queue_fifo_13_empty ? queue_13_enq_bits_store : queue_dataOut_13_store;
  assign queue_13_deq_bits_special = _queue_fifo_13_empty ? queue_13_enq_bits_special : queue_dataOut_13_special;
  assign queue_13_deq_bits_lsWholeReg = _queue_fifo_13_empty ? queue_13_enq_bits_lsWholeReg : queue_dataOut_13_lsWholeReg;
  assign queue_13_deq_bits_vs1 = _queue_fifo_13_empty ? queue_13_enq_bits_vs1 : queue_dataOut_13_vs1;
  assign queue_13_deq_bits_vs2 = _queue_fifo_13_empty ? queue_13_enq_bits_vs2 : queue_dataOut_13_vs2;
  assign queue_13_deq_bits_vd = _queue_fifo_13_empty ? queue_13_enq_bits_vd : queue_dataOut_13_vd;
  assign queue_13_deq_bits_loadStoreEEW = _queue_fifo_13_empty ? queue_13_enq_bits_loadStoreEEW : queue_dataOut_13_loadStoreEEW;
  assign queue_13_deq_bits_mask = _queue_fifo_13_empty ? queue_13_enq_bits_mask : queue_dataOut_13_mask;
  assign queue_13_deq_bits_segment = _queue_fifo_13_empty ? queue_13_enq_bits_segment : queue_dataOut_13_segment;
  assign queue_13_deq_bits_readFromScalar = _queue_fifo_13_empty ? queue_13_enq_bits_readFromScalar : queue_dataOut_13_readFromScalar;
  assign queue_13_deq_bits_csrInterface_vl = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vl : queue_dataOut_13_csrInterface_vl;
  assign queue_13_deq_bits_csrInterface_vStart = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vStart : queue_dataOut_13_csrInterface_vStart;
  assign queue_13_deq_bits_csrInterface_vlmul = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vlmul : queue_dataOut_13_csrInterface_vlmul;
  assign queue_13_deq_bits_csrInterface_vSew = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vSew : queue_dataOut_13_csrInterface_vSew;
  assign queue_13_deq_bits_csrInterface_vxrm = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vxrm : queue_dataOut_13_csrInterface_vxrm;
  assign queue_13_deq_bits_csrInterface_vta = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vta : queue_dataOut_13_csrInterface_vta;
  assign queue_13_deq_bits_csrInterface_vma = _queue_fifo_13_empty ? queue_13_enq_bits_csrInterface_vma : queue_dataOut_13_csrInterface_vma;
  wire         laneVec_13_laneRequest_bits_issueInst = laneRequestSinkWire_13_ready & laneRequestSinkWire_13_valid;
  reg          releasePipe_pipe_v_13;
  wire         releasePipe_pipe_out_13_valid = releasePipe_pipe_v_13;
  wire         laneRequestSourceWire_13_ready;
  wire         validSource_13_valid = laneRequestSourceWire_13_ready & laneRequestSourceWire_13_valid;
  reg  [2:0]   tokenCheck_counter_13;
  wire [2:0]   tokenCheck_counterChange_13 = validSource_13_valid ? 3'h1 : 3'h7;
  assign tokenCheck_13 = ~(tokenCheck_counter_13[2]);
  assign laneRequestSourceWire_13_ready = tokenCheck_13;
  assign queue_13_enq_valid = validSink_13_valid;
  assign queue_13_enq_bits_instructionIndex = validSink_13_bits_instructionIndex;
  assign queue_13_enq_bits_decodeResult_orderReduce = validSink_13_bits_decodeResult_orderReduce;
  assign queue_13_enq_bits_decodeResult_floatMul = validSink_13_bits_decodeResult_floatMul;
  assign queue_13_enq_bits_decodeResult_fpExecutionType = validSink_13_bits_decodeResult_fpExecutionType;
  assign queue_13_enq_bits_decodeResult_float = validSink_13_bits_decodeResult_float;
  assign queue_13_enq_bits_decodeResult_specialSlot = validSink_13_bits_decodeResult_specialSlot;
  assign queue_13_enq_bits_decodeResult_topUop = validSink_13_bits_decodeResult_topUop;
  assign queue_13_enq_bits_decodeResult_popCount = validSink_13_bits_decodeResult_popCount;
  assign queue_13_enq_bits_decodeResult_ffo = validSink_13_bits_decodeResult_ffo;
  assign queue_13_enq_bits_decodeResult_average = validSink_13_bits_decodeResult_average;
  assign queue_13_enq_bits_decodeResult_reverse = validSink_13_bits_decodeResult_reverse;
  assign queue_13_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_13_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_13_enq_bits_decodeResult_scheduler = validSink_13_bits_decodeResult_scheduler;
  assign queue_13_enq_bits_decodeResult_sReadVD = validSink_13_bits_decodeResult_sReadVD;
  assign queue_13_enq_bits_decodeResult_vtype = validSink_13_bits_decodeResult_vtype;
  assign queue_13_enq_bits_decodeResult_sWrite = validSink_13_bits_decodeResult_sWrite;
  assign queue_13_enq_bits_decodeResult_crossRead = validSink_13_bits_decodeResult_crossRead;
  assign queue_13_enq_bits_decodeResult_crossWrite = validSink_13_bits_decodeResult_crossWrite;
  assign queue_13_enq_bits_decodeResult_maskUnit = validSink_13_bits_decodeResult_maskUnit;
  assign queue_13_enq_bits_decodeResult_special = validSink_13_bits_decodeResult_special;
  assign queue_13_enq_bits_decodeResult_saturate = validSink_13_bits_decodeResult_saturate;
  assign queue_13_enq_bits_decodeResult_vwmacc = validSink_13_bits_decodeResult_vwmacc;
  assign queue_13_enq_bits_decodeResult_readOnly = validSink_13_bits_decodeResult_readOnly;
  assign queue_13_enq_bits_decodeResult_maskSource = validSink_13_bits_decodeResult_maskSource;
  assign queue_13_enq_bits_decodeResult_maskDestination = validSink_13_bits_decodeResult_maskDestination;
  assign queue_13_enq_bits_decodeResult_maskLogic = validSink_13_bits_decodeResult_maskLogic;
  assign queue_13_enq_bits_decodeResult_uop = validSink_13_bits_decodeResult_uop;
  assign queue_13_enq_bits_decodeResult_iota = validSink_13_bits_decodeResult_iota;
  assign queue_13_enq_bits_decodeResult_mv = validSink_13_bits_decodeResult_mv;
  assign queue_13_enq_bits_decodeResult_extend = validSink_13_bits_decodeResult_extend;
  assign queue_13_enq_bits_decodeResult_unOrderWrite = validSink_13_bits_decodeResult_unOrderWrite;
  assign queue_13_enq_bits_decodeResult_compress = validSink_13_bits_decodeResult_compress;
  assign queue_13_enq_bits_decodeResult_gather16 = validSink_13_bits_decodeResult_gather16;
  assign queue_13_enq_bits_decodeResult_gather = validSink_13_bits_decodeResult_gather;
  assign queue_13_enq_bits_decodeResult_slid = validSink_13_bits_decodeResult_slid;
  assign queue_13_enq_bits_decodeResult_targetRd = validSink_13_bits_decodeResult_targetRd;
  assign queue_13_enq_bits_decodeResult_widenReduce = validSink_13_bits_decodeResult_widenReduce;
  assign queue_13_enq_bits_decodeResult_red = validSink_13_bits_decodeResult_red;
  assign queue_13_enq_bits_decodeResult_nr = validSink_13_bits_decodeResult_nr;
  assign queue_13_enq_bits_decodeResult_itype = validSink_13_bits_decodeResult_itype;
  assign queue_13_enq_bits_decodeResult_unsigned1 = validSink_13_bits_decodeResult_unsigned1;
  assign queue_13_enq_bits_decodeResult_unsigned0 = validSink_13_bits_decodeResult_unsigned0;
  assign queue_13_enq_bits_decodeResult_other = validSink_13_bits_decodeResult_other;
  assign queue_13_enq_bits_decodeResult_multiCycle = validSink_13_bits_decodeResult_multiCycle;
  assign queue_13_enq_bits_decodeResult_divider = validSink_13_bits_decodeResult_divider;
  assign queue_13_enq_bits_decodeResult_multiplier = validSink_13_bits_decodeResult_multiplier;
  assign queue_13_enq_bits_decodeResult_shift = validSink_13_bits_decodeResult_shift;
  assign queue_13_enq_bits_decodeResult_adder = validSink_13_bits_decodeResult_adder;
  assign queue_13_enq_bits_decodeResult_logic = validSink_13_bits_decodeResult_logic;
  assign queue_13_enq_bits_loadStore = validSink_13_bits_loadStore;
  assign queue_13_enq_bits_issueInst = validSink_13_bits_issueInst;
  assign queue_13_enq_bits_store = validSink_13_bits_store;
  assign queue_13_enq_bits_special = validSink_13_bits_special;
  assign queue_13_enq_bits_lsWholeReg = validSink_13_bits_lsWholeReg;
  assign queue_13_enq_bits_vs1 = validSink_13_bits_vs1;
  assign queue_13_enq_bits_vs2 = validSink_13_bits_vs2;
  assign queue_13_enq_bits_vd = validSink_13_bits_vd;
  assign queue_13_enq_bits_loadStoreEEW = validSink_13_bits_loadStoreEEW;
  assign queue_13_enq_bits_mask = validSink_13_bits_mask;
  assign queue_13_enq_bits_segment = validSink_13_bits_segment;
  assign queue_13_enq_bits_readFromScalar = validSink_13_bits_readFromScalar;
  assign queue_13_enq_bits_csrInterface_vl = validSink_13_bits_csrInterface_vl;
  assign queue_13_enq_bits_csrInterface_vStart = validSink_13_bits_csrInterface_vStart;
  assign queue_13_enq_bits_csrInterface_vlmul = validSink_13_bits_csrInterface_vlmul;
  assign queue_13_enq_bits_csrInterface_vSew = validSink_13_bits_csrInterface_vSew;
  assign queue_13_enq_bits_csrInterface_vxrm = validSink_13_bits_csrInterface_vxrm;
  assign queue_13_enq_bits_csrInterface_vta = validSink_13_bits_csrInterface_vta;
  assign queue_13_enq_bits_csrInterface_vma = validSink_13_bits_csrInterface_vma;
  reg          shifterReg_13_0_valid;
  assign validSink_13_valid = shifterReg_13_0_valid;
  reg  [2:0]   shifterReg_13_0_bits_instructionIndex;
  assign validSink_13_bits_instructionIndex = shifterReg_13_0_bits_instructionIndex;
  reg          shifterReg_13_0_bits_decodeResult_orderReduce;
  assign validSink_13_bits_decodeResult_orderReduce = shifterReg_13_0_bits_decodeResult_orderReduce;
  reg          shifterReg_13_0_bits_decodeResult_floatMul;
  assign validSink_13_bits_decodeResult_floatMul = shifterReg_13_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_13_0_bits_decodeResult_fpExecutionType;
  assign validSink_13_bits_decodeResult_fpExecutionType = shifterReg_13_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_13_0_bits_decodeResult_float;
  assign validSink_13_bits_decodeResult_float = shifterReg_13_0_bits_decodeResult_float;
  reg          shifterReg_13_0_bits_decodeResult_specialSlot;
  assign validSink_13_bits_decodeResult_specialSlot = shifterReg_13_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_13_0_bits_decodeResult_topUop;
  assign validSink_13_bits_decodeResult_topUop = shifterReg_13_0_bits_decodeResult_topUop;
  reg          shifterReg_13_0_bits_decodeResult_popCount;
  assign validSink_13_bits_decodeResult_popCount = shifterReg_13_0_bits_decodeResult_popCount;
  reg          shifterReg_13_0_bits_decodeResult_ffo;
  assign validSink_13_bits_decodeResult_ffo = shifterReg_13_0_bits_decodeResult_ffo;
  reg          shifterReg_13_0_bits_decodeResult_average;
  assign validSink_13_bits_decodeResult_average = shifterReg_13_0_bits_decodeResult_average;
  reg          shifterReg_13_0_bits_decodeResult_reverse;
  assign validSink_13_bits_decodeResult_reverse = shifterReg_13_0_bits_decodeResult_reverse;
  reg          shifterReg_13_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_13_bits_decodeResult_dontNeedExecuteInLane = shifterReg_13_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_13_0_bits_decodeResult_scheduler;
  assign validSink_13_bits_decodeResult_scheduler = shifterReg_13_0_bits_decodeResult_scheduler;
  reg          shifterReg_13_0_bits_decodeResult_sReadVD;
  assign validSink_13_bits_decodeResult_sReadVD = shifterReg_13_0_bits_decodeResult_sReadVD;
  reg          shifterReg_13_0_bits_decodeResult_vtype;
  assign validSink_13_bits_decodeResult_vtype = shifterReg_13_0_bits_decodeResult_vtype;
  reg          shifterReg_13_0_bits_decodeResult_sWrite;
  assign validSink_13_bits_decodeResult_sWrite = shifterReg_13_0_bits_decodeResult_sWrite;
  reg          shifterReg_13_0_bits_decodeResult_crossRead;
  assign validSink_13_bits_decodeResult_crossRead = shifterReg_13_0_bits_decodeResult_crossRead;
  reg          shifterReg_13_0_bits_decodeResult_crossWrite;
  assign validSink_13_bits_decodeResult_crossWrite = shifterReg_13_0_bits_decodeResult_crossWrite;
  reg          shifterReg_13_0_bits_decodeResult_maskUnit;
  assign validSink_13_bits_decodeResult_maskUnit = shifterReg_13_0_bits_decodeResult_maskUnit;
  reg          shifterReg_13_0_bits_decodeResult_special;
  assign validSink_13_bits_decodeResult_special = shifterReg_13_0_bits_decodeResult_special;
  reg          shifterReg_13_0_bits_decodeResult_saturate;
  assign validSink_13_bits_decodeResult_saturate = shifterReg_13_0_bits_decodeResult_saturate;
  reg          shifterReg_13_0_bits_decodeResult_vwmacc;
  assign validSink_13_bits_decodeResult_vwmacc = shifterReg_13_0_bits_decodeResult_vwmacc;
  reg          shifterReg_13_0_bits_decodeResult_readOnly;
  assign validSink_13_bits_decodeResult_readOnly = shifterReg_13_0_bits_decodeResult_readOnly;
  reg          shifterReg_13_0_bits_decodeResult_maskSource;
  assign validSink_13_bits_decodeResult_maskSource = shifterReg_13_0_bits_decodeResult_maskSource;
  reg          shifterReg_13_0_bits_decodeResult_maskDestination;
  assign validSink_13_bits_decodeResult_maskDestination = shifterReg_13_0_bits_decodeResult_maskDestination;
  reg          shifterReg_13_0_bits_decodeResult_maskLogic;
  assign validSink_13_bits_decodeResult_maskLogic = shifterReg_13_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_13_0_bits_decodeResult_uop;
  assign validSink_13_bits_decodeResult_uop = shifterReg_13_0_bits_decodeResult_uop;
  reg          shifterReg_13_0_bits_decodeResult_iota;
  assign validSink_13_bits_decodeResult_iota = shifterReg_13_0_bits_decodeResult_iota;
  reg          shifterReg_13_0_bits_decodeResult_mv;
  assign validSink_13_bits_decodeResult_mv = shifterReg_13_0_bits_decodeResult_mv;
  reg          shifterReg_13_0_bits_decodeResult_extend;
  assign validSink_13_bits_decodeResult_extend = shifterReg_13_0_bits_decodeResult_extend;
  reg          shifterReg_13_0_bits_decodeResult_unOrderWrite;
  assign validSink_13_bits_decodeResult_unOrderWrite = shifterReg_13_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_13_0_bits_decodeResult_compress;
  assign validSink_13_bits_decodeResult_compress = shifterReg_13_0_bits_decodeResult_compress;
  reg          shifterReg_13_0_bits_decodeResult_gather16;
  assign validSink_13_bits_decodeResult_gather16 = shifterReg_13_0_bits_decodeResult_gather16;
  reg          shifterReg_13_0_bits_decodeResult_gather;
  assign validSink_13_bits_decodeResult_gather = shifterReg_13_0_bits_decodeResult_gather;
  reg          shifterReg_13_0_bits_decodeResult_slid;
  assign validSink_13_bits_decodeResult_slid = shifterReg_13_0_bits_decodeResult_slid;
  reg          shifterReg_13_0_bits_decodeResult_targetRd;
  assign validSink_13_bits_decodeResult_targetRd = shifterReg_13_0_bits_decodeResult_targetRd;
  reg          shifterReg_13_0_bits_decodeResult_widenReduce;
  assign validSink_13_bits_decodeResult_widenReduce = shifterReg_13_0_bits_decodeResult_widenReduce;
  reg          shifterReg_13_0_bits_decodeResult_red;
  assign validSink_13_bits_decodeResult_red = shifterReg_13_0_bits_decodeResult_red;
  reg          shifterReg_13_0_bits_decodeResult_nr;
  assign validSink_13_bits_decodeResult_nr = shifterReg_13_0_bits_decodeResult_nr;
  reg          shifterReg_13_0_bits_decodeResult_itype;
  assign validSink_13_bits_decodeResult_itype = shifterReg_13_0_bits_decodeResult_itype;
  reg          shifterReg_13_0_bits_decodeResult_unsigned1;
  assign validSink_13_bits_decodeResult_unsigned1 = shifterReg_13_0_bits_decodeResult_unsigned1;
  reg          shifterReg_13_0_bits_decodeResult_unsigned0;
  assign validSink_13_bits_decodeResult_unsigned0 = shifterReg_13_0_bits_decodeResult_unsigned0;
  reg          shifterReg_13_0_bits_decodeResult_other;
  assign validSink_13_bits_decodeResult_other = shifterReg_13_0_bits_decodeResult_other;
  reg          shifterReg_13_0_bits_decodeResult_multiCycle;
  assign validSink_13_bits_decodeResult_multiCycle = shifterReg_13_0_bits_decodeResult_multiCycle;
  reg          shifterReg_13_0_bits_decodeResult_divider;
  assign validSink_13_bits_decodeResult_divider = shifterReg_13_0_bits_decodeResult_divider;
  reg          shifterReg_13_0_bits_decodeResult_multiplier;
  assign validSink_13_bits_decodeResult_multiplier = shifterReg_13_0_bits_decodeResult_multiplier;
  reg          shifterReg_13_0_bits_decodeResult_shift;
  assign validSink_13_bits_decodeResult_shift = shifterReg_13_0_bits_decodeResult_shift;
  reg          shifterReg_13_0_bits_decodeResult_adder;
  assign validSink_13_bits_decodeResult_adder = shifterReg_13_0_bits_decodeResult_adder;
  reg          shifterReg_13_0_bits_decodeResult_logic;
  assign validSink_13_bits_decodeResult_logic = shifterReg_13_0_bits_decodeResult_logic;
  reg          shifterReg_13_0_bits_loadStore;
  assign validSink_13_bits_loadStore = shifterReg_13_0_bits_loadStore;
  reg          shifterReg_13_0_bits_issueInst;
  assign validSink_13_bits_issueInst = shifterReg_13_0_bits_issueInst;
  reg          shifterReg_13_0_bits_store;
  assign validSink_13_bits_store = shifterReg_13_0_bits_store;
  reg          shifterReg_13_0_bits_special;
  assign validSink_13_bits_special = shifterReg_13_0_bits_special;
  reg          shifterReg_13_0_bits_lsWholeReg;
  assign validSink_13_bits_lsWholeReg = shifterReg_13_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_13_0_bits_vs1;
  assign validSink_13_bits_vs1 = shifterReg_13_0_bits_vs1;
  reg  [4:0]   shifterReg_13_0_bits_vs2;
  assign validSink_13_bits_vs2 = shifterReg_13_0_bits_vs2;
  reg  [4:0]   shifterReg_13_0_bits_vd;
  assign validSink_13_bits_vd = shifterReg_13_0_bits_vd;
  reg  [1:0]   shifterReg_13_0_bits_loadStoreEEW;
  assign validSink_13_bits_loadStoreEEW = shifterReg_13_0_bits_loadStoreEEW;
  reg          shifterReg_13_0_bits_mask;
  assign validSink_13_bits_mask = shifterReg_13_0_bits_mask;
  reg  [2:0]   shifterReg_13_0_bits_segment;
  assign validSink_13_bits_segment = shifterReg_13_0_bits_segment;
  reg  [31:0]  shifterReg_13_0_bits_readFromScalar;
  assign validSink_13_bits_readFromScalar = shifterReg_13_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_13_0_bits_csrInterface_vl;
  assign validSink_13_bits_csrInterface_vl = shifterReg_13_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_13_0_bits_csrInterface_vStart;
  assign validSink_13_bits_csrInterface_vStart = shifterReg_13_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_13_0_bits_csrInterface_vlmul;
  assign validSink_13_bits_csrInterface_vlmul = shifterReg_13_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_13_0_bits_csrInterface_vSew;
  assign validSink_13_bits_csrInterface_vSew = shifterReg_13_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_13_0_bits_csrInterface_vxrm;
  assign validSink_13_bits_csrInterface_vxrm = shifterReg_13_0_bits_csrInterface_vxrm;
  reg          shifterReg_13_0_bits_csrInterface_vta;
  assign validSink_13_bits_csrInterface_vta = shifterReg_13_0_bits_csrInterface_vta;
  reg          shifterReg_13_0_bits_csrInterface_vma;
  assign validSink_13_bits_csrInterface_vma = shifterReg_13_0_bits_csrInterface_vma;
  wire         shifterValid_13 = shifterReg_13_0_valid | validSource_13_valid;
  wire         validSink_14_valid;
  wire [2:0]   validSink_14_bits_instructionIndex;
  wire         validSink_14_bits_decodeResult_orderReduce;
  wire         validSink_14_bits_decodeResult_floatMul;
  wire [1:0]   validSink_14_bits_decodeResult_fpExecutionType;
  wire         validSink_14_bits_decodeResult_float;
  wire         validSink_14_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_14_bits_decodeResult_topUop;
  wire         validSink_14_bits_decodeResult_popCount;
  wire         validSink_14_bits_decodeResult_ffo;
  wire         validSink_14_bits_decodeResult_average;
  wire         validSink_14_bits_decodeResult_reverse;
  wire         validSink_14_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_14_bits_decodeResult_scheduler;
  wire         validSink_14_bits_decodeResult_sReadVD;
  wire         validSink_14_bits_decodeResult_vtype;
  wire         validSink_14_bits_decodeResult_sWrite;
  wire         validSink_14_bits_decodeResult_crossRead;
  wire         validSink_14_bits_decodeResult_crossWrite;
  wire         validSink_14_bits_decodeResult_maskUnit;
  wire         validSink_14_bits_decodeResult_special;
  wire         validSink_14_bits_decodeResult_saturate;
  wire         validSink_14_bits_decodeResult_vwmacc;
  wire         validSink_14_bits_decodeResult_readOnly;
  wire         validSink_14_bits_decodeResult_maskSource;
  wire         validSink_14_bits_decodeResult_maskDestination;
  wire         validSink_14_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_14_bits_decodeResult_uop;
  wire         validSink_14_bits_decodeResult_iota;
  wire         validSink_14_bits_decodeResult_mv;
  wire         validSink_14_bits_decodeResult_extend;
  wire         validSink_14_bits_decodeResult_unOrderWrite;
  wire         validSink_14_bits_decodeResult_compress;
  wire         validSink_14_bits_decodeResult_gather16;
  wire         validSink_14_bits_decodeResult_gather;
  wire         validSink_14_bits_decodeResult_slid;
  wire         validSink_14_bits_decodeResult_targetRd;
  wire         validSink_14_bits_decodeResult_widenReduce;
  wire         validSink_14_bits_decodeResult_red;
  wire         validSink_14_bits_decodeResult_nr;
  wire         validSink_14_bits_decodeResult_itype;
  wire         validSink_14_bits_decodeResult_unsigned1;
  wire         validSink_14_bits_decodeResult_unsigned0;
  wire         validSink_14_bits_decodeResult_other;
  wire         validSink_14_bits_decodeResult_multiCycle;
  wire         validSink_14_bits_decodeResult_divider;
  wire         validSink_14_bits_decodeResult_multiplier;
  wire         validSink_14_bits_decodeResult_shift;
  wire         validSink_14_bits_decodeResult_adder;
  wire         validSink_14_bits_decodeResult_logic;
  wire         validSink_14_bits_loadStore;
  wire         validSink_14_bits_issueInst;
  wire         validSink_14_bits_store;
  wire         validSink_14_bits_special;
  wire         validSink_14_bits_lsWholeReg;
  wire [4:0]   validSink_14_bits_vs1;
  wire [4:0]   validSink_14_bits_vs2;
  wire [4:0]   validSink_14_bits_vd;
  wire [1:0]   validSink_14_bits_loadStoreEEW;
  wire         validSink_14_bits_mask;
  wire [2:0]   validSink_14_bits_segment;
  wire [31:0]  validSink_14_bits_readFromScalar;
  wire [11:0]  validSink_14_bits_csrInterface_vl;
  wire [11:0]  validSink_14_bits_csrInterface_vStart;
  wire [2:0]   validSink_14_bits_csrInterface_vlmul;
  wire [1:0]   validSink_14_bits_csrInterface_vSew;
  wire [1:0]   validSink_14_bits_csrInterface_vxrm;
  wire         validSink_14_bits_csrInterface_vta;
  wire         validSink_14_bits_csrInterface_vma;
  wire         laneRequestSinkWire_14_valid = queue_14_deq_valid;
  wire [2:0]   laneRequestSinkWire_14_bits_instructionIndex = queue_14_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_14_bits_decodeResult_orderReduce = queue_14_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_14_bits_decodeResult_floatMul = queue_14_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_14_bits_decodeResult_fpExecutionType = queue_14_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_14_bits_decodeResult_float = queue_14_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_14_bits_decodeResult_specialSlot = queue_14_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_14_bits_decodeResult_topUop = queue_14_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_14_bits_decodeResult_popCount = queue_14_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_14_bits_decodeResult_ffo = queue_14_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_14_bits_decodeResult_average = queue_14_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_14_bits_decodeResult_reverse = queue_14_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_14_bits_decodeResult_dontNeedExecuteInLane = queue_14_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_14_bits_decodeResult_scheduler = queue_14_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_14_bits_decodeResult_sReadVD = queue_14_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_14_bits_decodeResult_vtype = queue_14_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_14_bits_decodeResult_sWrite = queue_14_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_14_bits_decodeResult_crossRead = queue_14_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_14_bits_decodeResult_crossWrite = queue_14_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_14_bits_decodeResult_maskUnit = queue_14_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_14_bits_decodeResult_special = queue_14_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_14_bits_decodeResult_saturate = queue_14_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_14_bits_decodeResult_vwmacc = queue_14_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_14_bits_decodeResult_readOnly = queue_14_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_14_bits_decodeResult_maskSource = queue_14_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_14_bits_decodeResult_maskDestination = queue_14_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_14_bits_decodeResult_maskLogic = queue_14_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_14_bits_decodeResult_uop = queue_14_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_14_bits_decodeResult_iota = queue_14_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_14_bits_decodeResult_mv = queue_14_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_14_bits_decodeResult_extend = queue_14_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_14_bits_decodeResult_unOrderWrite = queue_14_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_14_bits_decodeResult_compress = queue_14_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_14_bits_decodeResult_gather16 = queue_14_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_14_bits_decodeResult_gather = queue_14_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_14_bits_decodeResult_slid = queue_14_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_14_bits_decodeResult_targetRd = queue_14_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_14_bits_decodeResult_widenReduce = queue_14_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_14_bits_decodeResult_red = queue_14_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_14_bits_decodeResult_nr = queue_14_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_14_bits_decodeResult_itype = queue_14_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_14_bits_decodeResult_unsigned1 = queue_14_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_14_bits_decodeResult_unsigned0 = queue_14_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_14_bits_decodeResult_other = queue_14_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_14_bits_decodeResult_multiCycle = queue_14_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_14_bits_decodeResult_divider = queue_14_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_14_bits_decodeResult_multiplier = queue_14_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_14_bits_decodeResult_shift = queue_14_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_14_bits_decodeResult_adder = queue_14_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_14_bits_decodeResult_logic = queue_14_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_14_bits_loadStore = queue_14_deq_bits_loadStore;
  wire         laneRequestSinkWire_14_bits_issueInst = queue_14_deq_bits_issueInst;
  wire         laneRequestSinkWire_14_bits_store = queue_14_deq_bits_store;
  wire         laneRequestSinkWire_14_bits_special = queue_14_deq_bits_special;
  wire         laneRequestSinkWire_14_bits_lsWholeReg = queue_14_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_14_bits_vs1 = queue_14_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_14_bits_vs2 = queue_14_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_14_bits_vd = queue_14_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_14_bits_loadStoreEEW = queue_14_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_14_bits_mask = queue_14_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_14_bits_segment = queue_14_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_14_bits_readFromScalar = queue_14_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_14_bits_csrInterface_vl = queue_14_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_14_bits_csrInterface_vStart = queue_14_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_14_bits_csrInterface_vlmul = queue_14_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_14_bits_csrInterface_vSew = queue_14_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_14_bits_csrInterface_vxrm = queue_14_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_14_bits_csrInterface_vta = queue_14_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_14_bits_csrInterface_vma = queue_14_deq_bits_csrInterface_vma;
  wire [1:0]   queue_14_enq_bits_csrInterface_vxrm;
  wire         queue_14_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_42 = {queue_14_enq_bits_csrInterface_vxrm, queue_14_enq_bits_csrInterface_vta};
  wire         queue_14_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_42 = {queue_dataIn_lo_hi_42, queue_14_enq_bits_csrInterface_vma};
  wire [2:0]   queue_14_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_14_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_42 = {queue_14_enq_bits_csrInterface_vlmul, queue_14_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_14_enq_bits_csrInterface_vl;
  wire [11:0]  queue_14_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_42 = {queue_14_enq_bits_csrInterface_vl, queue_14_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_42 = {queue_dataIn_hi_hi_42, queue_dataIn_hi_lo_42};
  wire         queue_14_enq_bits_decodeResult_shift;
  wire         queue_14_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_14 = {queue_14_enq_bits_decodeResult_shift, queue_14_enq_bits_decodeResult_adder};
  wire         queue_14_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_14 = {queue_dataIn_lo_lo_lo_lo_hi_14, queue_14_enq_bits_decodeResult_logic};
  wire         queue_14_enq_bits_decodeResult_multiCycle;
  wire         queue_14_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_14 = {queue_14_enq_bits_decodeResult_multiCycle, queue_14_enq_bits_decodeResult_divider};
  wire         queue_14_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_14 = {queue_dataIn_lo_lo_lo_hi_hi_14, queue_14_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_14 = {queue_dataIn_lo_lo_lo_hi_14, queue_dataIn_lo_lo_lo_lo_14};
  wire         queue_14_enq_bits_decodeResult_unsigned1;
  wire         queue_14_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_14 = {queue_14_enq_bits_decodeResult_unsigned1, queue_14_enq_bits_decodeResult_unsigned0};
  wire         queue_14_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_14 = {queue_dataIn_lo_lo_hi_lo_hi_14, queue_14_enq_bits_decodeResult_other};
  wire         queue_14_enq_bits_decodeResult_red;
  wire         queue_14_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_14 = {queue_14_enq_bits_decodeResult_red, queue_14_enq_bits_decodeResult_nr};
  wire         queue_14_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_14 = {queue_dataIn_lo_lo_hi_hi_hi_14, queue_14_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_28 = {queue_dataIn_lo_lo_hi_hi_14, queue_dataIn_lo_lo_hi_lo_14};
  wire [11:0]  queue_dataIn_lo_lo_28 = {queue_dataIn_lo_lo_hi_28, queue_dataIn_lo_lo_lo_14};
  wire         queue_14_enq_bits_decodeResult_slid;
  wire         queue_14_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_14 = {queue_14_enq_bits_decodeResult_slid, queue_14_enq_bits_decodeResult_targetRd};
  wire         queue_14_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_14 = {queue_dataIn_lo_hi_lo_lo_hi_14, queue_14_enq_bits_decodeResult_widenReduce};
  wire         queue_14_enq_bits_decodeResult_compress;
  wire         queue_14_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_14 = {queue_14_enq_bits_decodeResult_compress, queue_14_enq_bits_decodeResult_gather16};
  wire         queue_14_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_14 = {queue_dataIn_lo_hi_lo_hi_hi_14, queue_14_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_28 = {queue_dataIn_lo_hi_lo_hi_14, queue_dataIn_lo_hi_lo_lo_14};
  wire         queue_14_enq_bits_decodeResult_mv;
  wire         queue_14_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_14 = {queue_14_enq_bits_decodeResult_mv, queue_14_enq_bits_decodeResult_extend};
  wire         queue_14_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_14 = {queue_dataIn_lo_hi_hi_lo_hi_14, queue_14_enq_bits_decodeResult_unOrderWrite};
  wire         queue_14_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_14_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_14 = {queue_14_enq_bits_decodeResult_maskLogic, queue_14_enq_bits_decodeResult_uop};
  wire         queue_14_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_14 = {queue_dataIn_lo_hi_hi_hi_hi_14, queue_14_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_28 = {queue_dataIn_lo_hi_hi_hi_14, queue_dataIn_lo_hi_hi_lo_14};
  wire [14:0]  queue_dataIn_lo_hi_43 = {queue_dataIn_lo_hi_hi_28, queue_dataIn_lo_hi_lo_28};
  wire [26:0]  queue_dataIn_lo_43 = {queue_dataIn_lo_hi_43, queue_dataIn_lo_lo_28};
  wire         queue_14_enq_bits_decodeResult_readOnly;
  wire         queue_14_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_14 = {queue_14_enq_bits_decodeResult_readOnly, queue_14_enq_bits_decodeResult_maskSource};
  wire         queue_14_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_14 = {queue_dataIn_hi_lo_lo_lo_hi_14, queue_14_enq_bits_decodeResult_maskDestination};
  wire         queue_14_enq_bits_decodeResult_special;
  wire         queue_14_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_14 = {queue_14_enq_bits_decodeResult_special, queue_14_enq_bits_decodeResult_saturate};
  wire         queue_14_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_14 = {queue_dataIn_hi_lo_lo_hi_hi_14, queue_14_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_28 = {queue_dataIn_hi_lo_lo_hi_14, queue_dataIn_hi_lo_lo_lo_14};
  wire         queue_14_enq_bits_decodeResult_crossRead;
  wire         queue_14_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_14 = {queue_14_enq_bits_decodeResult_crossRead, queue_14_enq_bits_decodeResult_crossWrite};
  wire         queue_14_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_14 = {queue_dataIn_hi_lo_hi_lo_hi_14, queue_14_enq_bits_decodeResult_maskUnit};
  wire         queue_14_enq_bits_decodeResult_sReadVD;
  wire         queue_14_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_14 = {queue_14_enq_bits_decodeResult_sReadVD, queue_14_enq_bits_decodeResult_vtype};
  wire         queue_14_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_14 = {queue_dataIn_hi_lo_hi_hi_hi_14, queue_14_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_28 = {queue_dataIn_hi_lo_hi_hi_14, queue_dataIn_hi_lo_hi_lo_14};
  wire [11:0]  queue_dataIn_hi_lo_43 = {queue_dataIn_hi_lo_hi_28, queue_dataIn_hi_lo_lo_28};
  wire         queue_14_enq_bits_decodeResult_reverse;
  wire         queue_14_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_14 = {queue_14_enq_bits_decodeResult_reverse, queue_14_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_14_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_14 = {queue_dataIn_hi_hi_lo_lo_hi_14, queue_14_enq_bits_decodeResult_scheduler};
  wire         queue_14_enq_bits_decodeResult_popCount;
  wire         queue_14_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_14 = {queue_14_enq_bits_decodeResult_popCount, queue_14_enq_bits_decodeResult_ffo};
  wire         queue_14_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_14 = {queue_dataIn_hi_hi_lo_hi_hi_14, queue_14_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_28 = {queue_dataIn_hi_hi_lo_hi_14, queue_dataIn_hi_hi_lo_lo_14};
  wire         queue_14_enq_bits_decodeResult_float;
  wire         queue_14_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_14 = {queue_14_enq_bits_decodeResult_float, queue_14_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_14_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_14 = {queue_dataIn_hi_hi_hi_lo_hi_14, queue_14_enq_bits_decodeResult_topUop};
  wire         queue_14_enq_bits_decodeResult_orderReduce;
  wire         queue_14_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_14 = {queue_14_enq_bits_decodeResult_orderReduce, queue_14_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_14_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_14 = {queue_dataIn_hi_hi_hi_hi_hi_14, queue_14_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_28 = {queue_dataIn_hi_hi_hi_hi_14, queue_dataIn_hi_hi_hi_lo_14};
  wire [16:0]  queue_dataIn_hi_hi_43 = {queue_dataIn_hi_hi_hi_28, queue_dataIn_hi_hi_lo_28};
  wire [28:0]  queue_dataIn_hi_43 = {queue_dataIn_hi_hi_43, queue_dataIn_hi_lo_43};
  wire [2:0]   queue_14_enq_bits_segment;
  wire [31:0]  queue_14_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_29 = {queue_14_enq_bits_segment, queue_14_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_29 = {queue_dataIn_lo_lo_hi_29, queue_dataIn_hi_42, queue_dataIn_lo_42};
  wire [1:0]   queue_14_enq_bits_loadStoreEEW;
  wire         queue_14_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_29 = {queue_14_enq_bits_loadStoreEEW, queue_14_enq_bits_mask};
  wire [4:0]   queue_14_enq_bits_vs2;
  wire [4:0]   queue_14_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_29 = {queue_14_enq_bits_vs2, queue_14_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_44 = {queue_dataIn_lo_hi_hi_29, queue_dataIn_lo_hi_lo_29};
  wire [80:0]  queue_dataIn_lo_44 = {queue_dataIn_lo_hi_44, queue_dataIn_lo_lo_29};
  wire         queue_14_enq_bits_lsWholeReg;
  wire [4:0]   queue_14_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_29 = {queue_14_enq_bits_lsWholeReg, queue_14_enq_bits_vs1};
  wire         queue_14_enq_bits_store;
  wire         queue_14_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_29 = {queue_14_enq_bits_store, queue_14_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_44 = {queue_dataIn_hi_lo_hi_29, queue_dataIn_hi_lo_lo_29};
  wire         queue_14_enq_bits_loadStore;
  wire         queue_14_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_29 = {queue_14_enq_bits_loadStore, queue_14_enq_bits_issueInst};
  wire [2:0]   queue_14_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_29 = {queue_14_enq_bits_instructionIndex, queue_dataIn_hi_43, queue_dataIn_lo_43};
  wire [60:0]  queue_dataIn_hi_hi_44 = {queue_dataIn_hi_hi_hi_29, queue_dataIn_hi_hi_lo_29};
  wire [68:0]  queue_dataIn_hi_44 = {queue_dataIn_hi_hi_44, queue_dataIn_hi_lo_44};
  wire [149:0] queue_dataIn_14 = {queue_dataIn_hi_44, queue_dataIn_lo_44};
  wire         queue_dataOut_14_csrInterface_vma = _queue_fifo_14_data_out[0];
  wire         queue_dataOut_14_csrInterface_vta = _queue_fifo_14_data_out[1];
  wire [1:0]   queue_dataOut_14_csrInterface_vxrm = _queue_fifo_14_data_out[3:2];
  wire [1:0]   queue_dataOut_14_csrInterface_vSew = _queue_fifo_14_data_out[5:4];
  wire [2:0]   queue_dataOut_14_csrInterface_vlmul = _queue_fifo_14_data_out[8:6];
  wire [11:0]  queue_dataOut_14_csrInterface_vStart = _queue_fifo_14_data_out[20:9];
  wire [11:0]  queue_dataOut_14_csrInterface_vl = _queue_fifo_14_data_out[32:21];
  wire [31:0]  queue_dataOut_14_readFromScalar = _queue_fifo_14_data_out[64:33];
  wire [2:0]   queue_dataOut_14_segment = _queue_fifo_14_data_out[67:65];
  wire         queue_dataOut_14_mask = _queue_fifo_14_data_out[68];
  wire [1:0]   queue_dataOut_14_loadStoreEEW = _queue_fifo_14_data_out[70:69];
  wire [4:0]   queue_dataOut_14_vd = _queue_fifo_14_data_out[75:71];
  wire [4:0]   queue_dataOut_14_vs2 = _queue_fifo_14_data_out[80:76];
  wire [4:0]   queue_dataOut_14_vs1 = _queue_fifo_14_data_out[85:81];
  wire         queue_dataOut_14_lsWholeReg = _queue_fifo_14_data_out[86];
  wire         queue_dataOut_14_special = _queue_fifo_14_data_out[87];
  wire         queue_dataOut_14_store = _queue_fifo_14_data_out[88];
  wire         queue_dataOut_14_issueInst = _queue_fifo_14_data_out[89];
  wire         queue_dataOut_14_loadStore = _queue_fifo_14_data_out[90];
  wire         queue_dataOut_14_decodeResult_logic = _queue_fifo_14_data_out[91];
  wire         queue_dataOut_14_decodeResult_adder = _queue_fifo_14_data_out[92];
  wire         queue_dataOut_14_decodeResult_shift = _queue_fifo_14_data_out[93];
  wire         queue_dataOut_14_decodeResult_multiplier = _queue_fifo_14_data_out[94];
  wire         queue_dataOut_14_decodeResult_divider = _queue_fifo_14_data_out[95];
  wire         queue_dataOut_14_decodeResult_multiCycle = _queue_fifo_14_data_out[96];
  wire         queue_dataOut_14_decodeResult_other = _queue_fifo_14_data_out[97];
  wire         queue_dataOut_14_decodeResult_unsigned0 = _queue_fifo_14_data_out[98];
  wire         queue_dataOut_14_decodeResult_unsigned1 = _queue_fifo_14_data_out[99];
  wire         queue_dataOut_14_decodeResult_itype = _queue_fifo_14_data_out[100];
  wire         queue_dataOut_14_decodeResult_nr = _queue_fifo_14_data_out[101];
  wire         queue_dataOut_14_decodeResult_red = _queue_fifo_14_data_out[102];
  wire         queue_dataOut_14_decodeResult_widenReduce = _queue_fifo_14_data_out[103];
  wire         queue_dataOut_14_decodeResult_targetRd = _queue_fifo_14_data_out[104];
  wire         queue_dataOut_14_decodeResult_slid = _queue_fifo_14_data_out[105];
  wire         queue_dataOut_14_decodeResult_gather = _queue_fifo_14_data_out[106];
  wire         queue_dataOut_14_decodeResult_gather16 = _queue_fifo_14_data_out[107];
  wire         queue_dataOut_14_decodeResult_compress = _queue_fifo_14_data_out[108];
  wire         queue_dataOut_14_decodeResult_unOrderWrite = _queue_fifo_14_data_out[109];
  wire         queue_dataOut_14_decodeResult_extend = _queue_fifo_14_data_out[110];
  wire         queue_dataOut_14_decodeResult_mv = _queue_fifo_14_data_out[111];
  wire         queue_dataOut_14_decodeResult_iota = _queue_fifo_14_data_out[112];
  wire [3:0]   queue_dataOut_14_decodeResult_uop = _queue_fifo_14_data_out[116:113];
  wire         queue_dataOut_14_decodeResult_maskLogic = _queue_fifo_14_data_out[117];
  wire         queue_dataOut_14_decodeResult_maskDestination = _queue_fifo_14_data_out[118];
  wire         queue_dataOut_14_decodeResult_maskSource = _queue_fifo_14_data_out[119];
  wire         queue_dataOut_14_decodeResult_readOnly = _queue_fifo_14_data_out[120];
  wire         queue_dataOut_14_decodeResult_vwmacc = _queue_fifo_14_data_out[121];
  wire         queue_dataOut_14_decodeResult_saturate = _queue_fifo_14_data_out[122];
  wire         queue_dataOut_14_decodeResult_special = _queue_fifo_14_data_out[123];
  wire         queue_dataOut_14_decodeResult_maskUnit = _queue_fifo_14_data_out[124];
  wire         queue_dataOut_14_decodeResult_crossWrite = _queue_fifo_14_data_out[125];
  wire         queue_dataOut_14_decodeResult_crossRead = _queue_fifo_14_data_out[126];
  wire         queue_dataOut_14_decodeResult_sWrite = _queue_fifo_14_data_out[127];
  wire         queue_dataOut_14_decodeResult_vtype = _queue_fifo_14_data_out[128];
  wire         queue_dataOut_14_decodeResult_sReadVD = _queue_fifo_14_data_out[129];
  wire         queue_dataOut_14_decodeResult_scheduler = _queue_fifo_14_data_out[130];
  wire         queue_dataOut_14_decodeResult_dontNeedExecuteInLane = _queue_fifo_14_data_out[131];
  wire         queue_dataOut_14_decodeResult_reverse = _queue_fifo_14_data_out[132];
  wire         queue_dataOut_14_decodeResult_average = _queue_fifo_14_data_out[133];
  wire         queue_dataOut_14_decodeResult_ffo = _queue_fifo_14_data_out[134];
  wire         queue_dataOut_14_decodeResult_popCount = _queue_fifo_14_data_out[135];
  wire [4:0]   queue_dataOut_14_decodeResult_topUop = _queue_fifo_14_data_out[140:136];
  wire         queue_dataOut_14_decodeResult_specialSlot = _queue_fifo_14_data_out[141];
  wire         queue_dataOut_14_decodeResult_float = _queue_fifo_14_data_out[142];
  wire [1:0]   queue_dataOut_14_decodeResult_fpExecutionType = _queue_fifo_14_data_out[144:143];
  wire         queue_dataOut_14_decodeResult_floatMul = _queue_fifo_14_data_out[145];
  wire         queue_dataOut_14_decodeResult_orderReduce = _queue_fifo_14_data_out[146];
  wire [2:0]   queue_dataOut_14_instructionIndex = _queue_fifo_14_data_out[149:147];
  wire         queue_14_enq_ready = ~_queue_fifo_14_full;
  wire         queue_14_enq_valid;
  assign queue_14_deq_valid = ~_queue_fifo_14_empty | queue_14_enq_valid;
  assign queue_14_deq_bits_instructionIndex = _queue_fifo_14_empty ? queue_14_enq_bits_instructionIndex : queue_dataOut_14_instructionIndex;
  assign queue_14_deq_bits_decodeResult_orderReduce = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_orderReduce : queue_dataOut_14_decodeResult_orderReduce;
  assign queue_14_deq_bits_decodeResult_floatMul = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_floatMul : queue_dataOut_14_decodeResult_floatMul;
  assign queue_14_deq_bits_decodeResult_fpExecutionType = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_fpExecutionType : queue_dataOut_14_decodeResult_fpExecutionType;
  assign queue_14_deq_bits_decodeResult_float = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_float : queue_dataOut_14_decodeResult_float;
  assign queue_14_deq_bits_decodeResult_specialSlot = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_specialSlot : queue_dataOut_14_decodeResult_specialSlot;
  assign queue_14_deq_bits_decodeResult_topUop = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_topUop : queue_dataOut_14_decodeResult_topUop;
  assign queue_14_deq_bits_decodeResult_popCount = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_popCount : queue_dataOut_14_decodeResult_popCount;
  assign queue_14_deq_bits_decodeResult_ffo = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_ffo : queue_dataOut_14_decodeResult_ffo;
  assign queue_14_deq_bits_decodeResult_average = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_average : queue_dataOut_14_decodeResult_average;
  assign queue_14_deq_bits_decodeResult_reverse = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_reverse : queue_dataOut_14_decodeResult_reverse;
  assign queue_14_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_14_decodeResult_dontNeedExecuteInLane;
  assign queue_14_deq_bits_decodeResult_scheduler = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_scheduler : queue_dataOut_14_decodeResult_scheduler;
  assign queue_14_deq_bits_decodeResult_sReadVD = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_sReadVD : queue_dataOut_14_decodeResult_sReadVD;
  assign queue_14_deq_bits_decodeResult_vtype = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_vtype : queue_dataOut_14_decodeResult_vtype;
  assign queue_14_deq_bits_decodeResult_sWrite = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_sWrite : queue_dataOut_14_decodeResult_sWrite;
  assign queue_14_deq_bits_decodeResult_crossRead = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_crossRead : queue_dataOut_14_decodeResult_crossRead;
  assign queue_14_deq_bits_decodeResult_crossWrite = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_crossWrite : queue_dataOut_14_decodeResult_crossWrite;
  assign queue_14_deq_bits_decodeResult_maskUnit = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_maskUnit : queue_dataOut_14_decodeResult_maskUnit;
  assign queue_14_deq_bits_decodeResult_special = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_special : queue_dataOut_14_decodeResult_special;
  assign queue_14_deq_bits_decodeResult_saturate = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_saturate : queue_dataOut_14_decodeResult_saturate;
  assign queue_14_deq_bits_decodeResult_vwmacc = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_vwmacc : queue_dataOut_14_decodeResult_vwmacc;
  assign queue_14_deq_bits_decodeResult_readOnly = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_readOnly : queue_dataOut_14_decodeResult_readOnly;
  assign queue_14_deq_bits_decodeResult_maskSource = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_maskSource : queue_dataOut_14_decodeResult_maskSource;
  assign queue_14_deq_bits_decodeResult_maskDestination = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_maskDestination : queue_dataOut_14_decodeResult_maskDestination;
  assign queue_14_deq_bits_decodeResult_maskLogic = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_maskLogic : queue_dataOut_14_decodeResult_maskLogic;
  assign queue_14_deq_bits_decodeResult_uop = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_uop : queue_dataOut_14_decodeResult_uop;
  assign queue_14_deq_bits_decodeResult_iota = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_iota : queue_dataOut_14_decodeResult_iota;
  assign queue_14_deq_bits_decodeResult_mv = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_mv : queue_dataOut_14_decodeResult_mv;
  assign queue_14_deq_bits_decodeResult_extend = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_extend : queue_dataOut_14_decodeResult_extend;
  assign queue_14_deq_bits_decodeResult_unOrderWrite = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_unOrderWrite : queue_dataOut_14_decodeResult_unOrderWrite;
  assign queue_14_deq_bits_decodeResult_compress = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_compress : queue_dataOut_14_decodeResult_compress;
  assign queue_14_deq_bits_decodeResult_gather16 = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_gather16 : queue_dataOut_14_decodeResult_gather16;
  assign queue_14_deq_bits_decodeResult_gather = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_gather : queue_dataOut_14_decodeResult_gather;
  assign queue_14_deq_bits_decodeResult_slid = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_slid : queue_dataOut_14_decodeResult_slid;
  assign queue_14_deq_bits_decodeResult_targetRd = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_targetRd : queue_dataOut_14_decodeResult_targetRd;
  assign queue_14_deq_bits_decodeResult_widenReduce = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_widenReduce : queue_dataOut_14_decodeResult_widenReduce;
  assign queue_14_deq_bits_decodeResult_red = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_red : queue_dataOut_14_decodeResult_red;
  assign queue_14_deq_bits_decodeResult_nr = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_nr : queue_dataOut_14_decodeResult_nr;
  assign queue_14_deq_bits_decodeResult_itype = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_itype : queue_dataOut_14_decodeResult_itype;
  assign queue_14_deq_bits_decodeResult_unsigned1 = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_unsigned1 : queue_dataOut_14_decodeResult_unsigned1;
  assign queue_14_deq_bits_decodeResult_unsigned0 = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_unsigned0 : queue_dataOut_14_decodeResult_unsigned0;
  assign queue_14_deq_bits_decodeResult_other = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_other : queue_dataOut_14_decodeResult_other;
  assign queue_14_deq_bits_decodeResult_multiCycle = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_multiCycle : queue_dataOut_14_decodeResult_multiCycle;
  assign queue_14_deq_bits_decodeResult_divider = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_divider : queue_dataOut_14_decodeResult_divider;
  assign queue_14_deq_bits_decodeResult_multiplier = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_multiplier : queue_dataOut_14_decodeResult_multiplier;
  assign queue_14_deq_bits_decodeResult_shift = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_shift : queue_dataOut_14_decodeResult_shift;
  assign queue_14_deq_bits_decodeResult_adder = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_adder : queue_dataOut_14_decodeResult_adder;
  assign queue_14_deq_bits_decodeResult_logic = _queue_fifo_14_empty ? queue_14_enq_bits_decodeResult_logic : queue_dataOut_14_decodeResult_logic;
  assign queue_14_deq_bits_loadStore = _queue_fifo_14_empty ? queue_14_enq_bits_loadStore : queue_dataOut_14_loadStore;
  assign queue_14_deq_bits_issueInst = _queue_fifo_14_empty ? queue_14_enq_bits_issueInst : queue_dataOut_14_issueInst;
  assign queue_14_deq_bits_store = _queue_fifo_14_empty ? queue_14_enq_bits_store : queue_dataOut_14_store;
  assign queue_14_deq_bits_special = _queue_fifo_14_empty ? queue_14_enq_bits_special : queue_dataOut_14_special;
  assign queue_14_deq_bits_lsWholeReg = _queue_fifo_14_empty ? queue_14_enq_bits_lsWholeReg : queue_dataOut_14_lsWholeReg;
  assign queue_14_deq_bits_vs1 = _queue_fifo_14_empty ? queue_14_enq_bits_vs1 : queue_dataOut_14_vs1;
  assign queue_14_deq_bits_vs2 = _queue_fifo_14_empty ? queue_14_enq_bits_vs2 : queue_dataOut_14_vs2;
  assign queue_14_deq_bits_vd = _queue_fifo_14_empty ? queue_14_enq_bits_vd : queue_dataOut_14_vd;
  assign queue_14_deq_bits_loadStoreEEW = _queue_fifo_14_empty ? queue_14_enq_bits_loadStoreEEW : queue_dataOut_14_loadStoreEEW;
  assign queue_14_deq_bits_mask = _queue_fifo_14_empty ? queue_14_enq_bits_mask : queue_dataOut_14_mask;
  assign queue_14_deq_bits_segment = _queue_fifo_14_empty ? queue_14_enq_bits_segment : queue_dataOut_14_segment;
  assign queue_14_deq_bits_readFromScalar = _queue_fifo_14_empty ? queue_14_enq_bits_readFromScalar : queue_dataOut_14_readFromScalar;
  assign queue_14_deq_bits_csrInterface_vl = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vl : queue_dataOut_14_csrInterface_vl;
  assign queue_14_deq_bits_csrInterface_vStart = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vStart : queue_dataOut_14_csrInterface_vStart;
  assign queue_14_deq_bits_csrInterface_vlmul = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vlmul : queue_dataOut_14_csrInterface_vlmul;
  assign queue_14_deq_bits_csrInterface_vSew = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vSew : queue_dataOut_14_csrInterface_vSew;
  assign queue_14_deq_bits_csrInterface_vxrm = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vxrm : queue_dataOut_14_csrInterface_vxrm;
  assign queue_14_deq_bits_csrInterface_vta = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vta : queue_dataOut_14_csrInterface_vta;
  assign queue_14_deq_bits_csrInterface_vma = _queue_fifo_14_empty ? queue_14_enq_bits_csrInterface_vma : queue_dataOut_14_csrInterface_vma;
  wire         laneVec_14_laneRequest_bits_issueInst = laneRequestSinkWire_14_ready & laneRequestSinkWire_14_valid;
  reg          releasePipe_pipe_v_14;
  wire         releasePipe_pipe_out_14_valid = releasePipe_pipe_v_14;
  wire         laneRequestSourceWire_14_ready;
  wire         validSource_14_valid = laneRequestSourceWire_14_ready & laneRequestSourceWire_14_valid;
  reg  [2:0]   tokenCheck_counter_14;
  wire [2:0]   tokenCheck_counterChange_14 = validSource_14_valid ? 3'h1 : 3'h7;
  assign tokenCheck_14 = ~(tokenCheck_counter_14[2]);
  assign laneRequestSourceWire_14_ready = tokenCheck_14;
  assign queue_14_enq_valid = validSink_14_valid;
  assign queue_14_enq_bits_instructionIndex = validSink_14_bits_instructionIndex;
  assign queue_14_enq_bits_decodeResult_orderReduce = validSink_14_bits_decodeResult_orderReduce;
  assign queue_14_enq_bits_decodeResult_floatMul = validSink_14_bits_decodeResult_floatMul;
  assign queue_14_enq_bits_decodeResult_fpExecutionType = validSink_14_bits_decodeResult_fpExecutionType;
  assign queue_14_enq_bits_decodeResult_float = validSink_14_bits_decodeResult_float;
  assign queue_14_enq_bits_decodeResult_specialSlot = validSink_14_bits_decodeResult_specialSlot;
  assign queue_14_enq_bits_decodeResult_topUop = validSink_14_bits_decodeResult_topUop;
  assign queue_14_enq_bits_decodeResult_popCount = validSink_14_bits_decodeResult_popCount;
  assign queue_14_enq_bits_decodeResult_ffo = validSink_14_bits_decodeResult_ffo;
  assign queue_14_enq_bits_decodeResult_average = validSink_14_bits_decodeResult_average;
  assign queue_14_enq_bits_decodeResult_reverse = validSink_14_bits_decodeResult_reverse;
  assign queue_14_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_14_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_14_enq_bits_decodeResult_scheduler = validSink_14_bits_decodeResult_scheduler;
  assign queue_14_enq_bits_decodeResult_sReadVD = validSink_14_bits_decodeResult_sReadVD;
  assign queue_14_enq_bits_decodeResult_vtype = validSink_14_bits_decodeResult_vtype;
  assign queue_14_enq_bits_decodeResult_sWrite = validSink_14_bits_decodeResult_sWrite;
  assign queue_14_enq_bits_decodeResult_crossRead = validSink_14_bits_decodeResult_crossRead;
  assign queue_14_enq_bits_decodeResult_crossWrite = validSink_14_bits_decodeResult_crossWrite;
  assign queue_14_enq_bits_decodeResult_maskUnit = validSink_14_bits_decodeResult_maskUnit;
  assign queue_14_enq_bits_decodeResult_special = validSink_14_bits_decodeResult_special;
  assign queue_14_enq_bits_decodeResult_saturate = validSink_14_bits_decodeResult_saturate;
  assign queue_14_enq_bits_decodeResult_vwmacc = validSink_14_bits_decodeResult_vwmacc;
  assign queue_14_enq_bits_decodeResult_readOnly = validSink_14_bits_decodeResult_readOnly;
  assign queue_14_enq_bits_decodeResult_maskSource = validSink_14_bits_decodeResult_maskSource;
  assign queue_14_enq_bits_decodeResult_maskDestination = validSink_14_bits_decodeResult_maskDestination;
  assign queue_14_enq_bits_decodeResult_maskLogic = validSink_14_bits_decodeResult_maskLogic;
  assign queue_14_enq_bits_decodeResult_uop = validSink_14_bits_decodeResult_uop;
  assign queue_14_enq_bits_decodeResult_iota = validSink_14_bits_decodeResult_iota;
  assign queue_14_enq_bits_decodeResult_mv = validSink_14_bits_decodeResult_mv;
  assign queue_14_enq_bits_decodeResult_extend = validSink_14_bits_decodeResult_extend;
  assign queue_14_enq_bits_decodeResult_unOrderWrite = validSink_14_bits_decodeResult_unOrderWrite;
  assign queue_14_enq_bits_decodeResult_compress = validSink_14_bits_decodeResult_compress;
  assign queue_14_enq_bits_decodeResult_gather16 = validSink_14_bits_decodeResult_gather16;
  assign queue_14_enq_bits_decodeResult_gather = validSink_14_bits_decodeResult_gather;
  assign queue_14_enq_bits_decodeResult_slid = validSink_14_bits_decodeResult_slid;
  assign queue_14_enq_bits_decodeResult_targetRd = validSink_14_bits_decodeResult_targetRd;
  assign queue_14_enq_bits_decodeResult_widenReduce = validSink_14_bits_decodeResult_widenReduce;
  assign queue_14_enq_bits_decodeResult_red = validSink_14_bits_decodeResult_red;
  assign queue_14_enq_bits_decodeResult_nr = validSink_14_bits_decodeResult_nr;
  assign queue_14_enq_bits_decodeResult_itype = validSink_14_bits_decodeResult_itype;
  assign queue_14_enq_bits_decodeResult_unsigned1 = validSink_14_bits_decodeResult_unsigned1;
  assign queue_14_enq_bits_decodeResult_unsigned0 = validSink_14_bits_decodeResult_unsigned0;
  assign queue_14_enq_bits_decodeResult_other = validSink_14_bits_decodeResult_other;
  assign queue_14_enq_bits_decodeResult_multiCycle = validSink_14_bits_decodeResult_multiCycle;
  assign queue_14_enq_bits_decodeResult_divider = validSink_14_bits_decodeResult_divider;
  assign queue_14_enq_bits_decodeResult_multiplier = validSink_14_bits_decodeResult_multiplier;
  assign queue_14_enq_bits_decodeResult_shift = validSink_14_bits_decodeResult_shift;
  assign queue_14_enq_bits_decodeResult_adder = validSink_14_bits_decodeResult_adder;
  assign queue_14_enq_bits_decodeResult_logic = validSink_14_bits_decodeResult_logic;
  assign queue_14_enq_bits_loadStore = validSink_14_bits_loadStore;
  assign queue_14_enq_bits_issueInst = validSink_14_bits_issueInst;
  assign queue_14_enq_bits_store = validSink_14_bits_store;
  assign queue_14_enq_bits_special = validSink_14_bits_special;
  assign queue_14_enq_bits_lsWholeReg = validSink_14_bits_lsWholeReg;
  assign queue_14_enq_bits_vs1 = validSink_14_bits_vs1;
  assign queue_14_enq_bits_vs2 = validSink_14_bits_vs2;
  assign queue_14_enq_bits_vd = validSink_14_bits_vd;
  assign queue_14_enq_bits_loadStoreEEW = validSink_14_bits_loadStoreEEW;
  assign queue_14_enq_bits_mask = validSink_14_bits_mask;
  assign queue_14_enq_bits_segment = validSink_14_bits_segment;
  assign queue_14_enq_bits_readFromScalar = validSink_14_bits_readFromScalar;
  assign queue_14_enq_bits_csrInterface_vl = validSink_14_bits_csrInterface_vl;
  assign queue_14_enq_bits_csrInterface_vStart = validSink_14_bits_csrInterface_vStart;
  assign queue_14_enq_bits_csrInterface_vlmul = validSink_14_bits_csrInterface_vlmul;
  assign queue_14_enq_bits_csrInterface_vSew = validSink_14_bits_csrInterface_vSew;
  assign queue_14_enq_bits_csrInterface_vxrm = validSink_14_bits_csrInterface_vxrm;
  assign queue_14_enq_bits_csrInterface_vta = validSink_14_bits_csrInterface_vta;
  assign queue_14_enq_bits_csrInterface_vma = validSink_14_bits_csrInterface_vma;
  reg          shifterReg_14_0_valid;
  assign validSink_14_valid = shifterReg_14_0_valid;
  reg  [2:0]   shifterReg_14_0_bits_instructionIndex;
  assign validSink_14_bits_instructionIndex = shifterReg_14_0_bits_instructionIndex;
  reg          shifterReg_14_0_bits_decodeResult_orderReduce;
  assign validSink_14_bits_decodeResult_orderReduce = shifterReg_14_0_bits_decodeResult_orderReduce;
  reg          shifterReg_14_0_bits_decodeResult_floatMul;
  assign validSink_14_bits_decodeResult_floatMul = shifterReg_14_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_14_0_bits_decodeResult_fpExecutionType;
  assign validSink_14_bits_decodeResult_fpExecutionType = shifterReg_14_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_14_0_bits_decodeResult_float;
  assign validSink_14_bits_decodeResult_float = shifterReg_14_0_bits_decodeResult_float;
  reg          shifterReg_14_0_bits_decodeResult_specialSlot;
  assign validSink_14_bits_decodeResult_specialSlot = shifterReg_14_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_14_0_bits_decodeResult_topUop;
  assign validSink_14_bits_decodeResult_topUop = shifterReg_14_0_bits_decodeResult_topUop;
  reg          shifterReg_14_0_bits_decodeResult_popCount;
  assign validSink_14_bits_decodeResult_popCount = shifterReg_14_0_bits_decodeResult_popCount;
  reg          shifterReg_14_0_bits_decodeResult_ffo;
  assign validSink_14_bits_decodeResult_ffo = shifterReg_14_0_bits_decodeResult_ffo;
  reg          shifterReg_14_0_bits_decodeResult_average;
  assign validSink_14_bits_decodeResult_average = shifterReg_14_0_bits_decodeResult_average;
  reg          shifterReg_14_0_bits_decodeResult_reverse;
  assign validSink_14_bits_decodeResult_reverse = shifterReg_14_0_bits_decodeResult_reverse;
  reg          shifterReg_14_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_14_bits_decodeResult_dontNeedExecuteInLane = shifterReg_14_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_14_0_bits_decodeResult_scheduler;
  assign validSink_14_bits_decodeResult_scheduler = shifterReg_14_0_bits_decodeResult_scheduler;
  reg          shifterReg_14_0_bits_decodeResult_sReadVD;
  assign validSink_14_bits_decodeResult_sReadVD = shifterReg_14_0_bits_decodeResult_sReadVD;
  reg          shifterReg_14_0_bits_decodeResult_vtype;
  assign validSink_14_bits_decodeResult_vtype = shifterReg_14_0_bits_decodeResult_vtype;
  reg          shifterReg_14_0_bits_decodeResult_sWrite;
  assign validSink_14_bits_decodeResult_sWrite = shifterReg_14_0_bits_decodeResult_sWrite;
  reg          shifterReg_14_0_bits_decodeResult_crossRead;
  assign validSink_14_bits_decodeResult_crossRead = shifterReg_14_0_bits_decodeResult_crossRead;
  reg          shifterReg_14_0_bits_decodeResult_crossWrite;
  assign validSink_14_bits_decodeResult_crossWrite = shifterReg_14_0_bits_decodeResult_crossWrite;
  reg          shifterReg_14_0_bits_decodeResult_maskUnit;
  assign validSink_14_bits_decodeResult_maskUnit = shifterReg_14_0_bits_decodeResult_maskUnit;
  reg          shifterReg_14_0_bits_decodeResult_special;
  assign validSink_14_bits_decodeResult_special = shifterReg_14_0_bits_decodeResult_special;
  reg          shifterReg_14_0_bits_decodeResult_saturate;
  assign validSink_14_bits_decodeResult_saturate = shifterReg_14_0_bits_decodeResult_saturate;
  reg          shifterReg_14_0_bits_decodeResult_vwmacc;
  assign validSink_14_bits_decodeResult_vwmacc = shifterReg_14_0_bits_decodeResult_vwmacc;
  reg          shifterReg_14_0_bits_decodeResult_readOnly;
  assign validSink_14_bits_decodeResult_readOnly = shifterReg_14_0_bits_decodeResult_readOnly;
  reg          shifterReg_14_0_bits_decodeResult_maskSource;
  assign validSink_14_bits_decodeResult_maskSource = shifterReg_14_0_bits_decodeResult_maskSource;
  reg          shifterReg_14_0_bits_decodeResult_maskDestination;
  assign validSink_14_bits_decodeResult_maskDestination = shifterReg_14_0_bits_decodeResult_maskDestination;
  reg          shifterReg_14_0_bits_decodeResult_maskLogic;
  assign validSink_14_bits_decodeResult_maskLogic = shifterReg_14_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_14_0_bits_decodeResult_uop;
  assign validSink_14_bits_decodeResult_uop = shifterReg_14_0_bits_decodeResult_uop;
  reg          shifterReg_14_0_bits_decodeResult_iota;
  assign validSink_14_bits_decodeResult_iota = shifterReg_14_0_bits_decodeResult_iota;
  reg          shifterReg_14_0_bits_decodeResult_mv;
  assign validSink_14_bits_decodeResult_mv = shifterReg_14_0_bits_decodeResult_mv;
  reg          shifterReg_14_0_bits_decodeResult_extend;
  assign validSink_14_bits_decodeResult_extend = shifterReg_14_0_bits_decodeResult_extend;
  reg          shifterReg_14_0_bits_decodeResult_unOrderWrite;
  assign validSink_14_bits_decodeResult_unOrderWrite = shifterReg_14_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_14_0_bits_decodeResult_compress;
  assign validSink_14_bits_decodeResult_compress = shifterReg_14_0_bits_decodeResult_compress;
  reg          shifterReg_14_0_bits_decodeResult_gather16;
  assign validSink_14_bits_decodeResult_gather16 = shifterReg_14_0_bits_decodeResult_gather16;
  reg          shifterReg_14_0_bits_decodeResult_gather;
  assign validSink_14_bits_decodeResult_gather = shifterReg_14_0_bits_decodeResult_gather;
  reg          shifterReg_14_0_bits_decodeResult_slid;
  assign validSink_14_bits_decodeResult_slid = shifterReg_14_0_bits_decodeResult_slid;
  reg          shifterReg_14_0_bits_decodeResult_targetRd;
  assign validSink_14_bits_decodeResult_targetRd = shifterReg_14_0_bits_decodeResult_targetRd;
  reg          shifterReg_14_0_bits_decodeResult_widenReduce;
  assign validSink_14_bits_decodeResult_widenReduce = shifterReg_14_0_bits_decodeResult_widenReduce;
  reg          shifterReg_14_0_bits_decodeResult_red;
  assign validSink_14_bits_decodeResult_red = shifterReg_14_0_bits_decodeResult_red;
  reg          shifterReg_14_0_bits_decodeResult_nr;
  assign validSink_14_bits_decodeResult_nr = shifterReg_14_0_bits_decodeResult_nr;
  reg          shifterReg_14_0_bits_decodeResult_itype;
  assign validSink_14_bits_decodeResult_itype = shifterReg_14_0_bits_decodeResult_itype;
  reg          shifterReg_14_0_bits_decodeResult_unsigned1;
  assign validSink_14_bits_decodeResult_unsigned1 = shifterReg_14_0_bits_decodeResult_unsigned1;
  reg          shifterReg_14_0_bits_decodeResult_unsigned0;
  assign validSink_14_bits_decodeResult_unsigned0 = shifterReg_14_0_bits_decodeResult_unsigned0;
  reg          shifterReg_14_0_bits_decodeResult_other;
  assign validSink_14_bits_decodeResult_other = shifterReg_14_0_bits_decodeResult_other;
  reg          shifterReg_14_0_bits_decodeResult_multiCycle;
  assign validSink_14_bits_decodeResult_multiCycle = shifterReg_14_0_bits_decodeResult_multiCycle;
  reg          shifterReg_14_0_bits_decodeResult_divider;
  assign validSink_14_bits_decodeResult_divider = shifterReg_14_0_bits_decodeResult_divider;
  reg          shifterReg_14_0_bits_decodeResult_multiplier;
  assign validSink_14_bits_decodeResult_multiplier = shifterReg_14_0_bits_decodeResult_multiplier;
  reg          shifterReg_14_0_bits_decodeResult_shift;
  assign validSink_14_bits_decodeResult_shift = shifterReg_14_0_bits_decodeResult_shift;
  reg          shifterReg_14_0_bits_decodeResult_adder;
  assign validSink_14_bits_decodeResult_adder = shifterReg_14_0_bits_decodeResult_adder;
  reg          shifterReg_14_0_bits_decodeResult_logic;
  assign validSink_14_bits_decodeResult_logic = shifterReg_14_0_bits_decodeResult_logic;
  reg          shifterReg_14_0_bits_loadStore;
  assign validSink_14_bits_loadStore = shifterReg_14_0_bits_loadStore;
  reg          shifterReg_14_0_bits_issueInst;
  assign validSink_14_bits_issueInst = shifterReg_14_0_bits_issueInst;
  reg          shifterReg_14_0_bits_store;
  assign validSink_14_bits_store = shifterReg_14_0_bits_store;
  reg          shifterReg_14_0_bits_special;
  assign validSink_14_bits_special = shifterReg_14_0_bits_special;
  reg          shifterReg_14_0_bits_lsWholeReg;
  assign validSink_14_bits_lsWholeReg = shifterReg_14_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_14_0_bits_vs1;
  assign validSink_14_bits_vs1 = shifterReg_14_0_bits_vs1;
  reg  [4:0]   shifterReg_14_0_bits_vs2;
  assign validSink_14_bits_vs2 = shifterReg_14_0_bits_vs2;
  reg  [4:0]   shifterReg_14_0_bits_vd;
  assign validSink_14_bits_vd = shifterReg_14_0_bits_vd;
  reg  [1:0]   shifterReg_14_0_bits_loadStoreEEW;
  assign validSink_14_bits_loadStoreEEW = shifterReg_14_0_bits_loadStoreEEW;
  reg          shifterReg_14_0_bits_mask;
  assign validSink_14_bits_mask = shifterReg_14_0_bits_mask;
  reg  [2:0]   shifterReg_14_0_bits_segment;
  assign validSink_14_bits_segment = shifterReg_14_0_bits_segment;
  reg  [31:0]  shifterReg_14_0_bits_readFromScalar;
  assign validSink_14_bits_readFromScalar = shifterReg_14_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_14_0_bits_csrInterface_vl;
  assign validSink_14_bits_csrInterface_vl = shifterReg_14_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_14_0_bits_csrInterface_vStart;
  assign validSink_14_bits_csrInterface_vStart = shifterReg_14_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_14_0_bits_csrInterface_vlmul;
  assign validSink_14_bits_csrInterface_vlmul = shifterReg_14_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_14_0_bits_csrInterface_vSew;
  assign validSink_14_bits_csrInterface_vSew = shifterReg_14_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_14_0_bits_csrInterface_vxrm;
  assign validSink_14_bits_csrInterface_vxrm = shifterReg_14_0_bits_csrInterface_vxrm;
  reg          shifterReg_14_0_bits_csrInterface_vta;
  assign validSink_14_bits_csrInterface_vta = shifterReg_14_0_bits_csrInterface_vta;
  reg          shifterReg_14_0_bits_csrInterface_vma;
  assign validSink_14_bits_csrInterface_vma = shifterReg_14_0_bits_csrInterface_vma;
  wire         shifterValid_14 = shifterReg_14_0_valid | validSource_14_valid;
  wire         validSink_15_valid;
  wire [2:0]   validSink_15_bits_instructionIndex;
  wire         validSink_15_bits_decodeResult_orderReduce;
  wire         validSink_15_bits_decodeResult_floatMul;
  wire [1:0]   validSink_15_bits_decodeResult_fpExecutionType;
  wire         validSink_15_bits_decodeResult_float;
  wire         validSink_15_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_15_bits_decodeResult_topUop;
  wire         validSink_15_bits_decodeResult_popCount;
  wire         validSink_15_bits_decodeResult_ffo;
  wire         validSink_15_bits_decodeResult_average;
  wire         validSink_15_bits_decodeResult_reverse;
  wire         validSink_15_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_15_bits_decodeResult_scheduler;
  wire         validSink_15_bits_decodeResult_sReadVD;
  wire         validSink_15_bits_decodeResult_vtype;
  wire         validSink_15_bits_decodeResult_sWrite;
  wire         validSink_15_bits_decodeResult_crossRead;
  wire         validSink_15_bits_decodeResult_crossWrite;
  wire         validSink_15_bits_decodeResult_maskUnit;
  wire         validSink_15_bits_decodeResult_special;
  wire         validSink_15_bits_decodeResult_saturate;
  wire         validSink_15_bits_decodeResult_vwmacc;
  wire         validSink_15_bits_decodeResult_readOnly;
  wire         validSink_15_bits_decodeResult_maskSource;
  wire         validSink_15_bits_decodeResult_maskDestination;
  wire         validSink_15_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_15_bits_decodeResult_uop;
  wire         validSink_15_bits_decodeResult_iota;
  wire         validSink_15_bits_decodeResult_mv;
  wire         validSink_15_bits_decodeResult_extend;
  wire         validSink_15_bits_decodeResult_unOrderWrite;
  wire         validSink_15_bits_decodeResult_compress;
  wire         validSink_15_bits_decodeResult_gather16;
  wire         validSink_15_bits_decodeResult_gather;
  wire         validSink_15_bits_decodeResult_slid;
  wire         validSink_15_bits_decodeResult_targetRd;
  wire         validSink_15_bits_decodeResult_widenReduce;
  wire         validSink_15_bits_decodeResult_red;
  wire         validSink_15_bits_decodeResult_nr;
  wire         validSink_15_bits_decodeResult_itype;
  wire         validSink_15_bits_decodeResult_unsigned1;
  wire         validSink_15_bits_decodeResult_unsigned0;
  wire         validSink_15_bits_decodeResult_other;
  wire         validSink_15_bits_decodeResult_multiCycle;
  wire         validSink_15_bits_decodeResult_divider;
  wire         validSink_15_bits_decodeResult_multiplier;
  wire         validSink_15_bits_decodeResult_shift;
  wire         validSink_15_bits_decodeResult_adder;
  wire         validSink_15_bits_decodeResult_logic;
  wire         validSink_15_bits_loadStore;
  wire         validSink_15_bits_issueInst;
  wire         validSink_15_bits_store;
  wire         validSink_15_bits_special;
  wire         validSink_15_bits_lsWholeReg;
  wire [4:0]   validSink_15_bits_vs1;
  wire [4:0]   validSink_15_bits_vs2;
  wire [4:0]   validSink_15_bits_vd;
  wire [1:0]   validSink_15_bits_loadStoreEEW;
  wire         validSink_15_bits_mask;
  wire [2:0]   validSink_15_bits_segment;
  wire [31:0]  validSink_15_bits_readFromScalar;
  wire [11:0]  validSink_15_bits_csrInterface_vl;
  wire [11:0]  validSink_15_bits_csrInterface_vStart;
  wire [2:0]   validSink_15_bits_csrInterface_vlmul;
  wire [1:0]   validSink_15_bits_csrInterface_vSew;
  wire [1:0]   validSink_15_bits_csrInterface_vxrm;
  wire         validSink_15_bits_csrInterface_vta;
  wire         validSink_15_bits_csrInterface_vma;
  wire         laneRequestSinkWire_15_valid = queue_15_deq_valid;
  wire [2:0]   laneRequestSinkWire_15_bits_instructionIndex = queue_15_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_15_bits_decodeResult_orderReduce = queue_15_deq_bits_decodeResult_orderReduce;
  wire         laneRequestSinkWire_15_bits_decodeResult_floatMul = queue_15_deq_bits_decodeResult_floatMul;
  wire [1:0]   laneRequestSinkWire_15_bits_decodeResult_fpExecutionType = queue_15_deq_bits_decodeResult_fpExecutionType;
  wire         laneRequestSinkWire_15_bits_decodeResult_float = queue_15_deq_bits_decodeResult_float;
  wire         laneRequestSinkWire_15_bits_decodeResult_specialSlot = queue_15_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_15_bits_decodeResult_topUop = queue_15_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_15_bits_decodeResult_popCount = queue_15_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_15_bits_decodeResult_ffo = queue_15_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_15_bits_decodeResult_average = queue_15_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_15_bits_decodeResult_reverse = queue_15_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_15_bits_decodeResult_dontNeedExecuteInLane = queue_15_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_15_bits_decodeResult_scheduler = queue_15_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_15_bits_decodeResult_sReadVD = queue_15_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_15_bits_decodeResult_vtype = queue_15_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_15_bits_decodeResult_sWrite = queue_15_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_15_bits_decodeResult_crossRead = queue_15_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_15_bits_decodeResult_crossWrite = queue_15_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_15_bits_decodeResult_maskUnit = queue_15_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_15_bits_decodeResult_special = queue_15_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_15_bits_decodeResult_saturate = queue_15_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_15_bits_decodeResult_vwmacc = queue_15_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_15_bits_decodeResult_readOnly = queue_15_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_15_bits_decodeResult_maskSource = queue_15_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_15_bits_decodeResult_maskDestination = queue_15_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_15_bits_decodeResult_maskLogic = queue_15_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_15_bits_decodeResult_uop = queue_15_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_15_bits_decodeResult_iota = queue_15_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_15_bits_decodeResult_mv = queue_15_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_15_bits_decodeResult_extend = queue_15_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_15_bits_decodeResult_unOrderWrite = queue_15_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_15_bits_decodeResult_compress = queue_15_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_15_bits_decodeResult_gather16 = queue_15_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_15_bits_decodeResult_gather = queue_15_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_15_bits_decodeResult_slid = queue_15_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_15_bits_decodeResult_targetRd = queue_15_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_15_bits_decodeResult_widenReduce = queue_15_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_15_bits_decodeResult_red = queue_15_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_15_bits_decodeResult_nr = queue_15_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_15_bits_decodeResult_itype = queue_15_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_15_bits_decodeResult_unsigned1 = queue_15_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_15_bits_decodeResult_unsigned0 = queue_15_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_15_bits_decodeResult_other = queue_15_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_15_bits_decodeResult_multiCycle = queue_15_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_15_bits_decodeResult_divider = queue_15_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_15_bits_decodeResult_multiplier = queue_15_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_15_bits_decodeResult_shift = queue_15_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_15_bits_decodeResult_adder = queue_15_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_15_bits_decodeResult_logic = queue_15_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_15_bits_loadStore = queue_15_deq_bits_loadStore;
  wire         laneRequestSinkWire_15_bits_issueInst = queue_15_deq_bits_issueInst;
  wire         laneRequestSinkWire_15_bits_store = queue_15_deq_bits_store;
  wire         laneRequestSinkWire_15_bits_special = queue_15_deq_bits_special;
  wire         laneRequestSinkWire_15_bits_lsWholeReg = queue_15_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_15_bits_vs1 = queue_15_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_15_bits_vs2 = queue_15_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_15_bits_vd = queue_15_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_15_bits_loadStoreEEW = queue_15_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_15_bits_mask = queue_15_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_15_bits_segment = queue_15_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_15_bits_readFromScalar = queue_15_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_15_bits_csrInterface_vl = queue_15_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_15_bits_csrInterface_vStart = queue_15_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_15_bits_csrInterface_vlmul = queue_15_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_15_bits_csrInterface_vSew = queue_15_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_15_bits_csrInterface_vxrm = queue_15_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_15_bits_csrInterface_vta = queue_15_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_15_bits_csrInterface_vma = queue_15_deq_bits_csrInterface_vma;
  wire [1:0]   queue_15_enq_bits_csrInterface_vxrm;
  wire         queue_15_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_45 = {queue_15_enq_bits_csrInterface_vxrm, queue_15_enq_bits_csrInterface_vta};
  wire         queue_15_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_45 = {queue_dataIn_lo_hi_45, queue_15_enq_bits_csrInterface_vma};
  wire [2:0]   queue_15_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_15_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_45 = {queue_15_enq_bits_csrInterface_vlmul, queue_15_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_15_enq_bits_csrInterface_vl;
  wire [11:0]  queue_15_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_45 = {queue_15_enq_bits_csrInterface_vl, queue_15_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_45 = {queue_dataIn_hi_hi_45, queue_dataIn_hi_lo_45};
  wire         queue_15_enq_bits_decodeResult_shift;
  wire         queue_15_enq_bits_decodeResult_adder;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_hi_15 = {queue_15_enq_bits_decodeResult_shift, queue_15_enq_bits_decodeResult_adder};
  wire         queue_15_enq_bits_decodeResult_logic;
  wire [2:0]   queue_dataIn_lo_lo_lo_lo_15 = {queue_dataIn_lo_lo_lo_lo_hi_15, queue_15_enq_bits_decodeResult_logic};
  wire         queue_15_enq_bits_decodeResult_multiCycle;
  wire         queue_15_enq_bits_decodeResult_divider;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_15 = {queue_15_enq_bits_decodeResult_multiCycle, queue_15_enq_bits_decodeResult_divider};
  wire         queue_15_enq_bits_decodeResult_multiplier;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_15 = {queue_dataIn_lo_lo_lo_hi_hi_15, queue_15_enq_bits_decodeResult_multiplier};
  wire [5:0]   queue_dataIn_lo_lo_lo_15 = {queue_dataIn_lo_lo_lo_hi_15, queue_dataIn_lo_lo_lo_lo_15};
  wire         queue_15_enq_bits_decodeResult_unsigned1;
  wire         queue_15_enq_bits_decodeResult_unsigned0;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_15 = {queue_15_enq_bits_decodeResult_unsigned1, queue_15_enq_bits_decodeResult_unsigned0};
  wire         queue_15_enq_bits_decodeResult_other;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_15 = {queue_dataIn_lo_lo_hi_lo_hi_15, queue_15_enq_bits_decodeResult_other};
  wire         queue_15_enq_bits_decodeResult_red;
  wire         queue_15_enq_bits_decodeResult_nr;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_15 = {queue_15_enq_bits_decodeResult_red, queue_15_enq_bits_decodeResult_nr};
  wire         queue_15_enq_bits_decodeResult_itype;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_15 = {queue_dataIn_lo_lo_hi_hi_hi_15, queue_15_enq_bits_decodeResult_itype};
  wire [5:0]   queue_dataIn_lo_lo_hi_30 = {queue_dataIn_lo_lo_hi_hi_15, queue_dataIn_lo_lo_hi_lo_15};
  wire [11:0]  queue_dataIn_lo_lo_30 = {queue_dataIn_lo_lo_hi_30, queue_dataIn_lo_lo_lo_15};
  wire         queue_15_enq_bits_decodeResult_slid;
  wire         queue_15_enq_bits_decodeResult_targetRd;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_hi_15 = {queue_15_enq_bits_decodeResult_slid, queue_15_enq_bits_decodeResult_targetRd};
  wire         queue_15_enq_bits_decodeResult_widenReduce;
  wire [2:0]   queue_dataIn_lo_hi_lo_lo_15 = {queue_dataIn_lo_hi_lo_lo_hi_15, queue_15_enq_bits_decodeResult_widenReduce};
  wire         queue_15_enq_bits_decodeResult_compress;
  wire         queue_15_enq_bits_decodeResult_gather16;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_15 = {queue_15_enq_bits_decodeResult_compress, queue_15_enq_bits_decodeResult_gather16};
  wire         queue_15_enq_bits_decodeResult_gather;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_15 = {queue_dataIn_lo_hi_lo_hi_hi_15, queue_15_enq_bits_decodeResult_gather};
  wire [5:0]   queue_dataIn_lo_hi_lo_30 = {queue_dataIn_lo_hi_lo_hi_15, queue_dataIn_lo_hi_lo_lo_15};
  wire         queue_15_enq_bits_decodeResult_mv;
  wire         queue_15_enq_bits_decodeResult_extend;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_15 = {queue_15_enq_bits_decodeResult_mv, queue_15_enq_bits_decodeResult_extend};
  wire         queue_15_enq_bits_decodeResult_unOrderWrite;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_15 = {queue_dataIn_lo_hi_hi_lo_hi_15, queue_15_enq_bits_decodeResult_unOrderWrite};
  wire         queue_15_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_15_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_lo_hi_hi_hi_hi_15 = {queue_15_enq_bits_decodeResult_maskLogic, queue_15_enq_bits_decodeResult_uop};
  wire         queue_15_enq_bits_decodeResult_iota;
  wire [5:0]   queue_dataIn_lo_hi_hi_hi_15 = {queue_dataIn_lo_hi_hi_hi_hi_15, queue_15_enq_bits_decodeResult_iota};
  wire [8:0]   queue_dataIn_lo_hi_hi_30 = {queue_dataIn_lo_hi_hi_hi_15, queue_dataIn_lo_hi_hi_lo_15};
  wire [14:0]  queue_dataIn_lo_hi_46 = {queue_dataIn_lo_hi_hi_30, queue_dataIn_lo_hi_lo_30};
  wire [26:0]  queue_dataIn_lo_46 = {queue_dataIn_lo_hi_46, queue_dataIn_lo_lo_30};
  wire         queue_15_enq_bits_decodeResult_readOnly;
  wire         queue_15_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_lo_hi_15 = {queue_15_enq_bits_decodeResult_readOnly, queue_15_enq_bits_decodeResult_maskSource};
  wire         queue_15_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_lo_15 = {queue_dataIn_hi_lo_lo_lo_hi_15, queue_15_enq_bits_decodeResult_maskDestination};
  wire         queue_15_enq_bits_decodeResult_special;
  wire         queue_15_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_15 = {queue_15_enq_bits_decodeResult_special, queue_15_enq_bits_decodeResult_saturate};
  wire         queue_15_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_15 = {queue_dataIn_hi_lo_lo_hi_hi_15, queue_15_enq_bits_decodeResult_vwmacc};
  wire [5:0]   queue_dataIn_hi_lo_lo_30 = {queue_dataIn_hi_lo_lo_hi_15, queue_dataIn_hi_lo_lo_lo_15};
  wire         queue_15_enq_bits_decodeResult_crossRead;
  wire         queue_15_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_15 = {queue_15_enq_bits_decodeResult_crossRead, queue_15_enq_bits_decodeResult_crossWrite};
  wire         queue_15_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_15 = {queue_dataIn_hi_lo_hi_lo_hi_15, queue_15_enq_bits_decodeResult_maskUnit};
  wire         queue_15_enq_bits_decodeResult_sReadVD;
  wire         queue_15_enq_bits_decodeResult_vtype;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_15 = {queue_15_enq_bits_decodeResult_sReadVD, queue_15_enq_bits_decodeResult_vtype};
  wire         queue_15_enq_bits_decodeResult_sWrite;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_15 = {queue_dataIn_hi_lo_hi_hi_hi_15, queue_15_enq_bits_decodeResult_sWrite};
  wire [5:0]   queue_dataIn_hi_lo_hi_30 = {queue_dataIn_hi_lo_hi_hi_15, queue_dataIn_hi_lo_hi_lo_15};
  wire [11:0]  queue_dataIn_hi_lo_46 = {queue_dataIn_hi_lo_hi_30, queue_dataIn_hi_lo_lo_30};
  wire         queue_15_enq_bits_decodeResult_reverse;
  wire         queue_15_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_hi_15 = {queue_15_enq_bits_decodeResult_reverse, queue_15_enq_bits_decodeResult_dontNeedExecuteInLane};
  wire         queue_15_enq_bits_decodeResult_scheduler;
  wire [2:0]   queue_dataIn_hi_hi_lo_lo_15 = {queue_dataIn_hi_hi_lo_lo_hi_15, queue_15_enq_bits_decodeResult_scheduler};
  wire         queue_15_enq_bits_decodeResult_popCount;
  wire         queue_15_enq_bits_decodeResult_ffo;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_15 = {queue_15_enq_bits_decodeResult_popCount, queue_15_enq_bits_decodeResult_ffo};
  wire         queue_15_enq_bits_decodeResult_average;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_15 = {queue_dataIn_hi_hi_lo_hi_hi_15, queue_15_enq_bits_decodeResult_average};
  wire [5:0]   queue_dataIn_hi_hi_lo_30 = {queue_dataIn_hi_hi_lo_hi_15, queue_dataIn_hi_hi_lo_lo_15};
  wire         queue_15_enq_bits_decodeResult_float;
  wire         queue_15_enq_bits_decodeResult_specialSlot;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_15 = {queue_15_enq_bits_decodeResult_float, queue_15_enq_bits_decodeResult_specialSlot};
  wire [4:0]   queue_15_enq_bits_decodeResult_topUop;
  wire [6:0]   queue_dataIn_hi_hi_hi_lo_15 = {queue_dataIn_hi_hi_hi_lo_hi_15, queue_15_enq_bits_decodeResult_topUop};
  wire         queue_15_enq_bits_decodeResult_orderReduce;
  wire         queue_15_enq_bits_decodeResult_floatMul;
  wire [1:0]   queue_dataIn_hi_hi_hi_hi_hi_15 = {queue_15_enq_bits_decodeResult_orderReduce, queue_15_enq_bits_decodeResult_floatMul};
  wire [1:0]   queue_15_enq_bits_decodeResult_fpExecutionType;
  wire [3:0]   queue_dataIn_hi_hi_hi_hi_15 = {queue_dataIn_hi_hi_hi_hi_hi_15, queue_15_enq_bits_decodeResult_fpExecutionType};
  wire [10:0]  queue_dataIn_hi_hi_hi_30 = {queue_dataIn_hi_hi_hi_hi_15, queue_dataIn_hi_hi_hi_lo_15};
  wire [16:0]  queue_dataIn_hi_hi_46 = {queue_dataIn_hi_hi_hi_30, queue_dataIn_hi_hi_lo_30};
  wire [28:0]  queue_dataIn_hi_46 = {queue_dataIn_hi_hi_46, queue_dataIn_hi_lo_46};
  wire [2:0]   queue_15_enq_bits_segment;
  wire [31:0]  queue_15_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_31 = {queue_15_enq_bits_segment, queue_15_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_31 = {queue_dataIn_lo_lo_hi_31, queue_dataIn_hi_45, queue_dataIn_lo_45};
  wire [1:0]   queue_15_enq_bits_loadStoreEEW;
  wire         queue_15_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_31 = {queue_15_enq_bits_loadStoreEEW, queue_15_enq_bits_mask};
  wire [4:0]   queue_15_enq_bits_vs2;
  wire [4:0]   queue_15_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_31 = {queue_15_enq_bits_vs2, queue_15_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_47 = {queue_dataIn_lo_hi_hi_31, queue_dataIn_lo_hi_lo_31};
  wire [80:0]  queue_dataIn_lo_47 = {queue_dataIn_lo_hi_47, queue_dataIn_lo_lo_31};
  wire         queue_15_enq_bits_lsWholeReg;
  wire [4:0]   queue_15_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_31 = {queue_15_enq_bits_lsWholeReg, queue_15_enq_bits_vs1};
  wire         queue_15_enq_bits_store;
  wire         queue_15_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_31 = {queue_15_enq_bits_store, queue_15_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_47 = {queue_dataIn_hi_lo_hi_31, queue_dataIn_hi_lo_lo_31};
  wire         queue_15_enq_bits_loadStore;
  wire         queue_15_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_31 = {queue_15_enq_bits_loadStore, queue_15_enq_bits_issueInst};
  wire [2:0]   queue_15_enq_bits_instructionIndex;
  wire [58:0]  queue_dataIn_hi_hi_hi_31 = {queue_15_enq_bits_instructionIndex, queue_dataIn_hi_46, queue_dataIn_lo_46};
  wire [60:0]  queue_dataIn_hi_hi_47 = {queue_dataIn_hi_hi_hi_31, queue_dataIn_hi_hi_lo_31};
  wire [68:0]  queue_dataIn_hi_47 = {queue_dataIn_hi_hi_47, queue_dataIn_hi_lo_47};
  wire [149:0] queue_dataIn_15 = {queue_dataIn_hi_47, queue_dataIn_lo_47};
  wire         queue_dataOut_15_csrInterface_vma = _queue_fifo_15_data_out[0];
  wire         queue_dataOut_15_csrInterface_vta = _queue_fifo_15_data_out[1];
  wire [1:0]   queue_dataOut_15_csrInterface_vxrm = _queue_fifo_15_data_out[3:2];
  wire [1:0]   queue_dataOut_15_csrInterface_vSew = _queue_fifo_15_data_out[5:4];
  wire [2:0]   queue_dataOut_15_csrInterface_vlmul = _queue_fifo_15_data_out[8:6];
  wire [11:0]  queue_dataOut_15_csrInterface_vStart = _queue_fifo_15_data_out[20:9];
  wire [11:0]  queue_dataOut_15_csrInterface_vl = _queue_fifo_15_data_out[32:21];
  wire [31:0]  queue_dataOut_15_readFromScalar = _queue_fifo_15_data_out[64:33];
  wire [2:0]   queue_dataOut_15_segment = _queue_fifo_15_data_out[67:65];
  wire         queue_dataOut_15_mask = _queue_fifo_15_data_out[68];
  wire [1:0]   queue_dataOut_15_loadStoreEEW = _queue_fifo_15_data_out[70:69];
  wire [4:0]   queue_dataOut_15_vd = _queue_fifo_15_data_out[75:71];
  wire [4:0]   queue_dataOut_15_vs2 = _queue_fifo_15_data_out[80:76];
  wire [4:0]   queue_dataOut_15_vs1 = _queue_fifo_15_data_out[85:81];
  wire         queue_dataOut_15_lsWholeReg = _queue_fifo_15_data_out[86];
  wire         queue_dataOut_15_special = _queue_fifo_15_data_out[87];
  wire         queue_dataOut_15_store = _queue_fifo_15_data_out[88];
  wire         queue_dataOut_15_issueInst = _queue_fifo_15_data_out[89];
  wire         queue_dataOut_15_loadStore = _queue_fifo_15_data_out[90];
  wire         queue_dataOut_15_decodeResult_logic = _queue_fifo_15_data_out[91];
  wire         queue_dataOut_15_decodeResult_adder = _queue_fifo_15_data_out[92];
  wire         queue_dataOut_15_decodeResult_shift = _queue_fifo_15_data_out[93];
  wire         queue_dataOut_15_decodeResult_multiplier = _queue_fifo_15_data_out[94];
  wire         queue_dataOut_15_decodeResult_divider = _queue_fifo_15_data_out[95];
  wire         queue_dataOut_15_decodeResult_multiCycle = _queue_fifo_15_data_out[96];
  wire         queue_dataOut_15_decodeResult_other = _queue_fifo_15_data_out[97];
  wire         queue_dataOut_15_decodeResult_unsigned0 = _queue_fifo_15_data_out[98];
  wire         queue_dataOut_15_decodeResult_unsigned1 = _queue_fifo_15_data_out[99];
  wire         queue_dataOut_15_decodeResult_itype = _queue_fifo_15_data_out[100];
  wire         queue_dataOut_15_decodeResult_nr = _queue_fifo_15_data_out[101];
  wire         queue_dataOut_15_decodeResult_red = _queue_fifo_15_data_out[102];
  wire         queue_dataOut_15_decodeResult_widenReduce = _queue_fifo_15_data_out[103];
  wire         queue_dataOut_15_decodeResult_targetRd = _queue_fifo_15_data_out[104];
  wire         queue_dataOut_15_decodeResult_slid = _queue_fifo_15_data_out[105];
  wire         queue_dataOut_15_decodeResult_gather = _queue_fifo_15_data_out[106];
  wire         queue_dataOut_15_decodeResult_gather16 = _queue_fifo_15_data_out[107];
  wire         queue_dataOut_15_decodeResult_compress = _queue_fifo_15_data_out[108];
  wire         queue_dataOut_15_decodeResult_unOrderWrite = _queue_fifo_15_data_out[109];
  wire         queue_dataOut_15_decodeResult_extend = _queue_fifo_15_data_out[110];
  wire         queue_dataOut_15_decodeResult_mv = _queue_fifo_15_data_out[111];
  wire         queue_dataOut_15_decodeResult_iota = _queue_fifo_15_data_out[112];
  wire [3:0]   queue_dataOut_15_decodeResult_uop = _queue_fifo_15_data_out[116:113];
  wire         queue_dataOut_15_decodeResult_maskLogic = _queue_fifo_15_data_out[117];
  wire         queue_dataOut_15_decodeResult_maskDestination = _queue_fifo_15_data_out[118];
  wire         queue_dataOut_15_decodeResult_maskSource = _queue_fifo_15_data_out[119];
  wire         queue_dataOut_15_decodeResult_readOnly = _queue_fifo_15_data_out[120];
  wire         queue_dataOut_15_decodeResult_vwmacc = _queue_fifo_15_data_out[121];
  wire         queue_dataOut_15_decodeResult_saturate = _queue_fifo_15_data_out[122];
  wire         queue_dataOut_15_decodeResult_special = _queue_fifo_15_data_out[123];
  wire         queue_dataOut_15_decodeResult_maskUnit = _queue_fifo_15_data_out[124];
  wire         queue_dataOut_15_decodeResult_crossWrite = _queue_fifo_15_data_out[125];
  wire         queue_dataOut_15_decodeResult_crossRead = _queue_fifo_15_data_out[126];
  wire         queue_dataOut_15_decodeResult_sWrite = _queue_fifo_15_data_out[127];
  wire         queue_dataOut_15_decodeResult_vtype = _queue_fifo_15_data_out[128];
  wire         queue_dataOut_15_decodeResult_sReadVD = _queue_fifo_15_data_out[129];
  wire         queue_dataOut_15_decodeResult_scheduler = _queue_fifo_15_data_out[130];
  wire         queue_dataOut_15_decodeResult_dontNeedExecuteInLane = _queue_fifo_15_data_out[131];
  wire         queue_dataOut_15_decodeResult_reverse = _queue_fifo_15_data_out[132];
  wire         queue_dataOut_15_decodeResult_average = _queue_fifo_15_data_out[133];
  wire         queue_dataOut_15_decodeResult_ffo = _queue_fifo_15_data_out[134];
  wire         queue_dataOut_15_decodeResult_popCount = _queue_fifo_15_data_out[135];
  wire [4:0]   queue_dataOut_15_decodeResult_topUop = _queue_fifo_15_data_out[140:136];
  wire         queue_dataOut_15_decodeResult_specialSlot = _queue_fifo_15_data_out[141];
  wire         queue_dataOut_15_decodeResult_float = _queue_fifo_15_data_out[142];
  wire [1:0]   queue_dataOut_15_decodeResult_fpExecutionType = _queue_fifo_15_data_out[144:143];
  wire         queue_dataOut_15_decodeResult_floatMul = _queue_fifo_15_data_out[145];
  wire         queue_dataOut_15_decodeResult_orderReduce = _queue_fifo_15_data_out[146];
  wire [2:0]   queue_dataOut_15_instructionIndex = _queue_fifo_15_data_out[149:147];
  wire         queue_15_enq_ready = ~_queue_fifo_15_full;
  wire         queue_15_enq_valid;
  assign queue_15_deq_valid = ~_queue_fifo_15_empty | queue_15_enq_valid;
  assign queue_15_deq_bits_instructionIndex = _queue_fifo_15_empty ? queue_15_enq_bits_instructionIndex : queue_dataOut_15_instructionIndex;
  assign queue_15_deq_bits_decodeResult_orderReduce = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_orderReduce : queue_dataOut_15_decodeResult_orderReduce;
  assign queue_15_deq_bits_decodeResult_floatMul = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_floatMul : queue_dataOut_15_decodeResult_floatMul;
  assign queue_15_deq_bits_decodeResult_fpExecutionType = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_fpExecutionType : queue_dataOut_15_decodeResult_fpExecutionType;
  assign queue_15_deq_bits_decodeResult_float = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_float : queue_dataOut_15_decodeResult_float;
  assign queue_15_deq_bits_decodeResult_specialSlot = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_specialSlot : queue_dataOut_15_decodeResult_specialSlot;
  assign queue_15_deq_bits_decodeResult_topUop = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_topUop : queue_dataOut_15_decodeResult_topUop;
  assign queue_15_deq_bits_decodeResult_popCount = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_popCount : queue_dataOut_15_decodeResult_popCount;
  assign queue_15_deq_bits_decodeResult_ffo = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_ffo : queue_dataOut_15_decodeResult_ffo;
  assign queue_15_deq_bits_decodeResult_average = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_average : queue_dataOut_15_decodeResult_average;
  assign queue_15_deq_bits_decodeResult_reverse = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_reverse : queue_dataOut_15_decodeResult_reverse;
  assign queue_15_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_15_decodeResult_dontNeedExecuteInLane;
  assign queue_15_deq_bits_decodeResult_scheduler = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_scheduler : queue_dataOut_15_decodeResult_scheduler;
  assign queue_15_deq_bits_decodeResult_sReadVD = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_sReadVD : queue_dataOut_15_decodeResult_sReadVD;
  assign queue_15_deq_bits_decodeResult_vtype = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_vtype : queue_dataOut_15_decodeResult_vtype;
  assign queue_15_deq_bits_decodeResult_sWrite = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_sWrite : queue_dataOut_15_decodeResult_sWrite;
  assign queue_15_deq_bits_decodeResult_crossRead = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_crossRead : queue_dataOut_15_decodeResult_crossRead;
  assign queue_15_deq_bits_decodeResult_crossWrite = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_crossWrite : queue_dataOut_15_decodeResult_crossWrite;
  assign queue_15_deq_bits_decodeResult_maskUnit = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_maskUnit : queue_dataOut_15_decodeResult_maskUnit;
  assign queue_15_deq_bits_decodeResult_special = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_special : queue_dataOut_15_decodeResult_special;
  assign queue_15_deq_bits_decodeResult_saturate = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_saturate : queue_dataOut_15_decodeResult_saturate;
  assign queue_15_deq_bits_decodeResult_vwmacc = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_vwmacc : queue_dataOut_15_decodeResult_vwmacc;
  assign queue_15_deq_bits_decodeResult_readOnly = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_readOnly : queue_dataOut_15_decodeResult_readOnly;
  assign queue_15_deq_bits_decodeResult_maskSource = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_maskSource : queue_dataOut_15_decodeResult_maskSource;
  assign queue_15_deq_bits_decodeResult_maskDestination = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_maskDestination : queue_dataOut_15_decodeResult_maskDestination;
  assign queue_15_deq_bits_decodeResult_maskLogic = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_maskLogic : queue_dataOut_15_decodeResult_maskLogic;
  assign queue_15_deq_bits_decodeResult_uop = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_uop : queue_dataOut_15_decodeResult_uop;
  assign queue_15_deq_bits_decodeResult_iota = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_iota : queue_dataOut_15_decodeResult_iota;
  assign queue_15_deq_bits_decodeResult_mv = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_mv : queue_dataOut_15_decodeResult_mv;
  assign queue_15_deq_bits_decodeResult_extend = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_extend : queue_dataOut_15_decodeResult_extend;
  assign queue_15_deq_bits_decodeResult_unOrderWrite = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_unOrderWrite : queue_dataOut_15_decodeResult_unOrderWrite;
  assign queue_15_deq_bits_decodeResult_compress = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_compress : queue_dataOut_15_decodeResult_compress;
  assign queue_15_deq_bits_decodeResult_gather16 = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_gather16 : queue_dataOut_15_decodeResult_gather16;
  assign queue_15_deq_bits_decodeResult_gather = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_gather : queue_dataOut_15_decodeResult_gather;
  assign queue_15_deq_bits_decodeResult_slid = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_slid : queue_dataOut_15_decodeResult_slid;
  assign queue_15_deq_bits_decodeResult_targetRd = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_targetRd : queue_dataOut_15_decodeResult_targetRd;
  assign queue_15_deq_bits_decodeResult_widenReduce = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_widenReduce : queue_dataOut_15_decodeResult_widenReduce;
  assign queue_15_deq_bits_decodeResult_red = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_red : queue_dataOut_15_decodeResult_red;
  assign queue_15_deq_bits_decodeResult_nr = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_nr : queue_dataOut_15_decodeResult_nr;
  assign queue_15_deq_bits_decodeResult_itype = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_itype : queue_dataOut_15_decodeResult_itype;
  assign queue_15_deq_bits_decodeResult_unsigned1 = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_unsigned1 : queue_dataOut_15_decodeResult_unsigned1;
  assign queue_15_deq_bits_decodeResult_unsigned0 = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_unsigned0 : queue_dataOut_15_decodeResult_unsigned0;
  assign queue_15_deq_bits_decodeResult_other = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_other : queue_dataOut_15_decodeResult_other;
  assign queue_15_deq_bits_decodeResult_multiCycle = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_multiCycle : queue_dataOut_15_decodeResult_multiCycle;
  assign queue_15_deq_bits_decodeResult_divider = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_divider : queue_dataOut_15_decodeResult_divider;
  assign queue_15_deq_bits_decodeResult_multiplier = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_multiplier : queue_dataOut_15_decodeResult_multiplier;
  assign queue_15_deq_bits_decodeResult_shift = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_shift : queue_dataOut_15_decodeResult_shift;
  assign queue_15_deq_bits_decodeResult_adder = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_adder : queue_dataOut_15_decodeResult_adder;
  assign queue_15_deq_bits_decodeResult_logic = _queue_fifo_15_empty ? queue_15_enq_bits_decodeResult_logic : queue_dataOut_15_decodeResult_logic;
  assign queue_15_deq_bits_loadStore = _queue_fifo_15_empty ? queue_15_enq_bits_loadStore : queue_dataOut_15_loadStore;
  assign queue_15_deq_bits_issueInst = _queue_fifo_15_empty ? queue_15_enq_bits_issueInst : queue_dataOut_15_issueInst;
  assign queue_15_deq_bits_store = _queue_fifo_15_empty ? queue_15_enq_bits_store : queue_dataOut_15_store;
  assign queue_15_deq_bits_special = _queue_fifo_15_empty ? queue_15_enq_bits_special : queue_dataOut_15_special;
  assign queue_15_deq_bits_lsWholeReg = _queue_fifo_15_empty ? queue_15_enq_bits_lsWholeReg : queue_dataOut_15_lsWholeReg;
  assign queue_15_deq_bits_vs1 = _queue_fifo_15_empty ? queue_15_enq_bits_vs1 : queue_dataOut_15_vs1;
  assign queue_15_deq_bits_vs2 = _queue_fifo_15_empty ? queue_15_enq_bits_vs2 : queue_dataOut_15_vs2;
  assign queue_15_deq_bits_vd = _queue_fifo_15_empty ? queue_15_enq_bits_vd : queue_dataOut_15_vd;
  assign queue_15_deq_bits_loadStoreEEW = _queue_fifo_15_empty ? queue_15_enq_bits_loadStoreEEW : queue_dataOut_15_loadStoreEEW;
  assign queue_15_deq_bits_mask = _queue_fifo_15_empty ? queue_15_enq_bits_mask : queue_dataOut_15_mask;
  assign queue_15_deq_bits_segment = _queue_fifo_15_empty ? queue_15_enq_bits_segment : queue_dataOut_15_segment;
  assign queue_15_deq_bits_readFromScalar = _queue_fifo_15_empty ? queue_15_enq_bits_readFromScalar : queue_dataOut_15_readFromScalar;
  assign queue_15_deq_bits_csrInterface_vl = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vl : queue_dataOut_15_csrInterface_vl;
  assign queue_15_deq_bits_csrInterface_vStart = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vStart : queue_dataOut_15_csrInterface_vStart;
  assign queue_15_deq_bits_csrInterface_vlmul = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vlmul : queue_dataOut_15_csrInterface_vlmul;
  assign queue_15_deq_bits_csrInterface_vSew = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vSew : queue_dataOut_15_csrInterface_vSew;
  assign queue_15_deq_bits_csrInterface_vxrm = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vxrm : queue_dataOut_15_csrInterface_vxrm;
  assign queue_15_deq_bits_csrInterface_vta = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vta : queue_dataOut_15_csrInterface_vta;
  assign queue_15_deq_bits_csrInterface_vma = _queue_fifo_15_empty ? queue_15_enq_bits_csrInterface_vma : queue_dataOut_15_csrInterface_vma;
  wire         laneVec_15_laneRequest_bits_issueInst = laneRequestSinkWire_15_ready & laneRequestSinkWire_15_valid;
  reg          releasePipe_pipe_v_15;
  wire         releasePipe_pipe_out_15_valid = releasePipe_pipe_v_15;
  wire         laneRequestSourceWire_15_ready;
  wire         validSource_15_valid = laneRequestSourceWire_15_ready & laneRequestSourceWire_15_valid;
  reg  [2:0]   tokenCheck_counter_15;
  wire [2:0]   tokenCheck_counterChange_15 = validSource_15_valid ? 3'h1 : 3'h7;
  assign tokenCheck_15 = ~(tokenCheck_counter_15[2]);
  assign laneRequestSourceWire_15_ready = tokenCheck_15;
  assign queue_15_enq_valid = validSink_15_valid;
  assign queue_15_enq_bits_instructionIndex = validSink_15_bits_instructionIndex;
  assign queue_15_enq_bits_decodeResult_orderReduce = validSink_15_bits_decodeResult_orderReduce;
  assign queue_15_enq_bits_decodeResult_floatMul = validSink_15_bits_decodeResult_floatMul;
  assign queue_15_enq_bits_decodeResult_fpExecutionType = validSink_15_bits_decodeResult_fpExecutionType;
  assign queue_15_enq_bits_decodeResult_float = validSink_15_bits_decodeResult_float;
  assign queue_15_enq_bits_decodeResult_specialSlot = validSink_15_bits_decodeResult_specialSlot;
  assign queue_15_enq_bits_decodeResult_topUop = validSink_15_bits_decodeResult_topUop;
  assign queue_15_enq_bits_decodeResult_popCount = validSink_15_bits_decodeResult_popCount;
  assign queue_15_enq_bits_decodeResult_ffo = validSink_15_bits_decodeResult_ffo;
  assign queue_15_enq_bits_decodeResult_average = validSink_15_bits_decodeResult_average;
  assign queue_15_enq_bits_decodeResult_reverse = validSink_15_bits_decodeResult_reverse;
  assign queue_15_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_15_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_15_enq_bits_decodeResult_scheduler = validSink_15_bits_decodeResult_scheduler;
  assign queue_15_enq_bits_decodeResult_sReadVD = validSink_15_bits_decodeResult_sReadVD;
  assign queue_15_enq_bits_decodeResult_vtype = validSink_15_bits_decodeResult_vtype;
  assign queue_15_enq_bits_decodeResult_sWrite = validSink_15_bits_decodeResult_sWrite;
  assign queue_15_enq_bits_decodeResult_crossRead = validSink_15_bits_decodeResult_crossRead;
  assign queue_15_enq_bits_decodeResult_crossWrite = validSink_15_bits_decodeResult_crossWrite;
  assign queue_15_enq_bits_decodeResult_maskUnit = validSink_15_bits_decodeResult_maskUnit;
  assign queue_15_enq_bits_decodeResult_special = validSink_15_bits_decodeResult_special;
  assign queue_15_enq_bits_decodeResult_saturate = validSink_15_bits_decodeResult_saturate;
  assign queue_15_enq_bits_decodeResult_vwmacc = validSink_15_bits_decodeResult_vwmacc;
  assign queue_15_enq_bits_decodeResult_readOnly = validSink_15_bits_decodeResult_readOnly;
  assign queue_15_enq_bits_decodeResult_maskSource = validSink_15_bits_decodeResult_maskSource;
  assign queue_15_enq_bits_decodeResult_maskDestination = validSink_15_bits_decodeResult_maskDestination;
  assign queue_15_enq_bits_decodeResult_maskLogic = validSink_15_bits_decodeResult_maskLogic;
  assign queue_15_enq_bits_decodeResult_uop = validSink_15_bits_decodeResult_uop;
  assign queue_15_enq_bits_decodeResult_iota = validSink_15_bits_decodeResult_iota;
  assign queue_15_enq_bits_decodeResult_mv = validSink_15_bits_decodeResult_mv;
  assign queue_15_enq_bits_decodeResult_extend = validSink_15_bits_decodeResult_extend;
  assign queue_15_enq_bits_decodeResult_unOrderWrite = validSink_15_bits_decodeResult_unOrderWrite;
  assign queue_15_enq_bits_decodeResult_compress = validSink_15_bits_decodeResult_compress;
  assign queue_15_enq_bits_decodeResult_gather16 = validSink_15_bits_decodeResult_gather16;
  assign queue_15_enq_bits_decodeResult_gather = validSink_15_bits_decodeResult_gather;
  assign queue_15_enq_bits_decodeResult_slid = validSink_15_bits_decodeResult_slid;
  assign queue_15_enq_bits_decodeResult_targetRd = validSink_15_bits_decodeResult_targetRd;
  assign queue_15_enq_bits_decodeResult_widenReduce = validSink_15_bits_decodeResult_widenReduce;
  assign queue_15_enq_bits_decodeResult_red = validSink_15_bits_decodeResult_red;
  assign queue_15_enq_bits_decodeResult_nr = validSink_15_bits_decodeResult_nr;
  assign queue_15_enq_bits_decodeResult_itype = validSink_15_bits_decodeResult_itype;
  assign queue_15_enq_bits_decodeResult_unsigned1 = validSink_15_bits_decodeResult_unsigned1;
  assign queue_15_enq_bits_decodeResult_unsigned0 = validSink_15_bits_decodeResult_unsigned0;
  assign queue_15_enq_bits_decodeResult_other = validSink_15_bits_decodeResult_other;
  assign queue_15_enq_bits_decodeResult_multiCycle = validSink_15_bits_decodeResult_multiCycle;
  assign queue_15_enq_bits_decodeResult_divider = validSink_15_bits_decodeResult_divider;
  assign queue_15_enq_bits_decodeResult_multiplier = validSink_15_bits_decodeResult_multiplier;
  assign queue_15_enq_bits_decodeResult_shift = validSink_15_bits_decodeResult_shift;
  assign queue_15_enq_bits_decodeResult_adder = validSink_15_bits_decodeResult_adder;
  assign queue_15_enq_bits_decodeResult_logic = validSink_15_bits_decodeResult_logic;
  assign queue_15_enq_bits_loadStore = validSink_15_bits_loadStore;
  assign queue_15_enq_bits_issueInst = validSink_15_bits_issueInst;
  assign queue_15_enq_bits_store = validSink_15_bits_store;
  assign queue_15_enq_bits_special = validSink_15_bits_special;
  assign queue_15_enq_bits_lsWholeReg = validSink_15_bits_lsWholeReg;
  assign queue_15_enq_bits_vs1 = validSink_15_bits_vs1;
  assign queue_15_enq_bits_vs2 = validSink_15_bits_vs2;
  assign queue_15_enq_bits_vd = validSink_15_bits_vd;
  assign queue_15_enq_bits_loadStoreEEW = validSink_15_bits_loadStoreEEW;
  assign queue_15_enq_bits_mask = validSink_15_bits_mask;
  assign queue_15_enq_bits_segment = validSink_15_bits_segment;
  assign queue_15_enq_bits_readFromScalar = validSink_15_bits_readFromScalar;
  assign queue_15_enq_bits_csrInterface_vl = validSink_15_bits_csrInterface_vl;
  assign queue_15_enq_bits_csrInterface_vStart = validSink_15_bits_csrInterface_vStart;
  assign queue_15_enq_bits_csrInterface_vlmul = validSink_15_bits_csrInterface_vlmul;
  assign queue_15_enq_bits_csrInterface_vSew = validSink_15_bits_csrInterface_vSew;
  assign queue_15_enq_bits_csrInterface_vxrm = validSink_15_bits_csrInterface_vxrm;
  assign queue_15_enq_bits_csrInterface_vta = validSink_15_bits_csrInterface_vta;
  assign queue_15_enq_bits_csrInterface_vma = validSink_15_bits_csrInterface_vma;
  reg          shifterReg_15_0_valid;
  assign validSink_15_valid = shifterReg_15_0_valid;
  reg  [2:0]   shifterReg_15_0_bits_instructionIndex;
  assign validSink_15_bits_instructionIndex = shifterReg_15_0_bits_instructionIndex;
  reg          shifterReg_15_0_bits_decodeResult_orderReduce;
  assign validSink_15_bits_decodeResult_orderReduce = shifterReg_15_0_bits_decodeResult_orderReduce;
  reg          shifterReg_15_0_bits_decodeResult_floatMul;
  assign validSink_15_bits_decodeResult_floatMul = shifterReg_15_0_bits_decodeResult_floatMul;
  reg  [1:0]   shifterReg_15_0_bits_decodeResult_fpExecutionType;
  assign validSink_15_bits_decodeResult_fpExecutionType = shifterReg_15_0_bits_decodeResult_fpExecutionType;
  reg          shifterReg_15_0_bits_decodeResult_float;
  assign validSink_15_bits_decodeResult_float = shifterReg_15_0_bits_decodeResult_float;
  reg          shifterReg_15_0_bits_decodeResult_specialSlot;
  assign validSink_15_bits_decodeResult_specialSlot = shifterReg_15_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_15_0_bits_decodeResult_topUop;
  assign validSink_15_bits_decodeResult_topUop = shifterReg_15_0_bits_decodeResult_topUop;
  reg          shifterReg_15_0_bits_decodeResult_popCount;
  assign validSink_15_bits_decodeResult_popCount = shifterReg_15_0_bits_decodeResult_popCount;
  reg          shifterReg_15_0_bits_decodeResult_ffo;
  assign validSink_15_bits_decodeResult_ffo = shifterReg_15_0_bits_decodeResult_ffo;
  reg          shifterReg_15_0_bits_decodeResult_average;
  assign validSink_15_bits_decodeResult_average = shifterReg_15_0_bits_decodeResult_average;
  reg          shifterReg_15_0_bits_decodeResult_reverse;
  assign validSink_15_bits_decodeResult_reverse = shifterReg_15_0_bits_decodeResult_reverse;
  reg          shifterReg_15_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_15_bits_decodeResult_dontNeedExecuteInLane = shifterReg_15_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_15_0_bits_decodeResult_scheduler;
  assign validSink_15_bits_decodeResult_scheduler = shifterReg_15_0_bits_decodeResult_scheduler;
  reg          shifterReg_15_0_bits_decodeResult_sReadVD;
  assign validSink_15_bits_decodeResult_sReadVD = shifterReg_15_0_bits_decodeResult_sReadVD;
  reg          shifterReg_15_0_bits_decodeResult_vtype;
  assign validSink_15_bits_decodeResult_vtype = shifterReg_15_0_bits_decodeResult_vtype;
  reg          shifterReg_15_0_bits_decodeResult_sWrite;
  assign validSink_15_bits_decodeResult_sWrite = shifterReg_15_0_bits_decodeResult_sWrite;
  reg          shifterReg_15_0_bits_decodeResult_crossRead;
  assign validSink_15_bits_decodeResult_crossRead = shifterReg_15_0_bits_decodeResult_crossRead;
  reg          shifterReg_15_0_bits_decodeResult_crossWrite;
  assign validSink_15_bits_decodeResult_crossWrite = shifterReg_15_0_bits_decodeResult_crossWrite;
  reg          shifterReg_15_0_bits_decodeResult_maskUnit;
  assign validSink_15_bits_decodeResult_maskUnit = shifterReg_15_0_bits_decodeResult_maskUnit;
  reg          shifterReg_15_0_bits_decodeResult_special;
  assign validSink_15_bits_decodeResult_special = shifterReg_15_0_bits_decodeResult_special;
  reg          shifterReg_15_0_bits_decodeResult_saturate;
  assign validSink_15_bits_decodeResult_saturate = shifterReg_15_0_bits_decodeResult_saturate;
  reg          shifterReg_15_0_bits_decodeResult_vwmacc;
  assign validSink_15_bits_decodeResult_vwmacc = shifterReg_15_0_bits_decodeResult_vwmacc;
  reg          shifterReg_15_0_bits_decodeResult_readOnly;
  assign validSink_15_bits_decodeResult_readOnly = shifterReg_15_0_bits_decodeResult_readOnly;
  reg          shifterReg_15_0_bits_decodeResult_maskSource;
  assign validSink_15_bits_decodeResult_maskSource = shifterReg_15_0_bits_decodeResult_maskSource;
  reg          shifterReg_15_0_bits_decodeResult_maskDestination;
  assign validSink_15_bits_decodeResult_maskDestination = shifterReg_15_0_bits_decodeResult_maskDestination;
  reg          shifterReg_15_0_bits_decodeResult_maskLogic;
  assign validSink_15_bits_decodeResult_maskLogic = shifterReg_15_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_15_0_bits_decodeResult_uop;
  assign validSink_15_bits_decodeResult_uop = shifterReg_15_0_bits_decodeResult_uop;
  reg          shifterReg_15_0_bits_decodeResult_iota;
  assign validSink_15_bits_decodeResult_iota = shifterReg_15_0_bits_decodeResult_iota;
  reg          shifterReg_15_0_bits_decodeResult_mv;
  assign validSink_15_bits_decodeResult_mv = shifterReg_15_0_bits_decodeResult_mv;
  reg          shifterReg_15_0_bits_decodeResult_extend;
  assign validSink_15_bits_decodeResult_extend = shifterReg_15_0_bits_decodeResult_extend;
  reg          shifterReg_15_0_bits_decodeResult_unOrderWrite;
  assign validSink_15_bits_decodeResult_unOrderWrite = shifterReg_15_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_15_0_bits_decodeResult_compress;
  assign validSink_15_bits_decodeResult_compress = shifterReg_15_0_bits_decodeResult_compress;
  reg          shifterReg_15_0_bits_decodeResult_gather16;
  assign validSink_15_bits_decodeResult_gather16 = shifterReg_15_0_bits_decodeResult_gather16;
  reg          shifterReg_15_0_bits_decodeResult_gather;
  assign validSink_15_bits_decodeResult_gather = shifterReg_15_0_bits_decodeResult_gather;
  reg          shifterReg_15_0_bits_decodeResult_slid;
  assign validSink_15_bits_decodeResult_slid = shifterReg_15_0_bits_decodeResult_slid;
  reg          shifterReg_15_0_bits_decodeResult_targetRd;
  assign validSink_15_bits_decodeResult_targetRd = shifterReg_15_0_bits_decodeResult_targetRd;
  reg          shifterReg_15_0_bits_decodeResult_widenReduce;
  assign validSink_15_bits_decodeResult_widenReduce = shifterReg_15_0_bits_decodeResult_widenReduce;
  reg          shifterReg_15_0_bits_decodeResult_red;
  assign validSink_15_bits_decodeResult_red = shifterReg_15_0_bits_decodeResult_red;
  reg          shifterReg_15_0_bits_decodeResult_nr;
  assign validSink_15_bits_decodeResult_nr = shifterReg_15_0_bits_decodeResult_nr;
  reg          shifterReg_15_0_bits_decodeResult_itype;
  assign validSink_15_bits_decodeResult_itype = shifterReg_15_0_bits_decodeResult_itype;
  reg          shifterReg_15_0_bits_decodeResult_unsigned1;
  assign validSink_15_bits_decodeResult_unsigned1 = shifterReg_15_0_bits_decodeResult_unsigned1;
  reg          shifterReg_15_0_bits_decodeResult_unsigned0;
  assign validSink_15_bits_decodeResult_unsigned0 = shifterReg_15_0_bits_decodeResult_unsigned0;
  reg          shifterReg_15_0_bits_decodeResult_other;
  assign validSink_15_bits_decodeResult_other = shifterReg_15_0_bits_decodeResult_other;
  reg          shifterReg_15_0_bits_decodeResult_multiCycle;
  assign validSink_15_bits_decodeResult_multiCycle = shifterReg_15_0_bits_decodeResult_multiCycle;
  reg          shifterReg_15_0_bits_decodeResult_divider;
  assign validSink_15_bits_decodeResult_divider = shifterReg_15_0_bits_decodeResult_divider;
  reg          shifterReg_15_0_bits_decodeResult_multiplier;
  assign validSink_15_bits_decodeResult_multiplier = shifterReg_15_0_bits_decodeResult_multiplier;
  reg          shifterReg_15_0_bits_decodeResult_shift;
  assign validSink_15_bits_decodeResult_shift = shifterReg_15_0_bits_decodeResult_shift;
  reg          shifterReg_15_0_bits_decodeResult_adder;
  assign validSink_15_bits_decodeResult_adder = shifterReg_15_0_bits_decodeResult_adder;
  reg          shifterReg_15_0_bits_decodeResult_logic;
  assign validSink_15_bits_decodeResult_logic = shifterReg_15_0_bits_decodeResult_logic;
  reg          shifterReg_15_0_bits_loadStore;
  assign validSink_15_bits_loadStore = shifterReg_15_0_bits_loadStore;
  reg          shifterReg_15_0_bits_issueInst;
  assign validSink_15_bits_issueInst = shifterReg_15_0_bits_issueInst;
  reg          shifterReg_15_0_bits_store;
  assign validSink_15_bits_store = shifterReg_15_0_bits_store;
  reg          shifterReg_15_0_bits_special;
  assign validSink_15_bits_special = shifterReg_15_0_bits_special;
  reg          shifterReg_15_0_bits_lsWholeReg;
  assign validSink_15_bits_lsWholeReg = shifterReg_15_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_15_0_bits_vs1;
  assign validSink_15_bits_vs1 = shifterReg_15_0_bits_vs1;
  reg  [4:0]   shifterReg_15_0_bits_vs2;
  assign validSink_15_bits_vs2 = shifterReg_15_0_bits_vs2;
  reg  [4:0]   shifterReg_15_0_bits_vd;
  assign validSink_15_bits_vd = shifterReg_15_0_bits_vd;
  reg  [1:0]   shifterReg_15_0_bits_loadStoreEEW;
  assign validSink_15_bits_loadStoreEEW = shifterReg_15_0_bits_loadStoreEEW;
  reg          shifterReg_15_0_bits_mask;
  assign validSink_15_bits_mask = shifterReg_15_0_bits_mask;
  reg  [2:0]   shifterReg_15_0_bits_segment;
  assign validSink_15_bits_segment = shifterReg_15_0_bits_segment;
  reg  [31:0]  shifterReg_15_0_bits_readFromScalar;
  assign validSink_15_bits_readFromScalar = shifterReg_15_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_15_0_bits_csrInterface_vl;
  assign validSink_15_bits_csrInterface_vl = shifterReg_15_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_15_0_bits_csrInterface_vStart;
  assign validSink_15_bits_csrInterface_vStart = shifterReg_15_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_15_0_bits_csrInterface_vlmul;
  assign validSink_15_bits_csrInterface_vlmul = shifterReg_15_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_15_0_bits_csrInterface_vSew;
  assign validSink_15_bits_csrInterface_vSew = shifterReg_15_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_15_0_bits_csrInterface_vxrm;
  assign validSink_15_bits_csrInterface_vxrm = shifterReg_15_0_bits_csrInterface_vxrm;
  reg          shifterReg_15_0_bits_csrInterface_vta;
  assign validSink_15_bits_csrInterface_vta = shifterReg_15_0_bits_csrInterface_vta;
  reg          shifterReg_15_0_bits_csrInterface_vma;
  assign validSink_15_bits_csrInterface_vma = shifterReg_15_0_bits_csrInterface_vma;
  wire         shifterValid_15 = shifterReg_15_0_valid | validSource_15_valid;
  wire [1:0]   allLaneReady_lo_lo_lo = {laneRequestSourceWire_1_ready, laneRequestSourceWire_0_ready};
  wire [1:0]   allLaneReady_lo_lo_hi = {laneRequestSourceWire_3_ready, laneRequestSourceWire_2_ready};
  wire [3:0]   allLaneReady_lo_lo = {allLaneReady_lo_lo_hi, allLaneReady_lo_lo_lo};
  wire [1:0]   allLaneReady_lo_hi_lo = {laneRequestSourceWire_5_ready, laneRequestSourceWire_4_ready};
  wire [1:0]   allLaneReady_lo_hi_hi = {laneRequestSourceWire_7_ready, laneRequestSourceWire_6_ready};
  wire [3:0]   allLaneReady_lo_hi = {allLaneReady_lo_hi_hi, allLaneReady_lo_hi_lo};
  wire [7:0]   allLaneReady_lo = {allLaneReady_lo_hi, allLaneReady_lo_lo};
  wire [1:0]   allLaneReady_hi_lo_lo = {laneRequestSourceWire_9_ready, laneRequestSourceWire_8_ready};
  wire [1:0]   allLaneReady_hi_lo_hi = {laneRequestSourceWire_11_ready, laneRequestSourceWire_10_ready};
  wire [3:0]   allLaneReady_hi_lo = {allLaneReady_hi_lo_hi, allLaneReady_hi_lo_lo};
  wire [1:0]   allLaneReady_hi_hi_lo = {laneRequestSourceWire_13_ready, laneRequestSourceWire_12_ready};
  wire [1:0]   allLaneReady_hi_hi_hi = {laneRequestSourceWire_15_ready, laneRequestSourceWire_14_ready};
  wire [3:0]   allLaneReady_hi_hi = {allLaneReady_hi_hi_hi, allLaneReady_hi_hi_lo};
  wire [7:0]   allLaneReady_hi = {allLaneReady_hi_hi, allLaneReady_hi_lo};
  wire         allLaneReady = &{allLaneReady_hi, allLaneReady_lo};
  wire         completeIndexInstruction = (|(8'h1 << _GEN_2 & _lsu_lastReport)) & ~slots_3_state_idle;
  wire [1:0]   _GEN_3 = {slots_1_state_idle, slots_0_state_idle};
  wire [1:0]   freeOR_lo;
  assign freeOR_lo = _GEN_3;
  wire [1:0]   free_lo;
  assign free_lo = _GEN_3;
  wire [1:0]   _GEN_4 = {slots_3_state_idle, slots_2_state_idle};
  wire [1:0]   freeOR_hi;
  assign freeOR_hi = _GEN_4;
  wire [1:0]   free_hi;
  assign free_hi = _GEN_4;
  wire         freeOR = |{freeOR_hi, freeOR_lo};
  wire         slotReady = specialInstruction ? slots_3_state_idle : freeOR;
  wire         olderCheck_notSameLSB = slots_0_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_1 = slots_1_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_2 = slots_2_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_3 = slots_3_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck =
    (slots_0_state_idle | (slots_0_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_0_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB)
    & (slots_1_state_idle | (slots_1_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_1_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_1)
    & (slots_2_state_idle | (slots_2_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_2_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_2)
    & (slots_3_state_idle | (slots_3_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_3_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_3);
  assign source1Select = requestReg_bits_decodeResult_gather ? _maskUnit_gatherData_bits : requestReg_bits_decodeResult_itype ? immSignExtend : source1Extend;
  assign laneRequestSourceWire_0_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_1_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_2_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_3_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_4_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_5_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_6_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_7_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_8_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_9_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_10_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_11_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_12_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_13_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_14_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_15_bits_readFromScalar = source1Select;
  wire         extendDataEEW = requestReg_bits_issue_vtype[3] - requestReg_bits_decodeResult_topUop[1];
  assign laneRequestSourceWire_0_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_1_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_2_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_3_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_4_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_5_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_6_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_7_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_8_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_9_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_10_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_11_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_12_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_13_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_14_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_15_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  wire [2:0]   vSewSelect =
    isLoadStoreType
      ? {1'h0, requestRegDequeue_bits_instruction[13:12]}
      : requestReg_bits_decodeResult_nr | requestReg_bits_decodeResult_maskLogic ? 3'h2 : requestReg_bits_decodeResult_gather16 ? 3'h1 : requestReg_bits_decodeResult_extend ? {2'h0, extendDataEEW} : requestReg_bits_issue_vtype[5:3];
  wire [31:0]  evlForLane = requestReg_bits_decodeResult_nr ? {22'h0, {1'h0, requestRegDequeue_bits_instruction[17:15]} + 4'h1, 6'h0} : requestReg_bits_issue_vl;
  wire [1:0]   vSewForLsu = lsWholeReg ? 2'h2 : requestRegDequeue_bits_instruction[13:12];
  wire [31:0]  evlForLsu = lsWholeReg ? {22'h0, {1'h0, requestRegDequeue_bits_instruction[31:29]} + 4'h1, 6'h0} : requestReg_bits_issue_vl;
  assign laneRequestSourceWire_0_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_1_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_2_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_3_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_4_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_5_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_6_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_7_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_8_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_9_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_10_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_11_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_12_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_13_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_14_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_15_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_0_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_1_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_2_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_3_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_4_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_5_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_6_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_7_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_8_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_9_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_10_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_11_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_12_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_13_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_14_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_15_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_0_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_0_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_0_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_1_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_2_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_3_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_4_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_5_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_6_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_7_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_8_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_9_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_10_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_11_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_12_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_13_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_14_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_15_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_0_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_1_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_2_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_3_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_4_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_5_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_6_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_7_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_8_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_9_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_10_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_11_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_12_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_13_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_14_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_15_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_1_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_1_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_2_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_2_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_3_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_3_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_4_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_4_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_5_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_5_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_6_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_6_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_7_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_7_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_8_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_8_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_9_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_9_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_10_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_10_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_11_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_11_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_12_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_12_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_13_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_13_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_14_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_14_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_15_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_15_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSinkWire_0_ready = ~laneRequestSinkWire_0_bits_issueInst | _laneVec_0_laneRequest_ready;
  wire         sinkVec_tokenCheck;
  wire [4:0]   sinkVec_validSource_bits_vs = x13_0_bits_vs;
  wire [1:0]   sinkVec_validSource_bits_offset = x13_0_bits_offset;
  wire [2:0]   sinkVec_validSource_bits_instructionIndex = x13_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_1;
  wire [4:0]   sinkVec_validSource_1_bits_vs = x13_1_bits_vs;
  wire [1:0]   sinkVec_validSource_1_bits_offset = x13_1_bits_offset;
  wire [2:0]   sinkVec_validSource_1_bits_instructionIndex = x13_1_bits_instructionIndex;
  wire         sinkVec_0_ready;
  wire         sinkVec_queue_deq_ready = sinkVec_sinkWire_ready;
  wire         sinkVec_queue_deq_valid;
  wire [4:0]   sinkVec_queue_deq_bits_vs;
  wire         sinkVec_0_valid = sinkVec_sinkWire_valid;
  wire [1:0]   sinkVec_queue_deq_bits_readSource;
  wire [4:0]   sinkVec_0_bits_vs = sinkVec_sinkWire_bits_vs;
  wire [1:0]   sinkVec_queue_deq_bits_offset;
  wire [1:0]   sinkVec_0_bits_readSource = sinkVec_sinkWire_bits_readSource;
  wire [2:0]   sinkVec_queue_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_0_bits_offset = sinkVec_sinkWire_bits_offset;
  wire [2:0]   sinkVec_0_bits_instructionIndex = sinkVec_sinkWire_bits_instructionIndex;
  wire         sinkVec_validSink_valid;
  wire [4:0]   sinkVec_validSink_bits_vs;
  wire [1:0]   sinkVec_validSink_bits_readSource;
  wire [1:0]   sinkVec_validSink_bits_offset;
  wire [2:0]   sinkVec_validSink_bits_instructionIndex;
  assign sinkVec_sinkWire_valid = sinkVec_queue_deq_valid;
  assign sinkVec_sinkWire_bits_vs = sinkVec_queue_deq_bits_vs;
  assign sinkVec_sinkWire_bits_readSource = sinkVec_queue_deq_bits_readSource;
  assign sinkVec_sinkWire_bits_offset = sinkVec_queue_deq_bits_offset;
  assign sinkVec_sinkWire_bits_instructionIndex = sinkVec_queue_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_enq_bits_offset;
  wire [2:0]   sinkVec_queue_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo = {sinkVec_queue_enq_bits_offset, sinkVec_queue_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_enq_bits_vs;
  wire [1:0]   sinkVec_queue_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi = {sinkVec_queue_enq_bits_vs, sinkVec_queue_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn = {sinkVec_queue_dataIn_hi, sinkVec_queue_dataIn_lo};
  wire [2:0]   sinkVec_queue_dataOut_instructionIndex = _sinkVec_queue_fifo_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_offset = _sinkVec_queue_fifo_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_readSource = _sinkVec_queue_fifo_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_vs = _sinkVec_queue_fifo_data_out[11:7];
  wire         sinkVec_queue_enq_ready = ~_sinkVec_queue_fifo_full;
  wire         sinkVec_queue_enq_valid;
  assign sinkVec_queue_deq_valid = ~_sinkVec_queue_fifo_empty | sinkVec_queue_enq_valid;
  assign sinkVec_queue_deq_bits_vs = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_vs : sinkVec_queue_dataOut_vs;
  assign sinkVec_queue_deq_bits_readSource = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_readSource : sinkVec_queue_dataOut_readSource;
  assign sinkVec_queue_deq_bits_offset = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_offset : sinkVec_queue_dataOut_offset;
  assign sinkVec_queue_deq_bits_instructionIndex = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_instructionIndex : sinkVec_queue_dataOut_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v;
  wire         sinkVec_releasePipe_pipe_out_valid = sinkVec_releasePipe_pipe_v;
  wire         x13_0_ready;
  wire         x13_0_valid;
  wire         sinkVec_validSource_valid = x13_0_ready & x13_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter;
  wire [2:0]   sinkVec_tokenCheck_counterChange = sinkVec_validSource_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck = ~(sinkVec_tokenCheck_counter[2]);
  assign x13_0_ready = sinkVec_tokenCheck;
  assign sinkVec_queue_enq_valid = sinkVec_validSink_valid;
  assign sinkVec_queue_enq_bits_vs = sinkVec_validSink_bits_vs;
  assign sinkVec_queue_enq_bits_readSource = sinkVec_validSink_bits_readSource;
  assign sinkVec_queue_enq_bits_offset = sinkVec_validSink_bits_offset;
  assign sinkVec_queue_enq_bits_instructionIndex = sinkVec_validSink_bits_instructionIndex;
  reg          sinkVec_shifterReg_0_valid;
  assign sinkVec_validSink_valid = sinkVec_shifterReg_0_valid;
  reg  [4:0]   sinkVec_shifterReg_0_bits_vs;
  assign sinkVec_validSink_bits_vs = sinkVec_shifterReg_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_0_bits_readSource;
  assign sinkVec_validSink_bits_readSource = sinkVec_shifterReg_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_0_bits_offset;
  assign sinkVec_validSink_bits_offset = sinkVec_shifterReg_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_0_bits_instructionIndex;
  assign sinkVec_validSink_bits_instructionIndex = sinkVec_shifterReg_0_bits_instructionIndex;
  wire         sinkVec_shifterValid = sinkVec_shifterReg_0_valid | sinkVec_validSource_valid;
  wire         sinkVec_1_ready;
  wire         sinkVec_queue_1_deq_ready = sinkVec_sinkWire_1_ready;
  wire         sinkVec_queue_1_deq_valid;
  wire [4:0]   sinkVec_queue_1_deq_bits_vs;
  wire         sinkVec_1_valid = sinkVec_sinkWire_1_valid;
  wire [1:0]   sinkVec_queue_1_deq_bits_readSource;
  wire [4:0]   sinkVec_1_bits_vs = sinkVec_sinkWire_1_bits_vs;
  wire [1:0]   sinkVec_queue_1_deq_bits_offset;
  wire [1:0]   sinkVec_1_bits_readSource = sinkVec_sinkWire_1_bits_readSource;
  wire [2:0]   sinkVec_queue_1_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_1_bits_offset = sinkVec_sinkWire_1_bits_offset;
  wire [2:0]   sinkVec_1_bits_instructionIndex = sinkVec_sinkWire_1_bits_instructionIndex;
  wire         sinkVec_validSink_1_valid;
  wire [4:0]   sinkVec_validSink_1_bits_vs;
  wire [1:0]   sinkVec_validSink_1_bits_readSource;
  wire [1:0]   sinkVec_validSink_1_bits_offset;
  wire [2:0]   sinkVec_validSink_1_bits_instructionIndex;
  assign sinkVec_sinkWire_1_valid = sinkVec_queue_1_deq_valid;
  assign sinkVec_sinkWire_1_bits_vs = sinkVec_queue_1_deq_bits_vs;
  assign sinkVec_sinkWire_1_bits_readSource = sinkVec_queue_1_deq_bits_readSource;
  assign sinkVec_sinkWire_1_bits_offset = sinkVec_queue_1_deq_bits_offset;
  assign sinkVec_sinkWire_1_bits_instructionIndex = sinkVec_queue_1_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_1_enq_bits_offset;
  wire [2:0]   sinkVec_queue_1_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_1 = {sinkVec_queue_1_enq_bits_offset, sinkVec_queue_1_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_1_enq_bits_vs;
  wire [1:0]   sinkVec_queue_1_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_1 = {sinkVec_queue_1_enq_bits_vs, sinkVec_queue_1_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_1 = {sinkVec_queue_dataIn_hi_1, sinkVec_queue_dataIn_lo_1};
  wire [2:0]   sinkVec_queue_dataOut_1_instructionIndex = _sinkVec_queue_fifo_1_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_1_offset = _sinkVec_queue_fifo_1_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_1_readSource = _sinkVec_queue_fifo_1_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_1_vs = _sinkVec_queue_fifo_1_data_out[11:7];
  wire         sinkVec_queue_1_enq_ready = ~_sinkVec_queue_fifo_1_full;
  wire         sinkVec_queue_1_enq_valid;
  assign sinkVec_queue_1_deq_valid = ~_sinkVec_queue_fifo_1_empty | sinkVec_queue_1_enq_valid;
  assign sinkVec_queue_1_deq_bits_vs = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_vs : sinkVec_queue_dataOut_1_vs;
  assign sinkVec_queue_1_deq_bits_readSource = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_readSource : sinkVec_queue_dataOut_1_readSource;
  assign sinkVec_queue_1_deq_bits_offset = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_offset : sinkVec_queue_dataOut_1_offset;
  assign sinkVec_queue_1_deq_bits_instructionIndex = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_instructionIndex : sinkVec_queue_dataOut_1_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_1;
  wire         sinkVec_releasePipe_pipe_out_1_valid = sinkVec_releasePipe_pipe_v_1;
  wire         x13_1_ready;
  wire         x13_1_valid;
  wire         sinkVec_validSource_1_valid = x13_1_ready & x13_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_1;
  wire [2:0]   sinkVec_tokenCheck_counterChange_1 = sinkVec_validSource_1_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_1 = ~(sinkVec_tokenCheck_counter_1[2]);
  assign x13_1_ready = sinkVec_tokenCheck_1;
  assign sinkVec_queue_1_enq_valid = sinkVec_validSink_1_valid;
  assign sinkVec_queue_1_enq_bits_vs = sinkVec_validSink_1_bits_vs;
  assign sinkVec_queue_1_enq_bits_readSource = sinkVec_validSink_1_bits_readSource;
  assign sinkVec_queue_1_enq_bits_offset = sinkVec_validSink_1_bits_offset;
  assign sinkVec_queue_1_enq_bits_instructionIndex = sinkVec_validSink_1_bits_instructionIndex;
  reg          sinkVec_shifterReg_1_0_valid;
  assign sinkVec_validSink_1_valid = sinkVec_shifterReg_1_0_valid;
  reg  [4:0]   sinkVec_shifterReg_1_0_bits_vs;
  assign sinkVec_validSink_1_bits_vs = sinkVec_shifterReg_1_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_1_0_bits_readSource;
  assign sinkVec_validSink_1_bits_readSource = sinkVec_shifterReg_1_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_1_0_bits_offset;
  assign sinkVec_validSink_1_bits_offset = sinkVec_shifterReg_1_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_1_0_bits_instructionIndex;
  assign sinkVec_validSink_1_bits_instructionIndex = sinkVec_shifterReg_1_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_1 = sinkVec_shifterReg_1_0_valid | sinkVec_validSource_1_valid;
  assign sinkVec_sinkWire_ready = sinkVec_0_ready;
  assign sinkVec_sinkWire_1_ready = sinkVec_1_ready;
  reg          maskUnitFirst;
  wire         tryToRead = sinkVec_0_valid | sinkVec_1_valid;
  wire         sinkWire_valid = maskUnitFirst ? sinkVec_0_valid : sinkVec_1_valid;
  wire [4:0]   sinkWire_bits_vs = maskUnitFirst ? sinkVec_0_bits_vs : sinkVec_1_bits_vs;
  wire [1:0]   sinkWire_bits_readSource = maskUnitFirst ? sinkVec_0_bits_readSource : sinkVec_1_bits_readSource;
  wire [1:0]   sinkWire_bits_offset = maskUnitFirst ? sinkVec_0_bits_offset : sinkVec_1_bits_offset;
  wire [2:0]   sinkWire_bits_instructionIndex = maskUnitFirst ? sinkVec_0_bits_instructionIndex : sinkVec_1_bits_instructionIndex;
  wire         sinkWire_ready;
  assign sinkVec_1_ready = sinkWire_ready & ~maskUnitFirst;
  assign sinkVec_0_ready = sinkWire_ready & maskUnitFirst;
  reg          accessDataValid_pipe_v;
  reg          accessDataValid_pipe_pipe_v;
  wire         accessDataValid_pipe_pipe_out_valid = accessDataValid_pipe_pipe_v;
  wire         accessDataSource_valid = accessDataValid_pipe_pipe_out_valid;
  reg          shifterReg_16_0_valid;
  reg  [31:0]  shifterReg_16_0_bits;
  wire         shifterValid_16 = shifterReg_16_0_valid | accessDataSource_valid;
  reg          accessDataValid_pipe_v_1;
  reg          accessDataValid_pipe_pipe_v_1;
  wire         accessDataValid_pipe_pipe_out_1_valid = accessDataValid_pipe_pipe_v_1;
  wire         accessDataSource_1_valid = accessDataValid_pipe_pipe_out_1_valid;
  reg          shifterReg_17_0_valid;
  reg  [31:0]  shifterReg_17_0_bits;
  wire         shifterValid_17 = shifterReg_17_0_valid | accessDataSource_1_valid;
  wire         sinkVec_tokenCheck_2;
  wire [4:0]   sinkVec_validSource_2_bits_vd = x22_0_bits_vd;
  wire [1:0]   sinkVec_validSource_2_bits_offset = x22_0_bits_offset;
  wire [3:0]   sinkVec_validSource_2_bits_mask = x22_0_bits_mask;
  wire [31:0]  sinkVec_validSource_2_bits_data = x22_0_bits_data;
  wire [2:0]   sinkVec_validSource_2_bits_instructionIndex = x22_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_3;
  wire [4:0]   sinkVec_validSource_3_bits_vd = x22_1_bits_vd;
  wire [1:0]   sinkVec_validSource_3_bits_offset = x22_1_bits_offset;
  wire [3:0]   sinkVec_validSource_3_bits_mask = x22_1_bits_mask;
  wire [31:0]  sinkVec_validSource_3_bits_data = x22_1_bits_data;
  wire         sinkVec_validSource_3_bits_last = x22_1_bits_last;
  wire [2:0]   sinkVec_validSource_3_bits_instructionIndex = x22_1_bits_instructionIndex;
  wire         sinkVec_1_0_ready;
  wire         sinkVec_queue_2_deq_ready = sinkVec_sinkWire_2_ready;
  wire         sinkVec_queue_2_deq_valid;
  wire [4:0]   sinkVec_queue_2_deq_bits_vd;
  wire         sinkVec_1_0_valid = sinkVec_sinkWire_2_valid;
  wire [1:0]   sinkVec_queue_2_deq_bits_offset;
  wire [4:0]   sinkVec_1_0_bits_vd = sinkVec_sinkWire_2_bits_vd;
  wire [3:0]   sinkVec_queue_2_deq_bits_mask;
  wire [1:0]   sinkVec_1_0_bits_offset = sinkVec_sinkWire_2_bits_offset;
  wire [31:0]  sinkVec_queue_2_deq_bits_data;
  wire [3:0]   sinkVec_1_0_bits_mask = sinkVec_sinkWire_2_bits_mask;
  wire         sinkVec_queue_2_deq_bits_last;
  wire [31:0]  sinkVec_1_0_bits_data = sinkVec_sinkWire_2_bits_data;
  wire [2:0]   sinkVec_queue_2_deq_bits_instructionIndex;
  wire         sinkVec_1_0_bits_last = sinkVec_sinkWire_2_bits_last;
  wire [2:0]   sinkVec_1_0_bits_instructionIndex = sinkVec_sinkWire_2_bits_instructionIndex;
  wire         sinkVec_validSink_2_valid;
  wire [4:0]   sinkVec_validSink_2_bits_vd;
  wire [1:0]   sinkVec_validSink_2_bits_offset;
  wire [3:0]   sinkVec_validSink_2_bits_mask;
  wire [31:0]  sinkVec_validSink_2_bits_data;
  wire [2:0]   sinkVec_validSink_2_bits_instructionIndex;
  assign sinkVec_sinkWire_2_valid = sinkVec_queue_2_deq_valid;
  assign sinkVec_sinkWire_2_bits_vd = sinkVec_queue_2_deq_bits_vd;
  assign sinkVec_sinkWire_2_bits_offset = sinkVec_queue_2_deq_bits_offset;
  assign sinkVec_sinkWire_2_bits_mask = sinkVec_queue_2_deq_bits_mask;
  assign sinkVec_sinkWire_2_bits_data = sinkVec_queue_2_deq_bits_data;
  assign sinkVec_sinkWire_2_bits_last = sinkVec_queue_2_deq_bits_last;
  assign sinkVec_sinkWire_2_bits_instructionIndex = sinkVec_queue_2_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_2_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi = {sinkVec_queue_2_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_2_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_2 = {sinkVec_queue_dataIn_lo_hi, sinkVec_queue_2_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_2_enq_bits_vd;
  wire [1:0]   sinkVec_queue_2_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi = {sinkVec_queue_2_enq_bits_vd, sinkVec_queue_2_enq_bits_offset};
  wire [3:0]   sinkVec_queue_2_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_2 = {sinkVec_queue_dataIn_hi_hi, sinkVec_queue_2_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_2 = {sinkVec_queue_dataIn_hi_2, sinkVec_queue_dataIn_lo_2};
  wire [2:0]   sinkVec_queue_dataOut_2_instructionIndex = _sinkVec_queue_fifo_2_data_out[2:0];
  wire         sinkVec_queue_dataOut_2_last = _sinkVec_queue_fifo_2_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_2_data = _sinkVec_queue_fifo_2_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_2_mask = _sinkVec_queue_fifo_2_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_2_offset = _sinkVec_queue_fifo_2_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_2_vd = _sinkVec_queue_fifo_2_data_out[46:42];
  wire         sinkVec_queue_2_enq_ready = ~_sinkVec_queue_fifo_2_full;
  wire         sinkVec_queue_2_enq_valid;
  assign sinkVec_queue_2_deq_valid = ~_sinkVec_queue_fifo_2_empty | sinkVec_queue_2_enq_valid;
  assign sinkVec_queue_2_deq_bits_vd = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_vd : sinkVec_queue_dataOut_2_vd;
  assign sinkVec_queue_2_deq_bits_offset = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_offset : sinkVec_queue_dataOut_2_offset;
  assign sinkVec_queue_2_deq_bits_mask = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_mask : sinkVec_queue_dataOut_2_mask;
  assign sinkVec_queue_2_deq_bits_data = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_data : sinkVec_queue_dataOut_2_data;
  assign sinkVec_queue_2_deq_bits_last = ~_sinkVec_queue_fifo_2_empty & sinkVec_queue_dataOut_2_last;
  assign sinkVec_queue_2_deq_bits_instructionIndex = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_instructionIndex : sinkVec_queue_dataOut_2_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_2;
  wire         sinkVec_releasePipe_pipe_out_2_valid = sinkVec_releasePipe_pipe_v_2;
  wire         x22_0_ready;
  wire         x22_0_valid;
  wire         sinkVec_validSource_2_valid = x22_0_ready & x22_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_2;
  wire [2:0]   sinkVec_tokenCheck_counterChange_2 = sinkVec_validSource_2_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_2 = ~(sinkVec_tokenCheck_counter_2[2]);
  assign x22_0_ready = sinkVec_tokenCheck_2;
  assign sinkVec_queue_2_enq_valid = sinkVec_validSink_2_valid;
  assign sinkVec_queue_2_enq_bits_vd = sinkVec_validSink_2_bits_vd;
  assign sinkVec_queue_2_enq_bits_offset = sinkVec_validSink_2_bits_offset;
  assign sinkVec_queue_2_enq_bits_mask = sinkVec_validSink_2_bits_mask;
  assign sinkVec_queue_2_enq_bits_data = sinkVec_validSink_2_bits_data;
  assign sinkVec_queue_2_enq_bits_instructionIndex = sinkVec_validSink_2_bits_instructionIndex;
  reg          sinkVec_shifterReg_2_0_valid;
  assign sinkVec_validSink_2_valid = sinkVec_shifterReg_2_0_valid;
  reg  [4:0]   sinkVec_shifterReg_2_0_bits_vd;
  assign sinkVec_validSink_2_bits_vd = sinkVec_shifterReg_2_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_2_0_bits_offset;
  assign sinkVec_validSink_2_bits_offset = sinkVec_shifterReg_2_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_2_0_bits_mask;
  assign sinkVec_validSink_2_bits_mask = sinkVec_shifterReg_2_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_2_0_bits_data;
  assign sinkVec_validSink_2_bits_data = sinkVec_shifterReg_2_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_2_0_bits_instructionIndex;
  assign sinkVec_validSink_2_bits_instructionIndex = sinkVec_shifterReg_2_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_2 = sinkVec_shifterReg_2_0_valid | sinkVec_validSource_2_valid;
  wire         sinkVec_1_1_ready;
  wire         sinkVec_queue_3_deq_ready = sinkVec_sinkWire_3_ready;
  wire         sinkVec_queue_3_deq_valid;
  wire [4:0]   sinkVec_queue_3_deq_bits_vd;
  wire         sinkVec_1_1_valid = sinkVec_sinkWire_3_valid;
  wire [1:0]   sinkVec_queue_3_deq_bits_offset;
  wire [4:0]   sinkVec_1_1_bits_vd = sinkVec_sinkWire_3_bits_vd;
  wire [3:0]   sinkVec_queue_3_deq_bits_mask;
  wire [1:0]   sinkVec_1_1_bits_offset = sinkVec_sinkWire_3_bits_offset;
  wire [31:0]  sinkVec_queue_3_deq_bits_data;
  wire [3:0]   sinkVec_1_1_bits_mask = sinkVec_sinkWire_3_bits_mask;
  wire         sinkVec_queue_3_deq_bits_last;
  wire [31:0]  sinkVec_1_1_bits_data = sinkVec_sinkWire_3_bits_data;
  wire [2:0]   sinkVec_queue_3_deq_bits_instructionIndex;
  wire         sinkVec_1_1_bits_last = sinkVec_sinkWire_3_bits_last;
  wire [2:0]   sinkVec_1_1_bits_instructionIndex = sinkVec_sinkWire_3_bits_instructionIndex;
  wire         sinkVec_validSink_3_valid;
  wire [4:0]   sinkVec_validSink_3_bits_vd;
  wire [1:0]   sinkVec_validSink_3_bits_offset;
  wire [3:0]   sinkVec_validSink_3_bits_mask;
  wire [31:0]  sinkVec_validSink_3_bits_data;
  wire         sinkVec_validSink_3_bits_last;
  wire [2:0]   sinkVec_validSink_3_bits_instructionIndex;
  assign sinkVec_sinkWire_3_valid = sinkVec_queue_3_deq_valid;
  assign sinkVec_sinkWire_3_bits_vd = sinkVec_queue_3_deq_bits_vd;
  assign sinkVec_sinkWire_3_bits_offset = sinkVec_queue_3_deq_bits_offset;
  assign sinkVec_sinkWire_3_bits_mask = sinkVec_queue_3_deq_bits_mask;
  assign sinkVec_sinkWire_3_bits_data = sinkVec_queue_3_deq_bits_data;
  assign sinkVec_sinkWire_3_bits_last = sinkVec_queue_3_deq_bits_last;
  assign sinkVec_sinkWire_3_bits_instructionIndex = sinkVec_queue_3_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_3_enq_bits_data;
  wire         sinkVec_queue_3_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_1 = {sinkVec_queue_3_enq_bits_data, sinkVec_queue_3_enq_bits_last};
  wire [2:0]   sinkVec_queue_3_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_3 = {sinkVec_queue_dataIn_lo_hi_1, sinkVec_queue_3_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_3_enq_bits_vd;
  wire [1:0]   sinkVec_queue_3_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_1 = {sinkVec_queue_3_enq_bits_vd, sinkVec_queue_3_enq_bits_offset};
  wire [3:0]   sinkVec_queue_3_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_3 = {sinkVec_queue_dataIn_hi_hi_1, sinkVec_queue_3_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_3 = {sinkVec_queue_dataIn_hi_3, sinkVec_queue_dataIn_lo_3};
  wire [2:0]   sinkVec_queue_dataOut_3_instructionIndex = _sinkVec_queue_fifo_3_data_out[2:0];
  wire         sinkVec_queue_dataOut_3_last = _sinkVec_queue_fifo_3_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_3_data = _sinkVec_queue_fifo_3_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_3_mask = _sinkVec_queue_fifo_3_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_3_offset = _sinkVec_queue_fifo_3_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_3_vd = _sinkVec_queue_fifo_3_data_out[46:42];
  wire         sinkVec_queue_3_enq_ready = ~_sinkVec_queue_fifo_3_full;
  wire         sinkVec_queue_3_enq_valid;
  assign sinkVec_queue_3_deq_valid = ~_sinkVec_queue_fifo_3_empty | sinkVec_queue_3_enq_valid;
  assign sinkVec_queue_3_deq_bits_vd = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_vd : sinkVec_queue_dataOut_3_vd;
  assign sinkVec_queue_3_deq_bits_offset = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_offset : sinkVec_queue_dataOut_3_offset;
  assign sinkVec_queue_3_deq_bits_mask = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_mask : sinkVec_queue_dataOut_3_mask;
  assign sinkVec_queue_3_deq_bits_data = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_data : sinkVec_queue_dataOut_3_data;
  assign sinkVec_queue_3_deq_bits_last = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_last : sinkVec_queue_dataOut_3_last;
  assign sinkVec_queue_3_deq_bits_instructionIndex = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_instructionIndex : sinkVec_queue_dataOut_3_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_3;
  wire         sinkVec_releasePipe_pipe_out_3_valid = sinkVec_releasePipe_pipe_v_3;
  wire         x22_1_ready;
  wire         x22_1_valid;
  wire         sinkVec_validSource_3_valid = x22_1_ready & x22_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_3;
  wire [2:0]   sinkVec_tokenCheck_counterChange_3 = sinkVec_validSource_3_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_3 = ~(sinkVec_tokenCheck_counter_3[2]);
  assign x22_1_ready = sinkVec_tokenCheck_3;
  assign sinkVec_queue_3_enq_valid = sinkVec_validSink_3_valid;
  assign sinkVec_queue_3_enq_bits_vd = sinkVec_validSink_3_bits_vd;
  assign sinkVec_queue_3_enq_bits_offset = sinkVec_validSink_3_bits_offset;
  assign sinkVec_queue_3_enq_bits_mask = sinkVec_validSink_3_bits_mask;
  assign sinkVec_queue_3_enq_bits_data = sinkVec_validSink_3_bits_data;
  assign sinkVec_queue_3_enq_bits_last = sinkVec_validSink_3_bits_last;
  assign sinkVec_queue_3_enq_bits_instructionIndex = sinkVec_validSink_3_bits_instructionIndex;
  reg          sinkVec_shifterReg_3_0_valid;
  assign sinkVec_validSink_3_valid = sinkVec_shifterReg_3_0_valid;
  reg  [4:0]   sinkVec_shifterReg_3_0_bits_vd;
  assign sinkVec_validSink_3_bits_vd = sinkVec_shifterReg_3_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_3_0_bits_offset;
  assign sinkVec_validSink_3_bits_offset = sinkVec_shifterReg_3_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_3_0_bits_mask;
  assign sinkVec_validSink_3_bits_mask = sinkVec_shifterReg_3_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_3_0_bits_data;
  assign sinkVec_validSink_3_bits_data = sinkVec_shifterReg_3_0_bits_data;
  reg          sinkVec_shifterReg_3_0_bits_last;
  assign sinkVec_validSink_3_bits_last = sinkVec_shifterReg_3_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_3_0_bits_instructionIndex;
  assign sinkVec_validSink_3_bits_instructionIndex = sinkVec_shifterReg_3_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_3 = sinkVec_shifterReg_3_0_valid | sinkVec_validSource_3_valid;
  assign sinkVec_sinkWire_2_ready = sinkVec_1_0_ready;
  assign sinkVec_sinkWire_3_ready = sinkVec_1_1_ready;
  reg          maskUnitFirst_1;
  wire         tryToRead_1 = sinkVec_1_0_valid | sinkVec_1_1_valid;
  wire         sinkWire_1_valid = maskUnitFirst_1 ? sinkVec_1_0_valid : sinkVec_1_1_valid;
  wire [4:0]   sinkWire_1_bits_vd = maskUnitFirst_1 ? sinkVec_1_0_bits_vd : sinkVec_1_1_bits_vd;
  wire [1:0]   sinkWire_1_bits_offset = maskUnitFirst_1 ? sinkVec_1_0_bits_offset : sinkVec_1_1_bits_offset;
  wire [3:0]   sinkWire_1_bits_mask = maskUnitFirst_1 ? sinkVec_1_0_bits_mask : sinkVec_1_1_bits_mask;
  wire [31:0]  sinkWire_1_bits_data = maskUnitFirst_1 ? sinkVec_1_0_bits_data : sinkVec_1_1_bits_data;
  wire         sinkWire_1_bits_last = maskUnitFirst_1 ? sinkVec_1_0_bits_last : sinkVec_1_1_bits_last;
  wire [2:0]   sinkWire_1_bits_instructionIndex = maskUnitFirst_1 ? sinkVec_1_0_bits_instructionIndex : sinkVec_1_1_bits_instructionIndex;
  wire         sinkWire_1_ready;
  assign sinkVec_1_1_ready = sinkWire_1_ready & ~maskUnitFirst_1;
  assign sinkVec_1_0_ready = sinkWire_1_ready & maskUnitFirst_1;
  reg          view__writeRelease_0_pipe_v;
  wire         view__writeRelease_0_pipe_out_valid = view__writeRelease_0_pipe_v;
  reg          pipe_v;
  wire         pipe_out_valid = pipe_v;
  wire         _probeWire_writeQueueEnqVec_0_valid_T = x22_0_ready & _maskUnit_exeResp_0_valid;
  reg          instructionFinishedPipe_pipe_v;
  wire         instructionFinishedPipe_pipe_out_valid = instructionFinishedPipe_pipe_v;
  reg  [7:0]   instructionFinishedPipe_pipe_b;
  wire [7:0]   instructionFinishedPipe_pipe_out_bits = instructionFinishedPipe_pipe_b;
  wire         instructionFinished_0_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_bits);
  assign vxsatReportVec_0 = _laneVec_0_vxsatReport[3:0];
  reg          pipe_v_1;
  reg  [31:0]  pipe_b_1;
  reg          pipe_pipe_v;
  wire         pipe_pipe_out_valid = pipe_pipe_v;
  reg  [31:0]  pipe_pipe_b;
  wire [31:0]  pipe_pipe_out_bits = pipe_pipe_b;
  reg          view__laneMaskSelect_0_pipe_v;
  reg  [5:0]   view__laneMaskSelect_0_pipe_b;
  reg          view__laneMaskSelect_0_pipe_pipe_v;
  wire         view__laneMaskSelect_0_pipe_pipe_out_valid = view__laneMaskSelect_0_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_0_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_0_pipe_pipe_out_bits = view__laneMaskSelect_0_pipe_pipe_b;
  reg          view__laneMaskSewSelect_0_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_0_pipe_b;
  reg          view__laneMaskSewSelect_0_pipe_pipe_v;
  wire         view__laneMaskSewSelect_0_pipe_pipe_out_valid = view__laneMaskSewSelect_0_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_0_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_0_pipe_pipe_out_bits = view__laneMaskSewSelect_0_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v;
  wire         lsuLastPipe_pipe_out_valid = lsuLastPipe_pipe_v;
  reg  [7:0]   lsuLastPipe_pipe_b;
  wire [7:0]   lsuLastPipe_pipe_out_bits = lsuLastPipe_pipe_b;
  reg          maskLastPipe_pipe_v;
  wire         maskLastPipe_pipe_out_valid = maskLastPipe_pipe_v;
  reg  [7:0]   maskLastPipe_pipe_b;
  wire [7:0]   maskLastPipe_pipe_out_bits = maskLastPipe_pipe_b;
  wire [5:0]   writeCounter = requestReg_bits_writeByte[11:6] + {5'h0, |(requestReg_bits_writeByte[5:0])};
  reg          pipe_v_2;
  wire         pipe_out_1_valid = pipe_v_2;
  reg  [5:0]   pipe_b_2;
  wire [5:0]   pipe_out_1_bits = pipe_b_2;
  assign laneRequestSinkWire_1_ready = ~laneRequestSinkWire_1_bits_issueInst | _laneVec_1_laneRequest_ready;
  wire         sinkVec_tokenCheck_4;
  wire [4:0]   sinkVec_validSource_4_bits_vs = x13_1_0_bits_vs;
  wire [1:0]   sinkVec_validSource_4_bits_offset = x13_1_0_bits_offset;
  wire [2:0]   sinkVec_validSource_4_bits_instructionIndex = x13_1_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_5;
  wire [4:0]   sinkVec_validSource_5_bits_vs = x13_1_1_bits_vs;
  wire [1:0]   sinkVec_validSource_5_bits_offset = x13_1_1_bits_offset;
  wire [2:0]   sinkVec_validSource_5_bits_instructionIndex = x13_1_1_bits_instructionIndex;
  wire         sinkVec_2_0_ready;
  wire         sinkVec_queue_4_deq_ready = sinkVec_sinkWire_4_ready;
  wire         sinkVec_queue_4_deq_valid;
  wire [4:0]   sinkVec_queue_4_deq_bits_vs;
  wire         sinkVec_2_0_valid = sinkVec_sinkWire_4_valid;
  wire [1:0]   sinkVec_queue_4_deq_bits_readSource;
  wire [4:0]   sinkVec_2_0_bits_vs = sinkVec_sinkWire_4_bits_vs;
  wire [1:0]   sinkVec_queue_4_deq_bits_offset;
  wire [1:0]   sinkVec_2_0_bits_readSource = sinkVec_sinkWire_4_bits_readSource;
  wire [2:0]   sinkVec_queue_4_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_2_0_bits_offset = sinkVec_sinkWire_4_bits_offset;
  wire [2:0]   sinkVec_2_0_bits_instructionIndex = sinkVec_sinkWire_4_bits_instructionIndex;
  wire         sinkVec_validSink_4_valid;
  wire [4:0]   sinkVec_validSink_4_bits_vs;
  wire [1:0]   sinkVec_validSink_4_bits_readSource;
  wire [1:0]   sinkVec_validSink_4_bits_offset;
  wire [2:0]   sinkVec_validSink_4_bits_instructionIndex;
  assign sinkVec_sinkWire_4_valid = sinkVec_queue_4_deq_valid;
  assign sinkVec_sinkWire_4_bits_vs = sinkVec_queue_4_deq_bits_vs;
  assign sinkVec_sinkWire_4_bits_readSource = sinkVec_queue_4_deq_bits_readSource;
  assign sinkVec_sinkWire_4_bits_offset = sinkVec_queue_4_deq_bits_offset;
  assign sinkVec_sinkWire_4_bits_instructionIndex = sinkVec_queue_4_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_4_enq_bits_offset;
  wire [2:0]   sinkVec_queue_4_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_4 = {sinkVec_queue_4_enq_bits_offset, sinkVec_queue_4_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_4_enq_bits_vs;
  wire [1:0]   sinkVec_queue_4_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_4 = {sinkVec_queue_4_enq_bits_vs, sinkVec_queue_4_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_4 = {sinkVec_queue_dataIn_hi_4, sinkVec_queue_dataIn_lo_4};
  wire [2:0]   sinkVec_queue_dataOut_4_instructionIndex = _sinkVec_queue_fifo_4_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_4_offset = _sinkVec_queue_fifo_4_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_4_readSource = _sinkVec_queue_fifo_4_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_4_vs = _sinkVec_queue_fifo_4_data_out[11:7];
  wire         sinkVec_queue_4_enq_ready = ~_sinkVec_queue_fifo_4_full;
  wire         sinkVec_queue_4_enq_valid;
  assign sinkVec_queue_4_deq_valid = ~_sinkVec_queue_fifo_4_empty | sinkVec_queue_4_enq_valid;
  assign sinkVec_queue_4_deq_bits_vs = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_vs : sinkVec_queue_dataOut_4_vs;
  assign sinkVec_queue_4_deq_bits_readSource = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_readSource : sinkVec_queue_dataOut_4_readSource;
  assign sinkVec_queue_4_deq_bits_offset = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_offset : sinkVec_queue_dataOut_4_offset;
  assign sinkVec_queue_4_deq_bits_instructionIndex = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_instructionIndex : sinkVec_queue_dataOut_4_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_4;
  wire         sinkVec_releasePipe_pipe_out_4_valid = sinkVec_releasePipe_pipe_v_4;
  wire         x13_1_0_ready;
  wire         x13_1_0_valid;
  wire         sinkVec_validSource_4_valid = x13_1_0_ready & x13_1_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_4;
  wire [2:0]   sinkVec_tokenCheck_counterChange_4 = sinkVec_validSource_4_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_4 = ~(sinkVec_tokenCheck_counter_4[2]);
  assign x13_1_0_ready = sinkVec_tokenCheck_4;
  assign sinkVec_queue_4_enq_valid = sinkVec_validSink_4_valid;
  assign sinkVec_queue_4_enq_bits_vs = sinkVec_validSink_4_bits_vs;
  assign sinkVec_queue_4_enq_bits_readSource = sinkVec_validSink_4_bits_readSource;
  assign sinkVec_queue_4_enq_bits_offset = sinkVec_validSink_4_bits_offset;
  assign sinkVec_queue_4_enq_bits_instructionIndex = sinkVec_validSink_4_bits_instructionIndex;
  reg          sinkVec_shifterReg_4_0_valid;
  assign sinkVec_validSink_4_valid = sinkVec_shifterReg_4_0_valid;
  reg  [4:0]   sinkVec_shifterReg_4_0_bits_vs;
  assign sinkVec_validSink_4_bits_vs = sinkVec_shifterReg_4_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_4_0_bits_readSource;
  assign sinkVec_validSink_4_bits_readSource = sinkVec_shifterReg_4_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_4_0_bits_offset;
  assign sinkVec_validSink_4_bits_offset = sinkVec_shifterReg_4_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_4_0_bits_instructionIndex;
  assign sinkVec_validSink_4_bits_instructionIndex = sinkVec_shifterReg_4_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_4 = sinkVec_shifterReg_4_0_valid | sinkVec_validSource_4_valid;
  wire         sinkVec_2_1_ready;
  wire         sinkVec_queue_5_deq_ready = sinkVec_sinkWire_5_ready;
  wire         sinkVec_queue_5_deq_valid;
  wire [4:0]   sinkVec_queue_5_deq_bits_vs;
  wire         sinkVec_2_1_valid = sinkVec_sinkWire_5_valid;
  wire [1:0]   sinkVec_queue_5_deq_bits_readSource;
  wire [4:0]   sinkVec_2_1_bits_vs = sinkVec_sinkWire_5_bits_vs;
  wire [1:0]   sinkVec_queue_5_deq_bits_offset;
  wire [1:0]   sinkVec_2_1_bits_readSource = sinkVec_sinkWire_5_bits_readSource;
  wire [2:0]   sinkVec_queue_5_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_2_1_bits_offset = sinkVec_sinkWire_5_bits_offset;
  wire [2:0]   sinkVec_2_1_bits_instructionIndex = sinkVec_sinkWire_5_bits_instructionIndex;
  wire         sinkVec_validSink_5_valid;
  wire [4:0]   sinkVec_validSink_5_bits_vs;
  wire [1:0]   sinkVec_validSink_5_bits_readSource;
  wire [1:0]   sinkVec_validSink_5_bits_offset;
  wire [2:0]   sinkVec_validSink_5_bits_instructionIndex;
  assign sinkVec_sinkWire_5_valid = sinkVec_queue_5_deq_valid;
  assign sinkVec_sinkWire_5_bits_vs = sinkVec_queue_5_deq_bits_vs;
  assign sinkVec_sinkWire_5_bits_readSource = sinkVec_queue_5_deq_bits_readSource;
  assign sinkVec_sinkWire_5_bits_offset = sinkVec_queue_5_deq_bits_offset;
  assign sinkVec_sinkWire_5_bits_instructionIndex = sinkVec_queue_5_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_5_enq_bits_offset;
  wire [2:0]   sinkVec_queue_5_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_5 = {sinkVec_queue_5_enq_bits_offset, sinkVec_queue_5_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_5_enq_bits_vs;
  wire [1:0]   sinkVec_queue_5_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_5 = {sinkVec_queue_5_enq_bits_vs, sinkVec_queue_5_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_5 = {sinkVec_queue_dataIn_hi_5, sinkVec_queue_dataIn_lo_5};
  wire [2:0]   sinkVec_queue_dataOut_5_instructionIndex = _sinkVec_queue_fifo_5_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_5_offset = _sinkVec_queue_fifo_5_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_5_readSource = _sinkVec_queue_fifo_5_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_5_vs = _sinkVec_queue_fifo_5_data_out[11:7];
  wire         sinkVec_queue_5_enq_ready = ~_sinkVec_queue_fifo_5_full;
  wire         sinkVec_queue_5_enq_valid;
  assign sinkVec_queue_5_deq_valid = ~_sinkVec_queue_fifo_5_empty | sinkVec_queue_5_enq_valid;
  assign sinkVec_queue_5_deq_bits_vs = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_vs : sinkVec_queue_dataOut_5_vs;
  assign sinkVec_queue_5_deq_bits_readSource = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_readSource : sinkVec_queue_dataOut_5_readSource;
  assign sinkVec_queue_5_deq_bits_offset = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_offset : sinkVec_queue_dataOut_5_offset;
  assign sinkVec_queue_5_deq_bits_instructionIndex = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_instructionIndex : sinkVec_queue_dataOut_5_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_5;
  wire         sinkVec_releasePipe_pipe_out_5_valid = sinkVec_releasePipe_pipe_v_5;
  wire         x13_1_1_ready;
  wire         x13_1_1_valid;
  wire         sinkVec_validSource_5_valid = x13_1_1_ready & x13_1_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_5;
  wire [2:0]   sinkVec_tokenCheck_counterChange_5 = sinkVec_validSource_5_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_5 = ~(sinkVec_tokenCheck_counter_5[2]);
  assign x13_1_1_ready = sinkVec_tokenCheck_5;
  assign sinkVec_queue_5_enq_valid = sinkVec_validSink_5_valid;
  assign sinkVec_queue_5_enq_bits_vs = sinkVec_validSink_5_bits_vs;
  assign sinkVec_queue_5_enq_bits_readSource = sinkVec_validSink_5_bits_readSource;
  assign sinkVec_queue_5_enq_bits_offset = sinkVec_validSink_5_bits_offset;
  assign sinkVec_queue_5_enq_bits_instructionIndex = sinkVec_validSink_5_bits_instructionIndex;
  reg          sinkVec_shifterReg_5_0_valid;
  assign sinkVec_validSink_5_valid = sinkVec_shifterReg_5_0_valid;
  reg  [4:0]   sinkVec_shifterReg_5_0_bits_vs;
  assign sinkVec_validSink_5_bits_vs = sinkVec_shifterReg_5_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_5_0_bits_readSource;
  assign sinkVec_validSink_5_bits_readSource = sinkVec_shifterReg_5_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_5_0_bits_offset;
  assign sinkVec_validSink_5_bits_offset = sinkVec_shifterReg_5_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_5_0_bits_instructionIndex;
  assign sinkVec_validSink_5_bits_instructionIndex = sinkVec_shifterReg_5_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_5 = sinkVec_shifterReg_5_0_valid | sinkVec_validSource_5_valid;
  assign sinkVec_sinkWire_4_ready = sinkVec_2_0_ready;
  assign sinkVec_sinkWire_5_ready = sinkVec_2_1_ready;
  reg          maskUnitFirst_2;
  wire         tryToRead_2 = sinkVec_2_0_valid | sinkVec_2_1_valid;
  wire         sinkWire_2_valid = maskUnitFirst_2 ? sinkVec_2_0_valid : sinkVec_2_1_valid;
  wire [4:0]   sinkWire_2_bits_vs = maskUnitFirst_2 ? sinkVec_2_0_bits_vs : sinkVec_2_1_bits_vs;
  wire [1:0]   sinkWire_2_bits_readSource = maskUnitFirst_2 ? sinkVec_2_0_bits_readSource : sinkVec_2_1_bits_readSource;
  wire [1:0]   sinkWire_2_bits_offset = maskUnitFirst_2 ? sinkVec_2_0_bits_offset : sinkVec_2_1_bits_offset;
  wire [2:0]   sinkWire_2_bits_instructionIndex = maskUnitFirst_2 ? sinkVec_2_0_bits_instructionIndex : sinkVec_2_1_bits_instructionIndex;
  wire         sinkWire_2_ready;
  assign sinkVec_2_1_ready = sinkWire_2_ready & ~maskUnitFirst_2;
  assign sinkVec_2_0_ready = sinkWire_2_ready & maskUnitFirst_2;
  reg          accessDataValid_pipe_v_2;
  reg          accessDataValid_pipe_pipe_v_2;
  wire         accessDataValid_pipe_pipe_out_2_valid = accessDataValid_pipe_pipe_v_2;
  wire         accessDataSource_2_valid = accessDataValid_pipe_pipe_out_2_valid;
  reg          shifterReg_18_0_valid;
  reg  [31:0]  shifterReg_18_0_bits;
  wire         shifterValid_18 = shifterReg_18_0_valid | accessDataSource_2_valid;
  reg          accessDataValid_pipe_v_3;
  reg          accessDataValid_pipe_pipe_v_3;
  wire         accessDataValid_pipe_pipe_out_3_valid = accessDataValid_pipe_pipe_v_3;
  wire         accessDataSource_3_valid = accessDataValid_pipe_pipe_out_3_valid;
  reg          shifterReg_19_0_valid;
  reg  [31:0]  shifterReg_19_0_bits;
  wire         shifterValid_19 = shifterReg_19_0_valid | accessDataSource_3_valid;
  wire         sinkVec_tokenCheck_6;
  wire [4:0]   sinkVec_validSource_6_bits_vd = x22_1_0_bits_vd;
  wire [1:0]   sinkVec_validSource_6_bits_offset = x22_1_0_bits_offset;
  wire [3:0]   sinkVec_validSource_6_bits_mask = x22_1_0_bits_mask;
  wire [31:0]  sinkVec_validSource_6_bits_data = x22_1_0_bits_data;
  wire [2:0]   sinkVec_validSource_6_bits_instructionIndex = x22_1_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_7;
  wire [4:0]   sinkVec_validSource_7_bits_vd = x22_1_1_bits_vd;
  wire [1:0]   sinkVec_validSource_7_bits_offset = x22_1_1_bits_offset;
  wire [3:0]   sinkVec_validSource_7_bits_mask = x22_1_1_bits_mask;
  wire [31:0]  sinkVec_validSource_7_bits_data = x22_1_1_bits_data;
  wire         sinkVec_validSource_7_bits_last = x22_1_1_bits_last;
  wire [2:0]   sinkVec_validSource_7_bits_instructionIndex = x22_1_1_bits_instructionIndex;
  wire         sinkVec_3_0_ready;
  wire         sinkVec_queue_6_deq_ready = sinkVec_sinkWire_6_ready;
  wire         sinkVec_queue_6_deq_valid;
  wire [4:0]   sinkVec_queue_6_deq_bits_vd;
  wire         sinkVec_3_0_valid = sinkVec_sinkWire_6_valid;
  wire [1:0]   sinkVec_queue_6_deq_bits_offset;
  wire [4:0]   sinkVec_3_0_bits_vd = sinkVec_sinkWire_6_bits_vd;
  wire [3:0]   sinkVec_queue_6_deq_bits_mask;
  wire [1:0]   sinkVec_3_0_bits_offset = sinkVec_sinkWire_6_bits_offset;
  wire [31:0]  sinkVec_queue_6_deq_bits_data;
  wire [3:0]   sinkVec_3_0_bits_mask = sinkVec_sinkWire_6_bits_mask;
  wire         sinkVec_queue_6_deq_bits_last;
  wire [31:0]  sinkVec_3_0_bits_data = sinkVec_sinkWire_6_bits_data;
  wire [2:0]   sinkVec_queue_6_deq_bits_instructionIndex;
  wire         sinkVec_3_0_bits_last = sinkVec_sinkWire_6_bits_last;
  wire [2:0]   sinkVec_3_0_bits_instructionIndex = sinkVec_sinkWire_6_bits_instructionIndex;
  wire         sinkVec_validSink_6_valid;
  wire [4:0]   sinkVec_validSink_6_bits_vd;
  wire [1:0]   sinkVec_validSink_6_bits_offset;
  wire [3:0]   sinkVec_validSink_6_bits_mask;
  wire [31:0]  sinkVec_validSink_6_bits_data;
  wire [2:0]   sinkVec_validSink_6_bits_instructionIndex;
  assign sinkVec_sinkWire_6_valid = sinkVec_queue_6_deq_valid;
  assign sinkVec_sinkWire_6_bits_vd = sinkVec_queue_6_deq_bits_vd;
  assign sinkVec_sinkWire_6_bits_offset = sinkVec_queue_6_deq_bits_offset;
  assign sinkVec_sinkWire_6_bits_mask = sinkVec_queue_6_deq_bits_mask;
  assign sinkVec_sinkWire_6_bits_data = sinkVec_queue_6_deq_bits_data;
  assign sinkVec_sinkWire_6_bits_last = sinkVec_queue_6_deq_bits_last;
  assign sinkVec_sinkWire_6_bits_instructionIndex = sinkVec_queue_6_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_6_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_2 = {sinkVec_queue_6_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_6_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_6 = {sinkVec_queue_dataIn_lo_hi_2, sinkVec_queue_6_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_6_enq_bits_vd;
  wire [1:0]   sinkVec_queue_6_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_2 = {sinkVec_queue_6_enq_bits_vd, sinkVec_queue_6_enq_bits_offset};
  wire [3:0]   sinkVec_queue_6_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_6 = {sinkVec_queue_dataIn_hi_hi_2, sinkVec_queue_6_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_6 = {sinkVec_queue_dataIn_hi_6, sinkVec_queue_dataIn_lo_6};
  wire [2:0]   sinkVec_queue_dataOut_6_instructionIndex = _sinkVec_queue_fifo_6_data_out[2:0];
  wire         sinkVec_queue_dataOut_6_last = _sinkVec_queue_fifo_6_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_6_data = _sinkVec_queue_fifo_6_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_6_mask = _sinkVec_queue_fifo_6_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_6_offset = _sinkVec_queue_fifo_6_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_6_vd = _sinkVec_queue_fifo_6_data_out[46:42];
  wire         sinkVec_queue_6_enq_ready = ~_sinkVec_queue_fifo_6_full;
  wire         sinkVec_queue_6_enq_valid;
  assign sinkVec_queue_6_deq_valid = ~_sinkVec_queue_fifo_6_empty | sinkVec_queue_6_enq_valid;
  assign sinkVec_queue_6_deq_bits_vd = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_vd : sinkVec_queue_dataOut_6_vd;
  assign sinkVec_queue_6_deq_bits_offset = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_offset : sinkVec_queue_dataOut_6_offset;
  assign sinkVec_queue_6_deq_bits_mask = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_mask : sinkVec_queue_dataOut_6_mask;
  assign sinkVec_queue_6_deq_bits_data = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_data : sinkVec_queue_dataOut_6_data;
  assign sinkVec_queue_6_deq_bits_last = ~_sinkVec_queue_fifo_6_empty & sinkVec_queue_dataOut_6_last;
  assign sinkVec_queue_6_deq_bits_instructionIndex = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_instructionIndex : sinkVec_queue_dataOut_6_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_6;
  wire         sinkVec_releasePipe_pipe_out_6_valid = sinkVec_releasePipe_pipe_v_6;
  wire         x22_1_0_ready;
  wire         x22_1_0_valid;
  wire         sinkVec_validSource_6_valid = x22_1_0_ready & x22_1_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_6;
  wire [2:0]   sinkVec_tokenCheck_counterChange_6 = sinkVec_validSource_6_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_6 = ~(sinkVec_tokenCheck_counter_6[2]);
  assign x22_1_0_ready = sinkVec_tokenCheck_6;
  assign sinkVec_queue_6_enq_valid = sinkVec_validSink_6_valid;
  assign sinkVec_queue_6_enq_bits_vd = sinkVec_validSink_6_bits_vd;
  assign sinkVec_queue_6_enq_bits_offset = sinkVec_validSink_6_bits_offset;
  assign sinkVec_queue_6_enq_bits_mask = sinkVec_validSink_6_bits_mask;
  assign sinkVec_queue_6_enq_bits_data = sinkVec_validSink_6_bits_data;
  assign sinkVec_queue_6_enq_bits_instructionIndex = sinkVec_validSink_6_bits_instructionIndex;
  reg          sinkVec_shifterReg_6_0_valid;
  assign sinkVec_validSink_6_valid = sinkVec_shifterReg_6_0_valid;
  reg  [4:0]   sinkVec_shifterReg_6_0_bits_vd;
  assign sinkVec_validSink_6_bits_vd = sinkVec_shifterReg_6_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_6_0_bits_offset;
  assign sinkVec_validSink_6_bits_offset = sinkVec_shifterReg_6_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_6_0_bits_mask;
  assign sinkVec_validSink_6_bits_mask = sinkVec_shifterReg_6_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_6_0_bits_data;
  assign sinkVec_validSink_6_bits_data = sinkVec_shifterReg_6_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_6_0_bits_instructionIndex;
  assign sinkVec_validSink_6_bits_instructionIndex = sinkVec_shifterReg_6_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_6 = sinkVec_shifterReg_6_0_valid | sinkVec_validSource_6_valid;
  wire         sinkVec_3_1_ready;
  wire         sinkVec_queue_7_deq_ready = sinkVec_sinkWire_7_ready;
  wire         sinkVec_queue_7_deq_valid;
  wire [4:0]   sinkVec_queue_7_deq_bits_vd;
  wire         sinkVec_3_1_valid = sinkVec_sinkWire_7_valid;
  wire [1:0]   sinkVec_queue_7_deq_bits_offset;
  wire [4:0]   sinkVec_3_1_bits_vd = sinkVec_sinkWire_7_bits_vd;
  wire [3:0]   sinkVec_queue_7_deq_bits_mask;
  wire [1:0]   sinkVec_3_1_bits_offset = sinkVec_sinkWire_7_bits_offset;
  wire [31:0]  sinkVec_queue_7_deq_bits_data;
  wire [3:0]   sinkVec_3_1_bits_mask = sinkVec_sinkWire_7_bits_mask;
  wire         sinkVec_queue_7_deq_bits_last;
  wire [31:0]  sinkVec_3_1_bits_data = sinkVec_sinkWire_7_bits_data;
  wire [2:0]   sinkVec_queue_7_deq_bits_instructionIndex;
  wire         sinkVec_3_1_bits_last = sinkVec_sinkWire_7_bits_last;
  wire [2:0]   sinkVec_3_1_bits_instructionIndex = sinkVec_sinkWire_7_bits_instructionIndex;
  wire         sinkVec_validSink_7_valid;
  wire [4:0]   sinkVec_validSink_7_bits_vd;
  wire [1:0]   sinkVec_validSink_7_bits_offset;
  wire [3:0]   sinkVec_validSink_7_bits_mask;
  wire [31:0]  sinkVec_validSink_7_bits_data;
  wire         sinkVec_validSink_7_bits_last;
  wire [2:0]   sinkVec_validSink_7_bits_instructionIndex;
  assign sinkVec_sinkWire_7_valid = sinkVec_queue_7_deq_valid;
  assign sinkVec_sinkWire_7_bits_vd = sinkVec_queue_7_deq_bits_vd;
  assign sinkVec_sinkWire_7_bits_offset = sinkVec_queue_7_deq_bits_offset;
  assign sinkVec_sinkWire_7_bits_mask = sinkVec_queue_7_deq_bits_mask;
  assign sinkVec_sinkWire_7_bits_data = sinkVec_queue_7_deq_bits_data;
  assign sinkVec_sinkWire_7_bits_last = sinkVec_queue_7_deq_bits_last;
  assign sinkVec_sinkWire_7_bits_instructionIndex = sinkVec_queue_7_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_7_enq_bits_data;
  wire         sinkVec_queue_7_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_3 = {sinkVec_queue_7_enq_bits_data, sinkVec_queue_7_enq_bits_last};
  wire [2:0]   sinkVec_queue_7_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_7 = {sinkVec_queue_dataIn_lo_hi_3, sinkVec_queue_7_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_7_enq_bits_vd;
  wire [1:0]   sinkVec_queue_7_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_3 = {sinkVec_queue_7_enq_bits_vd, sinkVec_queue_7_enq_bits_offset};
  wire [3:0]   sinkVec_queue_7_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_7 = {sinkVec_queue_dataIn_hi_hi_3, sinkVec_queue_7_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_7 = {sinkVec_queue_dataIn_hi_7, sinkVec_queue_dataIn_lo_7};
  wire [2:0]   sinkVec_queue_dataOut_7_instructionIndex = _sinkVec_queue_fifo_7_data_out[2:0];
  wire         sinkVec_queue_dataOut_7_last = _sinkVec_queue_fifo_7_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_7_data = _sinkVec_queue_fifo_7_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_7_mask = _sinkVec_queue_fifo_7_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_7_offset = _sinkVec_queue_fifo_7_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_7_vd = _sinkVec_queue_fifo_7_data_out[46:42];
  wire         sinkVec_queue_7_enq_ready = ~_sinkVec_queue_fifo_7_full;
  wire         sinkVec_queue_7_enq_valid;
  assign sinkVec_queue_7_deq_valid = ~_sinkVec_queue_fifo_7_empty | sinkVec_queue_7_enq_valid;
  assign sinkVec_queue_7_deq_bits_vd = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_vd : sinkVec_queue_dataOut_7_vd;
  assign sinkVec_queue_7_deq_bits_offset = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_offset : sinkVec_queue_dataOut_7_offset;
  assign sinkVec_queue_7_deq_bits_mask = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_mask : sinkVec_queue_dataOut_7_mask;
  assign sinkVec_queue_7_deq_bits_data = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_data : sinkVec_queue_dataOut_7_data;
  assign sinkVec_queue_7_deq_bits_last = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_last : sinkVec_queue_dataOut_7_last;
  assign sinkVec_queue_7_deq_bits_instructionIndex = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_instructionIndex : sinkVec_queue_dataOut_7_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_7;
  wire         sinkVec_releasePipe_pipe_out_7_valid = sinkVec_releasePipe_pipe_v_7;
  wire         x22_1_1_ready;
  wire         x22_1_1_valid;
  wire         sinkVec_validSource_7_valid = x22_1_1_ready & x22_1_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_7;
  wire [2:0]   sinkVec_tokenCheck_counterChange_7 = sinkVec_validSource_7_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_7 = ~(sinkVec_tokenCheck_counter_7[2]);
  assign x22_1_1_ready = sinkVec_tokenCheck_7;
  assign sinkVec_queue_7_enq_valid = sinkVec_validSink_7_valid;
  assign sinkVec_queue_7_enq_bits_vd = sinkVec_validSink_7_bits_vd;
  assign sinkVec_queue_7_enq_bits_offset = sinkVec_validSink_7_bits_offset;
  assign sinkVec_queue_7_enq_bits_mask = sinkVec_validSink_7_bits_mask;
  assign sinkVec_queue_7_enq_bits_data = sinkVec_validSink_7_bits_data;
  assign sinkVec_queue_7_enq_bits_last = sinkVec_validSink_7_bits_last;
  assign sinkVec_queue_7_enq_bits_instructionIndex = sinkVec_validSink_7_bits_instructionIndex;
  reg          sinkVec_shifterReg_7_0_valid;
  assign sinkVec_validSink_7_valid = sinkVec_shifterReg_7_0_valid;
  reg  [4:0]   sinkVec_shifterReg_7_0_bits_vd;
  assign sinkVec_validSink_7_bits_vd = sinkVec_shifterReg_7_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_7_0_bits_offset;
  assign sinkVec_validSink_7_bits_offset = sinkVec_shifterReg_7_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_7_0_bits_mask;
  assign sinkVec_validSink_7_bits_mask = sinkVec_shifterReg_7_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_7_0_bits_data;
  assign sinkVec_validSink_7_bits_data = sinkVec_shifterReg_7_0_bits_data;
  reg          sinkVec_shifterReg_7_0_bits_last;
  assign sinkVec_validSink_7_bits_last = sinkVec_shifterReg_7_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_7_0_bits_instructionIndex;
  assign sinkVec_validSink_7_bits_instructionIndex = sinkVec_shifterReg_7_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_7 = sinkVec_shifterReg_7_0_valid | sinkVec_validSource_7_valid;
  assign sinkVec_sinkWire_6_ready = sinkVec_3_0_ready;
  assign sinkVec_sinkWire_7_ready = sinkVec_3_1_ready;
  reg          maskUnitFirst_3;
  wire         tryToRead_3 = sinkVec_3_0_valid | sinkVec_3_1_valid;
  wire         sinkWire_3_valid = maskUnitFirst_3 ? sinkVec_3_0_valid : sinkVec_3_1_valid;
  wire [4:0]   sinkWire_3_bits_vd = maskUnitFirst_3 ? sinkVec_3_0_bits_vd : sinkVec_3_1_bits_vd;
  wire [1:0]   sinkWire_3_bits_offset = maskUnitFirst_3 ? sinkVec_3_0_bits_offset : sinkVec_3_1_bits_offset;
  wire [3:0]   sinkWire_3_bits_mask = maskUnitFirst_3 ? sinkVec_3_0_bits_mask : sinkVec_3_1_bits_mask;
  wire [31:0]  sinkWire_3_bits_data = maskUnitFirst_3 ? sinkVec_3_0_bits_data : sinkVec_3_1_bits_data;
  wire         sinkWire_3_bits_last = maskUnitFirst_3 ? sinkVec_3_0_bits_last : sinkVec_3_1_bits_last;
  wire [2:0]   sinkWire_3_bits_instructionIndex = maskUnitFirst_3 ? sinkVec_3_0_bits_instructionIndex : sinkVec_3_1_bits_instructionIndex;
  wire         sinkWire_3_ready;
  assign sinkVec_3_1_ready = sinkWire_3_ready & ~maskUnitFirst_3;
  assign sinkVec_3_0_ready = sinkWire_3_ready & maskUnitFirst_3;
  reg          view__writeRelease_1_pipe_v;
  wire         view__writeRelease_1_pipe_out_valid = view__writeRelease_1_pipe_v;
  reg          pipe_v_3;
  wire         pipe_out_2_valid = pipe_v_3;
  wire         _probeWire_writeQueueEnqVec_1_valid_T = x22_1_0_ready & _maskUnit_exeResp_1_valid;
  reg          instructionFinishedPipe_pipe_v_1;
  wire         instructionFinishedPipe_pipe_out_1_valid = instructionFinishedPipe_pipe_v_1;
  reg  [7:0]   instructionFinishedPipe_pipe_b_1;
  wire [7:0]   instructionFinishedPipe_pipe_out_1_bits = instructionFinishedPipe_pipe_b_1;
  wire         instructionFinished_1_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_1_bits);
  assign vxsatReportVec_1 = _laneVec_1_vxsatReport[3:0];
  reg          pipe_v_4;
  reg  [31:0]  pipe_b_4;
  reg          pipe_pipe_v_1;
  wire         pipe_pipe_out_1_valid = pipe_pipe_v_1;
  reg  [31:0]  pipe_pipe_b_1;
  wire [31:0]  pipe_pipe_out_1_bits = pipe_pipe_b_1;
  reg          view__laneMaskSelect_1_pipe_v;
  reg  [5:0]   view__laneMaskSelect_1_pipe_b;
  reg          view__laneMaskSelect_1_pipe_pipe_v;
  wire         view__laneMaskSelect_1_pipe_pipe_out_valid = view__laneMaskSelect_1_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_1_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_1_pipe_pipe_out_bits = view__laneMaskSelect_1_pipe_pipe_b;
  reg          view__laneMaskSewSelect_1_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_1_pipe_b;
  reg          view__laneMaskSewSelect_1_pipe_pipe_v;
  wire         view__laneMaskSewSelect_1_pipe_pipe_out_valid = view__laneMaskSewSelect_1_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_1_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_1_pipe_pipe_out_bits = view__laneMaskSewSelect_1_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_1;
  wire         lsuLastPipe_pipe_out_1_valid = lsuLastPipe_pipe_v_1;
  reg  [7:0]   lsuLastPipe_pipe_b_1;
  wire [7:0]   lsuLastPipe_pipe_out_1_bits = lsuLastPipe_pipe_b_1;
  reg          maskLastPipe_pipe_v_1;
  wire         maskLastPipe_pipe_out_1_valid = maskLastPipe_pipe_v_1;
  reg  [7:0]   maskLastPipe_pipe_b_1;
  wire [7:0]   maskLastPipe_pipe_out_1_bits = maskLastPipe_pipe_b_1;
  wire [5:0]   writeCounter_1 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h4};
  reg          pipe_v_5;
  wire         pipe_out_3_valid = pipe_v_5;
  reg  [5:0]   pipe_b_5;
  wire [5:0]   pipe_out_3_bits = pipe_b_5;
  assign laneRequestSinkWire_2_ready = ~laneRequestSinkWire_2_bits_issueInst | _laneVec_2_laneRequest_ready;
  wire         sinkVec_tokenCheck_8;
  wire [4:0]   sinkVec_validSource_8_bits_vs = x13_2_0_bits_vs;
  wire [1:0]   sinkVec_validSource_8_bits_offset = x13_2_0_bits_offset;
  wire [2:0]   sinkVec_validSource_8_bits_instructionIndex = x13_2_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_9;
  wire [4:0]   sinkVec_validSource_9_bits_vs = x13_2_1_bits_vs;
  wire [1:0]   sinkVec_validSource_9_bits_offset = x13_2_1_bits_offset;
  wire [2:0]   sinkVec_validSource_9_bits_instructionIndex = x13_2_1_bits_instructionIndex;
  wire         sinkVec_4_0_ready;
  wire         sinkVec_queue_8_deq_ready = sinkVec_sinkWire_8_ready;
  wire         sinkVec_queue_8_deq_valid;
  wire [4:0]   sinkVec_queue_8_deq_bits_vs;
  wire         sinkVec_4_0_valid = sinkVec_sinkWire_8_valid;
  wire [1:0]   sinkVec_queue_8_deq_bits_readSource;
  wire [4:0]   sinkVec_4_0_bits_vs = sinkVec_sinkWire_8_bits_vs;
  wire [1:0]   sinkVec_queue_8_deq_bits_offset;
  wire [1:0]   sinkVec_4_0_bits_readSource = sinkVec_sinkWire_8_bits_readSource;
  wire [2:0]   sinkVec_queue_8_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_4_0_bits_offset = sinkVec_sinkWire_8_bits_offset;
  wire [2:0]   sinkVec_4_0_bits_instructionIndex = sinkVec_sinkWire_8_bits_instructionIndex;
  wire         sinkVec_validSink_8_valid;
  wire [4:0]   sinkVec_validSink_8_bits_vs;
  wire [1:0]   sinkVec_validSink_8_bits_readSource;
  wire [1:0]   sinkVec_validSink_8_bits_offset;
  wire [2:0]   sinkVec_validSink_8_bits_instructionIndex;
  assign sinkVec_sinkWire_8_valid = sinkVec_queue_8_deq_valid;
  assign sinkVec_sinkWire_8_bits_vs = sinkVec_queue_8_deq_bits_vs;
  assign sinkVec_sinkWire_8_bits_readSource = sinkVec_queue_8_deq_bits_readSource;
  assign sinkVec_sinkWire_8_bits_offset = sinkVec_queue_8_deq_bits_offset;
  assign sinkVec_sinkWire_8_bits_instructionIndex = sinkVec_queue_8_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_8_enq_bits_offset;
  wire [2:0]   sinkVec_queue_8_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_8 = {sinkVec_queue_8_enq_bits_offset, sinkVec_queue_8_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_8_enq_bits_vs;
  wire [1:0]   sinkVec_queue_8_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_8 = {sinkVec_queue_8_enq_bits_vs, sinkVec_queue_8_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_8 = {sinkVec_queue_dataIn_hi_8, sinkVec_queue_dataIn_lo_8};
  wire [2:0]   sinkVec_queue_dataOut_8_instructionIndex = _sinkVec_queue_fifo_8_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_8_offset = _sinkVec_queue_fifo_8_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_8_readSource = _sinkVec_queue_fifo_8_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_8_vs = _sinkVec_queue_fifo_8_data_out[11:7];
  wire         sinkVec_queue_8_enq_ready = ~_sinkVec_queue_fifo_8_full;
  wire         sinkVec_queue_8_enq_valid;
  assign sinkVec_queue_8_deq_valid = ~_sinkVec_queue_fifo_8_empty | sinkVec_queue_8_enq_valid;
  assign sinkVec_queue_8_deq_bits_vs = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_vs : sinkVec_queue_dataOut_8_vs;
  assign sinkVec_queue_8_deq_bits_readSource = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_readSource : sinkVec_queue_dataOut_8_readSource;
  assign sinkVec_queue_8_deq_bits_offset = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_offset : sinkVec_queue_dataOut_8_offset;
  assign sinkVec_queue_8_deq_bits_instructionIndex = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_instructionIndex : sinkVec_queue_dataOut_8_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_8;
  wire         sinkVec_releasePipe_pipe_out_8_valid = sinkVec_releasePipe_pipe_v_8;
  wire         x13_2_0_ready;
  wire         x13_2_0_valid;
  wire         sinkVec_validSource_8_valid = x13_2_0_ready & x13_2_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_8;
  wire [2:0]   sinkVec_tokenCheck_counterChange_8 = sinkVec_validSource_8_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_8 = ~(sinkVec_tokenCheck_counter_8[2]);
  assign x13_2_0_ready = sinkVec_tokenCheck_8;
  assign sinkVec_queue_8_enq_valid = sinkVec_validSink_8_valid;
  assign sinkVec_queue_8_enq_bits_vs = sinkVec_validSink_8_bits_vs;
  assign sinkVec_queue_8_enq_bits_readSource = sinkVec_validSink_8_bits_readSource;
  assign sinkVec_queue_8_enq_bits_offset = sinkVec_validSink_8_bits_offset;
  assign sinkVec_queue_8_enq_bits_instructionIndex = sinkVec_validSink_8_bits_instructionIndex;
  reg          sinkVec_shifterReg_8_0_valid;
  assign sinkVec_validSink_8_valid = sinkVec_shifterReg_8_0_valid;
  reg  [4:0]   sinkVec_shifterReg_8_0_bits_vs;
  assign sinkVec_validSink_8_bits_vs = sinkVec_shifterReg_8_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_8_0_bits_readSource;
  assign sinkVec_validSink_8_bits_readSource = sinkVec_shifterReg_8_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_8_0_bits_offset;
  assign sinkVec_validSink_8_bits_offset = sinkVec_shifterReg_8_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_8_0_bits_instructionIndex;
  assign sinkVec_validSink_8_bits_instructionIndex = sinkVec_shifterReg_8_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_8 = sinkVec_shifterReg_8_0_valid | sinkVec_validSource_8_valid;
  wire         sinkVec_4_1_ready;
  wire         sinkVec_queue_9_deq_ready = sinkVec_sinkWire_9_ready;
  wire         sinkVec_queue_9_deq_valid;
  wire [4:0]   sinkVec_queue_9_deq_bits_vs;
  wire         sinkVec_4_1_valid = sinkVec_sinkWire_9_valid;
  wire [1:0]   sinkVec_queue_9_deq_bits_readSource;
  wire [4:0]   sinkVec_4_1_bits_vs = sinkVec_sinkWire_9_bits_vs;
  wire [1:0]   sinkVec_queue_9_deq_bits_offset;
  wire [1:0]   sinkVec_4_1_bits_readSource = sinkVec_sinkWire_9_bits_readSource;
  wire [2:0]   sinkVec_queue_9_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_4_1_bits_offset = sinkVec_sinkWire_9_bits_offset;
  wire [2:0]   sinkVec_4_1_bits_instructionIndex = sinkVec_sinkWire_9_bits_instructionIndex;
  wire         sinkVec_validSink_9_valid;
  wire [4:0]   sinkVec_validSink_9_bits_vs;
  wire [1:0]   sinkVec_validSink_9_bits_readSource;
  wire [1:0]   sinkVec_validSink_9_bits_offset;
  wire [2:0]   sinkVec_validSink_9_bits_instructionIndex;
  assign sinkVec_sinkWire_9_valid = sinkVec_queue_9_deq_valid;
  assign sinkVec_sinkWire_9_bits_vs = sinkVec_queue_9_deq_bits_vs;
  assign sinkVec_sinkWire_9_bits_readSource = sinkVec_queue_9_deq_bits_readSource;
  assign sinkVec_sinkWire_9_bits_offset = sinkVec_queue_9_deq_bits_offset;
  assign sinkVec_sinkWire_9_bits_instructionIndex = sinkVec_queue_9_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_9_enq_bits_offset;
  wire [2:0]   sinkVec_queue_9_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_9 = {sinkVec_queue_9_enq_bits_offset, sinkVec_queue_9_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_9_enq_bits_vs;
  wire [1:0]   sinkVec_queue_9_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_9 = {sinkVec_queue_9_enq_bits_vs, sinkVec_queue_9_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_9 = {sinkVec_queue_dataIn_hi_9, sinkVec_queue_dataIn_lo_9};
  wire [2:0]   sinkVec_queue_dataOut_9_instructionIndex = _sinkVec_queue_fifo_9_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_9_offset = _sinkVec_queue_fifo_9_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_9_readSource = _sinkVec_queue_fifo_9_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_9_vs = _sinkVec_queue_fifo_9_data_out[11:7];
  wire         sinkVec_queue_9_enq_ready = ~_sinkVec_queue_fifo_9_full;
  wire         sinkVec_queue_9_enq_valid;
  assign sinkVec_queue_9_deq_valid = ~_sinkVec_queue_fifo_9_empty | sinkVec_queue_9_enq_valid;
  assign sinkVec_queue_9_deq_bits_vs = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_vs : sinkVec_queue_dataOut_9_vs;
  assign sinkVec_queue_9_deq_bits_readSource = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_readSource : sinkVec_queue_dataOut_9_readSource;
  assign sinkVec_queue_9_deq_bits_offset = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_offset : sinkVec_queue_dataOut_9_offset;
  assign sinkVec_queue_9_deq_bits_instructionIndex = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_instructionIndex : sinkVec_queue_dataOut_9_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_9;
  wire         sinkVec_releasePipe_pipe_out_9_valid = sinkVec_releasePipe_pipe_v_9;
  wire         x13_2_1_ready;
  wire         x13_2_1_valid;
  wire         sinkVec_validSource_9_valid = x13_2_1_ready & x13_2_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_9;
  wire [2:0]   sinkVec_tokenCheck_counterChange_9 = sinkVec_validSource_9_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_9 = ~(sinkVec_tokenCheck_counter_9[2]);
  assign x13_2_1_ready = sinkVec_tokenCheck_9;
  assign sinkVec_queue_9_enq_valid = sinkVec_validSink_9_valid;
  assign sinkVec_queue_9_enq_bits_vs = sinkVec_validSink_9_bits_vs;
  assign sinkVec_queue_9_enq_bits_readSource = sinkVec_validSink_9_bits_readSource;
  assign sinkVec_queue_9_enq_bits_offset = sinkVec_validSink_9_bits_offset;
  assign sinkVec_queue_9_enq_bits_instructionIndex = sinkVec_validSink_9_bits_instructionIndex;
  reg          sinkVec_shifterReg_9_0_valid;
  assign sinkVec_validSink_9_valid = sinkVec_shifterReg_9_0_valid;
  reg  [4:0]   sinkVec_shifterReg_9_0_bits_vs;
  assign sinkVec_validSink_9_bits_vs = sinkVec_shifterReg_9_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_9_0_bits_readSource;
  assign sinkVec_validSink_9_bits_readSource = sinkVec_shifterReg_9_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_9_0_bits_offset;
  assign sinkVec_validSink_9_bits_offset = sinkVec_shifterReg_9_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_9_0_bits_instructionIndex;
  assign sinkVec_validSink_9_bits_instructionIndex = sinkVec_shifterReg_9_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_9 = sinkVec_shifterReg_9_0_valid | sinkVec_validSource_9_valid;
  assign sinkVec_sinkWire_8_ready = sinkVec_4_0_ready;
  assign sinkVec_sinkWire_9_ready = sinkVec_4_1_ready;
  reg          maskUnitFirst_4;
  wire         tryToRead_4 = sinkVec_4_0_valid | sinkVec_4_1_valid;
  wire         sinkWire_4_valid = maskUnitFirst_4 ? sinkVec_4_0_valid : sinkVec_4_1_valid;
  wire [4:0]   sinkWire_4_bits_vs = maskUnitFirst_4 ? sinkVec_4_0_bits_vs : sinkVec_4_1_bits_vs;
  wire [1:0]   sinkWire_4_bits_readSource = maskUnitFirst_4 ? sinkVec_4_0_bits_readSource : sinkVec_4_1_bits_readSource;
  wire [1:0]   sinkWire_4_bits_offset = maskUnitFirst_4 ? sinkVec_4_0_bits_offset : sinkVec_4_1_bits_offset;
  wire [2:0]   sinkWire_4_bits_instructionIndex = maskUnitFirst_4 ? sinkVec_4_0_bits_instructionIndex : sinkVec_4_1_bits_instructionIndex;
  wire         sinkWire_4_ready;
  assign sinkVec_4_1_ready = sinkWire_4_ready & ~maskUnitFirst_4;
  assign sinkVec_4_0_ready = sinkWire_4_ready & maskUnitFirst_4;
  reg          accessDataValid_pipe_v_4;
  reg          accessDataValid_pipe_pipe_v_4;
  wire         accessDataValid_pipe_pipe_out_4_valid = accessDataValid_pipe_pipe_v_4;
  wire         accessDataSource_4_valid = accessDataValid_pipe_pipe_out_4_valid;
  reg          shifterReg_20_0_valid;
  reg  [31:0]  shifterReg_20_0_bits;
  wire         shifterValid_20 = shifterReg_20_0_valid | accessDataSource_4_valid;
  reg          accessDataValid_pipe_v_5;
  reg          accessDataValid_pipe_pipe_v_5;
  wire         accessDataValid_pipe_pipe_out_5_valid = accessDataValid_pipe_pipe_v_5;
  wire         accessDataSource_5_valid = accessDataValid_pipe_pipe_out_5_valid;
  reg          shifterReg_21_0_valid;
  reg  [31:0]  shifterReg_21_0_bits;
  wire         shifterValid_21 = shifterReg_21_0_valid | accessDataSource_5_valid;
  wire         sinkVec_tokenCheck_10;
  wire [4:0]   sinkVec_validSource_10_bits_vd = x22_2_0_bits_vd;
  wire [1:0]   sinkVec_validSource_10_bits_offset = x22_2_0_bits_offset;
  wire [3:0]   sinkVec_validSource_10_bits_mask = x22_2_0_bits_mask;
  wire [31:0]  sinkVec_validSource_10_bits_data = x22_2_0_bits_data;
  wire [2:0]   sinkVec_validSource_10_bits_instructionIndex = x22_2_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_11;
  wire [4:0]   sinkVec_validSource_11_bits_vd = x22_2_1_bits_vd;
  wire [1:0]   sinkVec_validSource_11_bits_offset = x22_2_1_bits_offset;
  wire [3:0]   sinkVec_validSource_11_bits_mask = x22_2_1_bits_mask;
  wire [31:0]  sinkVec_validSource_11_bits_data = x22_2_1_bits_data;
  wire         sinkVec_validSource_11_bits_last = x22_2_1_bits_last;
  wire [2:0]   sinkVec_validSource_11_bits_instructionIndex = x22_2_1_bits_instructionIndex;
  wire         sinkVec_5_0_ready;
  wire         sinkVec_queue_10_deq_ready = sinkVec_sinkWire_10_ready;
  wire         sinkVec_queue_10_deq_valid;
  wire [4:0]   sinkVec_queue_10_deq_bits_vd;
  wire         sinkVec_5_0_valid = sinkVec_sinkWire_10_valid;
  wire [1:0]   sinkVec_queue_10_deq_bits_offset;
  wire [4:0]   sinkVec_5_0_bits_vd = sinkVec_sinkWire_10_bits_vd;
  wire [3:0]   sinkVec_queue_10_deq_bits_mask;
  wire [1:0]   sinkVec_5_0_bits_offset = sinkVec_sinkWire_10_bits_offset;
  wire [31:0]  sinkVec_queue_10_deq_bits_data;
  wire [3:0]   sinkVec_5_0_bits_mask = sinkVec_sinkWire_10_bits_mask;
  wire         sinkVec_queue_10_deq_bits_last;
  wire [31:0]  sinkVec_5_0_bits_data = sinkVec_sinkWire_10_bits_data;
  wire [2:0]   sinkVec_queue_10_deq_bits_instructionIndex;
  wire         sinkVec_5_0_bits_last = sinkVec_sinkWire_10_bits_last;
  wire [2:0]   sinkVec_5_0_bits_instructionIndex = sinkVec_sinkWire_10_bits_instructionIndex;
  wire         sinkVec_validSink_10_valid;
  wire [4:0]   sinkVec_validSink_10_bits_vd;
  wire [1:0]   sinkVec_validSink_10_bits_offset;
  wire [3:0]   sinkVec_validSink_10_bits_mask;
  wire [31:0]  sinkVec_validSink_10_bits_data;
  wire [2:0]   sinkVec_validSink_10_bits_instructionIndex;
  assign sinkVec_sinkWire_10_valid = sinkVec_queue_10_deq_valid;
  assign sinkVec_sinkWire_10_bits_vd = sinkVec_queue_10_deq_bits_vd;
  assign sinkVec_sinkWire_10_bits_offset = sinkVec_queue_10_deq_bits_offset;
  assign sinkVec_sinkWire_10_bits_mask = sinkVec_queue_10_deq_bits_mask;
  assign sinkVec_sinkWire_10_bits_data = sinkVec_queue_10_deq_bits_data;
  assign sinkVec_sinkWire_10_bits_last = sinkVec_queue_10_deq_bits_last;
  assign sinkVec_sinkWire_10_bits_instructionIndex = sinkVec_queue_10_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_10_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_4 = {sinkVec_queue_10_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_10_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_10 = {sinkVec_queue_dataIn_lo_hi_4, sinkVec_queue_10_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_10_enq_bits_vd;
  wire [1:0]   sinkVec_queue_10_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_4 = {sinkVec_queue_10_enq_bits_vd, sinkVec_queue_10_enq_bits_offset};
  wire [3:0]   sinkVec_queue_10_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_10 = {sinkVec_queue_dataIn_hi_hi_4, sinkVec_queue_10_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_10 = {sinkVec_queue_dataIn_hi_10, sinkVec_queue_dataIn_lo_10};
  wire [2:0]   sinkVec_queue_dataOut_10_instructionIndex = _sinkVec_queue_fifo_10_data_out[2:0];
  wire         sinkVec_queue_dataOut_10_last = _sinkVec_queue_fifo_10_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_10_data = _sinkVec_queue_fifo_10_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_10_mask = _sinkVec_queue_fifo_10_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_10_offset = _sinkVec_queue_fifo_10_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_10_vd = _sinkVec_queue_fifo_10_data_out[46:42];
  wire         sinkVec_queue_10_enq_ready = ~_sinkVec_queue_fifo_10_full;
  wire         sinkVec_queue_10_enq_valid;
  assign sinkVec_queue_10_deq_valid = ~_sinkVec_queue_fifo_10_empty | sinkVec_queue_10_enq_valid;
  assign sinkVec_queue_10_deq_bits_vd = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_vd : sinkVec_queue_dataOut_10_vd;
  assign sinkVec_queue_10_deq_bits_offset = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_offset : sinkVec_queue_dataOut_10_offset;
  assign sinkVec_queue_10_deq_bits_mask = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_mask : sinkVec_queue_dataOut_10_mask;
  assign sinkVec_queue_10_deq_bits_data = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_data : sinkVec_queue_dataOut_10_data;
  assign sinkVec_queue_10_deq_bits_last = ~_sinkVec_queue_fifo_10_empty & sinkVec_queue_dataOut_10_last;
  assign sinkVec_queue_10_deq_bits_instructionIndex = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_instructionIndex : sinkVec_queue_dataOut_10_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_10;
  wire         sinkVec_releasePipe_pipe_out_10_valid = sinkVec_releasePipe_pipe_v_10;
  wire         x22_2_0_ready;
  wire         x22_2_0_valid;
  wire         sinkVec_validSource_10_valid = x22_2_0_ready & x22_2_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_10;
  wire [2:0]   sinkVec_tokenCheck_counterChange_10 = sinkVec_validSource_10_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_10 = ~(sinkVec_tokenCheck_counter_10[2]);
  assign x22_2_0_ready = sinkVec_tokenCheck_10;
  assign sinkVec_queue_10_enq_valid = sinkVec_validSink_10_valid;
  assign sinkVec_queue_10_enq_bits_vd = sinkVec_validSink_10_bits_vd;
  assign sinkVec_queue_10_enq_bits_offset = sinkVec_validSink_10_bits_offset;
  assign sinkVec_queue_10_enq_bits_mask = sinkVec_validSink_10_bits_mask;
  assign sinkVec_queue_10_enq_bits_data = sinkVec_validSink_10_bits_data;
  assign sinkVec_queue_10_enq_bits_instructionIndex = sinkVec_validSink_10_bits_instructionIndex;
  reg          sinkVec_shifterReg_10_0_valid;
  assign sinkVec_validSink_10_valid = sinkVec_shifterReg_10_0_valid;
  reg  [4:0]   sinkVec_shifterReg_10_0_bits_vd;
  assign sinkVec_validSink_10_bits_vd = sinkVec_shifterReg_10_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_10_0_bits_offset;
  assign sinkVec_validSink_10_bits_offset = sinkVec_shifterReg_10_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_10_0_bits_mask;
  assign sinkVec_validSink_10_bits_mask = sinkVec_shifterReg_10_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_10_0_bits_data;
  assign sinkVec_validSink_10_bits_data = sinkVec_shifterReg_10_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_10_0_bits_instructionIndex;
  assign sinkVec_validSink_10_bits_instructionIndex = sinkVec_shifterReg_10_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_10 = sinkVec_shifterReg_10_0_valid | sinkVec_validSource_10_valid;
  wire         sinkVec_5_1_ready;
  wire         sinkVec_queue_11_deq_ready = sinkVec_sinkWire_11_ready;
  wire         sinkVec_queue_11_deq_valid;
  wire [4:0]   sinkVec_queue_11_deq_bits_vd;
  wire         sinkVec_5_1_valid = sinkVec_sinkWire_11_valid;
  wire [1:0]   sinkVec_queue_11_deq_bits_offset;
  wire [4:0]   sinkVec_5_1_bits_vd = sinkVec_sinkWire_11_bits_vd;
  wire [3:0]   sinkVec_queue_11_deq_bits_mask;
  wire [1:0]   sinkVec_5_1_bits_offset = sinkVec_sinkWire_11_bits_offset;
  wire [31:0]  sinkVec_queue_11_deq_bits_data;
  wire [3:0]   sinkVec_5_1_bits_mask = sinkVec_sinkWire_11_bits_mask;
  wire         sinkVec_queue_11_deq_bits_last;
  wire [31:0]  sinkVec_5_1_bits_data = sinkVec_sinkWire_11_bits_data;
  wire [2:0]   sinkVec_queue_11_deq_bits_instructionIndex;
  wire         sinkVec_5_1_bits_last = sinkVec_sinkWire_11_bits_last;
  wire [2:0]   sinkVec_5_1_bits_instructionIndex = sinkVec_sinkWire_11_bits_instructionIndex;
  wire         sinkVec_validSink_11_valid;
  wire [4:0]   sinkVec_validSink_11_bits_vd;
  wire [1:0]   sinkVec_validSink_11_bits_offset;
  wire [3:0]   sinkVec_validSink_11_bits_mask;
  wire [31:0]  sinkVec_validSink_11_bits_data;
  wire         sinkVec_validSink_11_bits_last;
  wire [2:0]   sinkVec_validSink_11_bits_instructionIndex;
  assign sinkVec_sinkWire_11_valid = sinkVec_queue_11_deq_valid;
  assign sinkVec_sinkWire_11_bits_vd = sinkVec_queue_11_deq_bits_vd;
  assign sinkVec_sinkWire_11_bits_offset = sinkVec_queue_11_deq_bits_offset;
  assign sinkVec_sinkWire_11_bits_mask = sinkVec_queue_11_deq_bits_mask;
  assign sinkVec_sinkWire_11_bits_data = sinkVec_queue_11_deq_bits_data;
  assign sinkVec_sinkWire_11_bits_last = sinkVec_queue_11_deq_bits_last;
  assign sinkVec_sinkWire_11_bits_instructionIndex = sinkVec_queue_11_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_11_enq_bits_data;
  wire         sinkVec_queue_11_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_5 = {sinkVec_queue_11_enq_bits_data, sinkVec_queue_11_enq_bits_last};
  wire [2:0]   sinkVec_queue_11_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_11 = {sinkVec_queue_dataIn_lo_hi_5, sinkVec_queue_11_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_11_enq_bits_vd;
  wire [1:0]   sinkVec_queue_11_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_5 = {sinkVec_queue_11_enq_bits_vd, sinkVec_queue_11_enq_bits_offset};
  wire [3:0]   sinkVec_queue_11_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_11 = {sinkVec_queue_dataIn_hi_hi_5, sinkVec_queue_11_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_11 = {sinkVec_queue_dataIn_hi_11, sinkVec_queue_dataIn_lo_11};
  wire [2:0]   sinkVec_queue_dataOut_11_instructionIndex = _sinkVec_queue_fifo_11_data_out[2:0];
  wire         sinkVec_queue_dataOut_11_last = _sinkVec_queue_fifo_11_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_11_data = _sinkVec_queue_fifo_11_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_11_mask = _sinkVec_queue_fifo_11_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_11_offset = _sinkVec_queue_fifo_11_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_11_vd = _sinkVec_queue_fifo_11_data_out[46:42];
  wire         sinkVec_queue_11_enq_ready = ~_sinkVec_queue_fifo_11_full;
  wire         sinkVec_queue_11_enq_valid;
  assign sinkVec_queue_11_deq_valid = ~_sinkVec_queue_fifo_11_empty | sinkVec_queue_11_enq_valid;
  assign sinkVec_queue_11_deq_bits_vd = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_vd : sinkVec_queue_dataOut_11_vd;
  assign sinkVec_queue_11_deq_bits_offset = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_offset : sinkVec_queue_dataOut_11_offset;
  assign sinkVec_queue_11_deq_bits_mask = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_mask : sinkVec_queue_dataOut_11_mask;
  assign sinkVec_queue_11_deq_bits_data = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_data : sinkVec_queue_dataOut_11_data;
  assign sinkVec_queue_11_deq_bits_last = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_last : sinkVec_queue_dataOut_11_last;
  assign sinkVec_queue_11_deq_bits_instructionIndex = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_instructionIndex : sinkVec_queue_dataOut_11_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_11;
  wire         sinkVec_releasePipe_pipe_out_11_valid = sinkVec_releasePipe_pipe_v_11;
  wire         x22_2_1_ready;
  wire         x22_2_1_valid;
  wire         sinkVec_validSource_11_valid = x22_2_1_ready & x22_2_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_11;
  wire [2:0]   sinkVec_tokenCheck_counterChange_11 = sinkVec_validSource_11_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_11 = ~(sinkVec_tokenCheck_counter_11[2]);
  assign x22_2_1_ready = sinkVec_tokenCheck_11;
  assign sinkVec_queue_11_enq_valid = sinkVec_validSink_11_valid;
  assign sinkVec_queue_11_enq_bits_vd = sinkVec_validSink_11_bits_vd;
  assign sinkVec_queue_11_enq_bits_offset = sinkVec_validSink_11_bits_offset;
  assign sinkVec_queue_11_enq_bits_mask = sinkVec_validSink_11_bits_mask;
  assign sinkVec_queue_11_enq_bits_data = sinkVec_validSink_11_bits_data;
  assign sinkVec_queue_11_enq_bits_last = sinkVec_validSink_11_bits_last;
  assign sinkVec_queue_11_enq_bits_instructionIndex = sinkVec_validSink_11_bits_instructionIndex;
  reg          sinkVec_shifterReg_11_0_valid;
  assign sinkVec_validSink_11_valid = sinkVec_shifterReg_11_0_valid;
  reg  [4:0]   sinkVec_shifterReg_11_0_bits_vd;
  assign sinkVec_validSink_11_bits_vd = sinkVec_shifterReg_11_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_11_0_bits_offset;
  assign sinkVec_validSink_11_bits_offset = sinkVec_shifterReg_11_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_11_0_bits_mask;
  assign sinkVec_validSink_11_bits_mask = sinkVec_shifterReg_11_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_11_0_bits_data;
  assign sinkVec_validSink_11_bits_data = sinkVec_shifterReg_11_0_bits_data;
  reg          sinkVec_shifterReg_11_0_bits_last;
  assign sinkVec_validSink_11_bits_last = sinkVec_shifterReg_11_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_11_0_bits_instructionIndex;
  assign sinkVec_validSink_11_bits_instructionIndex = sinkVec_shifterReg_11_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_11 = sinkVec_shifterReg_11_0_valid | sinkVec_validSource_11_valid;
  assign sinkVec_sinkWire_10_ready = sinkVec_5_0_ready;
  assign sinkVec_sinkWire_11_ready = sinkVec_5_1_ready;
  reg          maskUnitFirst_5;
  wire         tryToRead_5 = sinkVec_5_0_valid | sinkVec_5_1_valid;
  wire         sinkWire_5_valid = maskUnitFirst_5 ? sinkVec_5_0_valid : sinkVec_5_1_valid;
  wire [4:0]   sinkWire_5_bits_vd = maskUnitFirst_5 ? sinkVec_5_0_bits_vd : sinkVec_5_1_bits_vd;
  wire [1:0]   sinkWire_5_bits_offset = maskUnitFirst_5 ? sinkVec_5_0_bits_offset : sinkVec_5_1_bits_offset;
  wire [3:0]   sinkWire_5_bits_mask = maskUnitFirst_5 ? sinkVec_5_0_bits_mask : sinkVec_5_1_bits_mask;
  wire [31:0]  sinkWire_5_bits_data = maskUnitFirst_5 ? sinkVec_5_0_bits_data : sinkVec_5_1_bits_data;
  wire         sinkWire_5_bits_last = maskUnitFirst_5 ? sinkVec_5_0_bits_last : sinkVec_5_1_bits_last;
  wire [2:0]   sinkWire_5_bits_instructionIndex = maskUnitFirst_5 ? sinkVec_5_0_bits_instructionIndex : sinkVec_5_1_bits_instructionIndex;
  wire         sinkWire_5_ready;
  assign sinkVec_5_1_ready = sinkWire_5_ready & ~maskUnitFirst_5;
  assign sinkVec_5_0_ready = sinkWire_5_ready & maskUnitFirst_5;
  reg          view__writeRelease_2_pipe_v;
  wire         view__writeRelease_2_pipe_out_valid = view__writeRelease_2_pipe_v;
  reg          pipe_v_6;
  wire         pipe_out_4_valid = pipe_v_6;
  wire         _probeWire_writeQueueEnqVec_2_valid_T = x22_2_0_ready & _maskUnit_exeResp_2_valid;
  reg          instructionFinishedPipe_pipe_v_2;
  wire         instructionFinishedPipe_pipe_out_2_valid = instructionFinishedPipe_pipe_v_2;
  reg  [7:0]   instructionFinishedPipe_pipe_b_2;
  wire [7:0]   instructionFinishedPipe_pipe_out_2_bits = instructionFinishedPipe_pipe_b_2;
  wire         instructionFinished_2_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_2_bits);
  assign vxsatReportVec_2 = _laneVec_2_vxsatReport[3:0];
  reg          pipe_v_7;
  reg  [31:0]  pipe_b_7;
  reg          pipe_pipe_v_2;
  wire         pipe_pipe_out_2_valid = pipe_pipe_v_2;
  reg  [31:0]  pipe_pipe_b_2;
  wire [31:0]  pipe_pipe_out_2_bits = pipe_pipe_b_2;
  reg          view__laneMaskSelect_2_pipe_v;
  reg  [5:0]   view__laneMaskSelect_2_pipe_b;
  reg          view__laneMaskSelect_2_pipe_pipe_v;
  wire         view__laneMaskSelect_2_pipe_pipe_out_valid = view__laneMaskSelect_2_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_2_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_2_pipe_pipe_out_bits = view__laneMaskSelect_2_pipe_pipe_b;
  reg          view__laneMaskSewSelect_2_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_2_pipe_b;
  reg          view__laneMaskSewSelect_2_pipe_pipe_v;
  wire         view__laneMaskSewSelect_2_pipe_pipe_out_valid = view__laneMaskSewSelect_2_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_2_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_2_pipe_pipe_out_bits = view__laneMaskSewSelect_2_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_2;
  wire         lsuLastPipe_pipe_out_2_valid = lsuLastPipe_pipe_v_2;
  reg  [7:0]   lsuLastPipe_pipe_b_2;
  wire [7:0]   lsuLastPipe_pipe_out_2_bits = lsuLastPipe_pipe_b_2;
  reg          maskLastPipe_pipe_v_2;
  wire         maskLastPipe_pipe_out_2_valid = maskLastPipe_pipe_v_2;
  reg  [7:0]   maskLastPipe_pipe_b_2;
  wire [7:0]   maskLastPipe_pipe_out_2_bits = maskLastPipe_pipe_b_2;
  wire [5:0]   writeCounter_2 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h8};
  reg          pipe_v_8;
  wire         pipe_out_5_valid = pipe_v_8;
  reg  [5:0]   pipe_b_8;
  wire [5:0]   pipe_out_5_bits = pipe_b_8;
  assign laneRequestSinkWire_3_ready = ~laneRequestSinkWire_3_bits_issueInst | _laneVec_3_laneRequest_ready;
  wire         sinkVec_tokenCheck_12;
  wire [4:0]   sinkVec_validSource_12_bits_vs = x13_3_0_bits_vs;
  wire [1:0]   sinkVec_validSource_12_bits_offset = x13_3_0_bits_offset;
  wire [2:0]   sinkVec_validSource_12_bits_instructionIndex = x13_3_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_13;
  wire [4:0]   sinkVec_validSource_13_bits_vs = x13_3_1_bits_vs;
  wire [1:0]   sinkVec_validSource_13_bits_offset = x13_3_1_bits_offset;
  wire [2:0]   sinkVec_validSource_13_bits_instructionIndex = x13_3_1_bits_instructionIndex;
  wire         sinkVec_6_0_ready;
  wire         sinkVec_queue_12_deq_ready = sinkVec_sinkWire_12_ready;
  wire         sinkVec_queue_12_deq_valid;
  wire [4:0]   sinkVec_queue_12_deq_bits_vs;
  wire         sinkVec_6_0_valid = sinkVec_sinkWire_12_valid;
  wire [1:0]   sinkVec_queue_12_deq_bits_readSource;
  wire [4:0]   sinkVec_6_0_bits_vs = sinkVec_sinkWire_12_bits_vs;
  wire [1:0]   sinkVec_queue_12_deq_bits_offset;
  wire [1:0]   sinkVec_6_0_bits_readSource = sinkVec_sinkWire_12_bits_readSource;
  wire [2:0]   sinkVec_queue_12_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_6_0_bits_offset = sinkVec_sinkWire_12_bits_offset;
  wire [2:0]   sinkVec_6_0_bits_instructionIndex = sinkVec_sinkWire_12_bits_instructionIndex;
  wire         sinkVec_validSink_12_valid;
  wire [4:0]   sinkVec_validSink_12_bits_vs;
  wire [1:0]   sinkVec_validSink_12_bits_readSource;
  wire [1:0]   sinkVec_validSink_12_bits_offset;
  wire [2:0]   sinkVec_validSink_12_bits_instructionIndex;
  assign sinkVec_sinkWire_12_valid = sinkVec_queue_12_deq_valid;
  assign sinkVec_sinkWire_12_bits_vs = sinkVec_queue_12_deq_bits_vs;
  assign sinkVec_sinkWire_12_bits_readSource = sinkVec_queue_12_deq_bits_readSource;
  assign sinkVec_sinkWire_12_bits_offset = sinkVec_queue_12_deq_bits_offset;
  assign sinkVec_sinkWire_12_bits_instructionIndex = sinkVec_queue_12_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_12_enq_bits_offset;
  wire [2:0]   sinkVec_queue_12_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_12 = {sinkVec_queue_12_enq_bits_offset, sinkVec_queue_12_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_12_enq_bits_vs;
  wire [1:0]   sinkVec_queue_12_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_12 = {sinkVec_queue_12_enq_bits_vs, sinkVec_queue_12_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_12 = {sinkVec_queue_dataIn_hi_12, sinkVec_queue_dataIn_lo_12};
  wire [2:0]   sinkVec_queue_dataOut_12_instructionIndex = _sinkVec_queue_fifo_12_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_12_offset = _sinkVec_queue_fifo_12_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_12_readSource = _sinkVec_queue_fifo_12_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_12_vs = _sinkVec_queue_fifo_12_data_out[11:7];
  wire         sinkVec_queue_12_enq_ready = ~_sinkVec_queue_fifo_12_full;
  wire         sinkVec_queue_12_enq_valid;
  assign sinkVec_queue_12_deq_valid = ~_sinkVec_queue_fifo_12_empty | sinkVec_queue_12_enq_valid;
  assign sinkVec_queue_12_deq_bits_vs = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_vs : sinkVec_queue_dataOut_12_vs;
  assign sinkVec_queue_12_deq_bits_readSource = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_readSource : sinkVec_queue_dataOut_12_readSource;
  assign sinkVec_queue_12_deq_bits_offset = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_offset : sinkVec_queue_dataOut_12_offset;
  assign sinkVec_queue_12_deq_bits_instructionIndex = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_instructionIndex : sinkVec_queue_dataOut_12_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_12;
  wire         sinkVec_releasePipe_pipe_out_12_valid = sinkVec_releasePipe_pipe_v_12;
  wire         x13_3_0_ready;
  wire         x13_3_0_valid;
  wire         sinkVec_validSource_12_valid = x13_3_0_ready & x13_3_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_12;
  wire [2:0]   sinkVec_tokenCheck_counterChange_12 = sinkVec_validSource_12_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_12 = ~(sinkVec_tokenCheck_counter_12[2]);
  assign x13_3_0_ready = sinkVec_tokenCheck_12;
  assign sinkVec_queue_12_enq_valid = sinkVec_validSink_12_valid;
  assign sinkVec_queue_12_enq_bits_vs = sinkVec_validSink_12_bits_vs;
  assign sinkVec_queue_12_enq_bits_readSource = sinkVec_validSink_12_bits_readSource;
  assign sinkVec_queue_12_enq_bits_offset = sinkVec_validSink_12_bits_offset;
  assign sinkVec_queue_12_enq_bits_instructionIndex = sinkVec_validSink_12_bits_instructionIndex;
  reg          sinkVec_shifterReg_12_0_valid;
  assign sinkVec_validSink_12_valid = sinkVec_shifterReg_12_0_valid;
  reg  [4:0]   sinkVec_shifterReg_12_0_bits_vs;
  assign sinkVec_validSink_12_bits_vs = sinkVec_shifterReg_12_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_12_0_bits_readSource;
  assign sinkVec_validSink_12_bits_readSource = sinkVec_shifterReg_12_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_12_0_bits_offset;
  assign sinkVec_validSink_12_bits_offset = sinkVec_shifterReg_12_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_12_0_bits_instructionIndex;
  assign sinkVec_validSink_12_bits_instructionIndex = sinkVec_shifterReg_12_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_12 = sinkVec_shifterReg_12_0_valid | sinkVec_validSource_12_valid;
  wire         sinkVec_6_1_ready;
  wire         sinkVec_queue_13_deq_ready = sinkVec_sinkWire_13_ready;
  wire         sinkVec_queue_13_deq_valid;
  wire [4:0]   sinkVec_queue_13_deq_bits_vs;
  wire         sinkVec_6_1_valid = sinkVec_sinkWire_13_valid;
  wire [1:0]   sinkVec_queue_13_deq_bits_readSource;
  wire [4:0]   sinkVec_6_1_bits_vs = sinkVec_sinkWire_13_bits_vs;
  wire [1:0]   sinkVec_queue_13_deq_bits_offset;
  wire [1:0]   sinkVec_6_1_bits_readSource = sinkVec_sinkWire_13_bits_readSource;
  wire [2:0]   sinkVec_queue_13_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_6_1_bits_offset = sinkVec_sinkWire_13_bits_offset;
  wire [2:0]   sinkVec_6_1_bits_instructionIndex = sinkVec_sinkWire_13_bits_instructionIndex;
  wire         sinkVec_validSink_13_valid;
  wire [4:0]   sinkVec_validSink_13_bits_vs;
  wire [1:0]   sinkVec_validSink_13_bits_readSource;
  wire [1:0]   sinkVec_validSink_13_bits_offset;
  wire [2:0]   sinkVec_validSink_13_bits_instructionIndex;
  assign sinkVec_sinkWire_13_valid = sinkVec_queue_13_deq_valid;
  assign sinkVec_sinkWire_13_bits_vs = sinkVec_queue_13_deq_bits_vs;
  assign sinkVec_sinkWire_13_bits_readSource = sinkVec_queue_13_deq_bits_readSource;
  assign sinkVec_sinkWire_13_bits_offset = sinkVec_queue_13_deq_bits_offset;
  assign sinkVec_sinkWire_13_bits_instructionIndex = sinkVec_queue_13_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_13_enq_bits_offset;
  wire [2:0]   sinkVec_queue_13_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_13 = {sinkVec_queue_13_enq_bits_offset, sinkVec_queue_13_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_13_enq_bits_vs;
  wire [1:0]   sinkVec_queue_13_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_13 = {sinkVec_queue_13_enq_bits_vs, sinkVec_queue_13_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_13 = {sinkVec_queue_dataIn_hi_13, sinkVec_queue_dataIn_lo_13};
  wire [2:0]   sinkVec_queue_dataOut_13_instructionIndex = _sinkVec_queue_fifo_13_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_13_offset = _sinkVec_queue_fifo_13_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_13_readSource = _sinkVec_queue_fifo_13_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_13_vs = _sinkVec_queue_fifo_13_data_out[11:7];
  wire         sinkVec_queue_13_enq_ready = ~_sinkVec_queue_fifo_13_full;
  wire         sinkVec_queue_13_enq_valid;
  assign sinkVec_queue_13_deq_valid = ~_sinkVec_queue_fifo_13_empty | sinkVec_queue_13_enq_valid;
  assign sinkVec_queue_13_deq_bits_vs = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_vs : sinkVec_queue_dataOut_13_vs;
  assign sinkVec_queue_13_deq_bits_readSource = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_readSource : sinkVec_queue_dataOut_13_readSource;
  assign sinkVec_queue_13_deq_bits_offset = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_offset : sinkVec_queue_dataOut_13_offset;
  assign sinkVec_queue_13_deq_bits_instructionIndex = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_instructionIndex : sinkVec_queue_dataOut_13_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_13;
  wire         sinkVec_releasePipe_pipe_out_13_valid = sinkVec_releasePipe_pipe_v_13;
  wire         x13_3_1_ready;
  wire         x13_3_1_valid;
  wire         sinkVec_validSource_13_valid = x13_3_1_ready & x13_3_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_13;
  wire [2:0]   sinkVec_tokenCheck_counterChange_13 = sinkVec_validSource_13_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_13 = ~(sinkVec_tokenCheck_counter_13[2]);
  assign x13_3_1_ready = sinkVec_tokenCheck_13;
  assign sinkVec_queue_13_enq_valid = sinkVec_validSink_13_valid;
  assign sinkVec_queue_13_enq_bits_vs = sinkVec_validSink_13_bits_vs;
  assign sinkVec_queue_13_enq_bits_readSource = sinkVec_validSink_13_bits_readSource;
  assign sinkVec_queue_13_enq_bits_offset = sinkVec_validSink_13_bits_offset;
  assign sinkVec_queue_13_enq_bits_instructionIndex = sinkVec_validSink_13_bits_instructionIndex;
  reg          sinkVec_shifterReg_13_0_valid;
  assign sinkVec_validSink_13_valid = sinkVec_shifterReg_13_0_valid;
  reg  [4:0]   sinkVec_shifterReg_13_0_bits_vs;
  assign sinkVec_validSink_13_bits_vs = sinkVec_shifterReg_13_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_13_0_bits_readSource;
  assign sinkVec_validSink_13_bits_readSource = sinkVec_shifterReg_13_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_13_0_bits_offset;
  assign sinkVec_validSink_13_bits_offset = sinkVec_shifterReg_13_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_13_0_bits_instructionIndex;
  assign sinkVec_validSink_13_bits_instructionIndex = sinkVec_shifterReg_13_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_13 = sinkVec_shifterReg_13_0_valid | sinkVec_validSource_13_valid;
  assign sinkVec_sinkWire_12_ready = sinkVec_6_0_ready;
  assign sinkVec_sinkWire_13_ready = sinkVec_6_1_ready;
  reg          maskUnitFirst_6;
  wire         tryToRead_6 = sinkVec_6_0_valid | sinkVec_6_1_valid;
  wire         sinkWire_6_valid = maskUnitFirst_6 ? sinkVec_6_0_valid : sinkVec_6_1_valid;
  wire [4:0]   sinkWire_6_bits_vs = maskUnitFirst_6 ? sinkVec_6_0_bits_vs : sinkVec_6_1_bits_vs;
  wire [1:0]   sinkWire_6_bits_readSource = maskUnitFirst_6 ? sinkVec_6_0_bits_readSource : sinkVec_6_1_bits_readSource;
  wire [1:0]   sinkWire_6_bits_offset = maskUnitFirst_6 ? sinkVec_6_0_bits_offset : sinkVec_6_1_bits_offset;
  wire [2:0]   sinkWire_6_bits_instructionIndex = maskUnitFirst_6 ? sinkVec_6_0_bits_instructionIndex : sinkVec_6_1_bits_instructionIndex;
  wire         sinkWire_6_ready;
  assign sinkVec_6_1_ready = sinkWire_6_ready & ~maskUnitFirst_6;
  assign sinkVec_6_0_ready = sinkWire_6_ready & maskUnitFirst_6;
  reg          accessDataValid_pipe_v_6;
  reg          accessDataValid_pipe_pipe_v_6;
  wire         accessDataValid_pipe_pipe_out_6_valid = accessDataValid_pipe_pipe_v_6;
  wire         accessDataSource_6_valid = accessDataValid_pipe_pipe_out_6_valid;
  reg          shifterReg_22_0_valid;
  reg  [31:0]  shifterReg_22_0_bits;
  wire         shifterValid_22 = shifterReg_22_0_valid | accessDataSource_6_valid;
  reg          accessDataValid_pipe_v_7;
  reg          accessDataValid_pipe_pipe_v_7;
  wire         accessDataValid_pipe_pipe_out_7_valid = accessDataValid_pipe_pipe_v_7;
  wire         accessDataSource_7_valid = accessDataValid_pipe_pipe_out_7_valid;
  reg          shifterReg_23_0_valid;
  reg  [31:0]  shifterReg_23_0_bits;
  wire         shifterValid_23 = shifterReg_23_0_valid | accessDataSource_7_valid;
  wire         sinkVec_tokenCheck_14;
  wire [4:0]   sinkVec_validSource_14_bits_vd = x22_3_0_bits_vd;
  wire [1:0]   sinkVec_validSource_14_bits_offset = x22_3_0_bits_offset;
  wire [3:0]   sinkVec_validSource_14_bits_mask = x22_3_0_bits_mask;
  wire [31:0]  sinkVec_validSource_14_bits_data = x22_3_0_bits_data;
  wire [2:0]   sinkVec_validSource_14_bits_instructionIndex = x22_3_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_15;
  wire [4:0]   sinkVec_validSource_15_bits_vd = x22_3_1_bits_vd;
  wire [1:0]   sinkVec_validSource_15_bits_offset = x22_3_1_bits_offset;
  wire [3:0]   sinkVec_validSource_15_bits_mask = x22_3_1_bits_mask;
  wire [31:0]  sinkVec_validSource_15_bits_data = x22_3_1_bits_data;
  wire         sinkVec_validSource_15_bits_last = x22_3_1_bits_last;
  wire [2:0]   sinkVec_validSource_15_bits_instructionIndex = x22_3_1_bits_instructionIndex;
  wire         sinkVec_7_0_ready;
  wire         sinkVec_queue_14_deq_ready = sinkVec_sinkWire_14_ready;
  wire         sinkVec_queue_14_deq_valid;
  wire [4:0]   sinkVec_queue_14_deq_bits_vd;
  wire         sinkVec_7_0_valid = sinkVec_sinkWire_14_valid;
  wire [1:0]   sinkVec_queue_14_deq_bits_offset;
  wire [4:0]   sinkVec_7_0_bits_vd = sinkVec_sinkWire_14_bits_vd;
  wire [3:0]   sinkVec_queue_14_deq_bits_mask;
  wire [1:0]   sinkVec_7_0_bits_offset = sinkVec_sinkWire_14_bits_offset;
  wire [31:0]  sinkVec_queue_14_deq_bits_data;
  wire [3:0]   sinkVec_7_0_bits_mask = sinkVec_sinkWire_14_bits_mask;
  wire         sinkVec_queue_14_deq_bits_last;
  wire [31:0]  sinkVec_7_0_bits_data = sinkVec_sinkWire_14_bits_data;
  wire [2:0]   sinkVec_queue_14_deq_bits_instructionIndex;
  wire         sinkVec_7_0_bits_last = sinkVec_sinkWire_14_bits_last;
  wire [2:0]   sinkVec_7_0_bits_instructionIndex = sinkVec_sinkWire_14_bits_instructionIndex;
  wire         sinkVec_validSink_14_valid;
  wire [4:0]   sinkVec_validSink_14_bits_vd;
  wire [1:0]   sinkVec_validSink_14_bits_offset;
  wire [3:0]   sinkVec_validSink_14_bits_mask;
  wire [31:0]  sinkVec_validSink_14_bits_data;
  wire [2:0]   sinkVec_validSink_14_bits_instructionIndex;
  assign sinkVec_sinkWire_14_valid = sinkVec_queue_14_deq_valid;
  assign sinkVec_sinkWire_14_bits_vd = sinkVec_queue_14_deq_bits_vd;
  assign sinkVec_sinkWire_14_bits_offset = sinkVec_queue_14_deq_bits_offset;
  assign sinkVec_sinkWire_14_bits_mask = sinkVec_queue_14_deq_bits_mask;
  assign sinkVec_sinkWire_14_bits_data = sinkVec_queue_14_deq_bits_data;
  assign sinkVec_sinkWire_14_bits_last = sinkVec_queue_14_deq_bits_last;
  assign sinkVec_sinkWire_14_bits_instructionIndex = sinkVec_queue_14_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_14_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_6 = {sinkVec_queue_14_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_14_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_14 = {sinkVec_queue_dataIn_lo_hi_6, sinkVec_queue_14_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_14_enq_bits_vd;
  wire [1:0]   sinkVec_queue_14_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_6 = {sinkVec_queue_14_enq_bits_vd, sinkVec_queue_14_enq_bits_offset};
  wire [3:0]   sinkVec_queue_14_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_14 = {sinkVec_queue_dataIn_hi_hi_6, sinkVec_queue_14_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_14 = {sinkVec_queue_dataIn_hi_14, sinkVec_queue_dataIn_lo_14};
  wire [2:0]   sinkVec_queue_dataOut_14_instructionIndex = _sinkVec_queue_fifo_14_data_out[2:0];
  wire         sinkVec_queue_dataOut_14_last = _sinkVec_queue_fifo_14_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_14_data = _sinkVec_queue_fifo_14_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_14_mask = _sinkVec_queue_fifo_14_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_14_offset = _sinkVec_queue_fifo_14_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_14_vd = _sinkVec_queue_fifo_14_data_out[46:42];
  wire         sinkVec_queue_14_enq_ready = ~_sinkVec_queue_fifo_14_full;
  wire         sinkVec_queue_14_enq_valid;
  assign sinkVec_queue_14_deq_valid = ~_sinkVec_queue_fifo_14_empty | sinkVec_queue_14_enq_valid;
  assign sinkVec_queue_14_deq_bits_vd = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_vd : sinkVec_queue_dataOut_14_vd;
  assign sinkVec_queue_14_deq_bits_offset = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_offset : sinkVec_queue_dataOut_14_offset;
  assign sinkVec_queue_14_deq_bits_mask = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_mask : sinkVec_queue_dataOut_14_mask;
  assign sinkVec_queue_14_deq_bits_data = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_data : sinkVec_queue_dataOut_14_data;
  assign sinkVec_queue_14_deq_bits_last = ~_sinkVec_queue_fifo_14_empty & sinkVec_queue_dataOut_14_last;
  assign sinkVec_queue_14_deq_bits_instructionIndex = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_instructionIndex : sinkVec_queue_dataOut_14_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_14;
  wire         sinkVec_releasePipe_pipe_out_14_valid = sinkVec_releasePipe_pipe_v_14;
  wire         x22_3_0_ready;
  wire         x22_3_0_valid;
  wire         sinkVec_validSource_14_valid = x22_3_0_ready & x22_3_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_14;
  wire [2:0]   sinkVec_tokenCheck_counterChange_14 = sinkVec_validSource_14_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_14 = ~(sinkVec_tokenCheck_counter_14[2]);
  assign x22_3_0_ready = sinkVec_tokenCheck_14;
  assign sinkVec_queue_14_enq_valid = sinkVec_validSink_14_valid;
  assign sinkVec_queue_14_enq_bits_vd = sinkVec_validSink_14_bits_vd;
  assign sinkVec_queue_14_enq_bits_offset = sinkVec_validSink_14_bits_offset;
  assign sinkVec_queue_14_enq_bits_mask = sinkVec_validSink_14_bits_mask;
  assign sinkVec_queue_14_enq_bits_data = sinkVec_validSink_14_bits_data;
  assign sinkVec_queue_14_enq_bits_instructionIndex = sinkVec_validSink_14_bits_instructionIndex;
  reg          sinkVec_shifterReg_14_0_valid;
  assign sinkVec_validSink_14_valid = sinkVec_shifterReg_14_0_valid;
  reg  [4:0]   sinkVec_shifterReg_14_0_bits_vd;
  assign sinkVec_validSink_14_bits_vd = sinkVec_shifterReg_14_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_14_0_bits_offset;
  assign sinkVec_validSink_14_bits_offset = sinkVec_shifterReg_14_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_14_0_bits_mask;
  assign sinkVec_validSink_14_bits_mask = sinkVec_shifterReg_14_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_14_0_bits_data;
  assign sinkVec_validSink_14_bits_data = sinkVec_shifterReg_14_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_14_0_bits_instructionIndex;
  assign sinkVec_validSink_14_bits_instructionIndex = sinkVec_shifterReg_14_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_14 = sinkVec_shifterReg_14_0_valid | sinkVec_validSource_14_valid;
  wire         sinkVec_7_1_ready;
  wire         sinkVec_queue_15_deq_ready = sinkVec_sinkWire_15_ready;
  wire         sinkVec_queue_15_deq_valid;
  wire [4:0]   sinkVec_queue_15_deq_bits_vd;
  wire         sinkVec_7_1_valid = sinkVec_sinkWire_15_valid;
  wire [1:0]   sinkVec_queue_15_deq_bits_offset;
  wire [4:0]   sinkVec_7_1_bits_vd = sinkVec_sinkWire_15_bits_vd;
  wire [3:0]   sinkVec_queue_15_deq_bits_mask;
  wire [1:0]   sinkVec_7_1_bits_offset = sinkVec_sinkWire_15_bits_offset;
  wire [31:0]  sinkVec_queue_15_deq_bits_data;
  wire [3:0]   sinkVec_7_1_bits_mask = sinkVec_sinkWire_15_bits_mask;
  wire         sinkVec_queue_15_deq_bits_last;
  wire [31:0]  sinkVec_7_1_bits_data = sinkVec_sinkWire_15_bits_data;
  wire [2:0]   sinkVec_queue_15_deq_bits_instructionIndex;
  wire         sinkVec_7_1_bits_last = sinkVec_sinkWire_15_bits_last;
  wire [2:0]   sinkVec_7_1_bits_instructionIndex = sinkVec_sinkWire_15_bits_instructionIndex;
  wire         sinkVec_validSink_15_valid;
  wire [4:0]   sinkVec_validSink_15_bits_vd;
  wire [1:0]   sinkVec_validSink_15_bits_offset;
  wire [3:0]   sinkVec_validSink_15_bits_mask;
  wire [31:0]  sinkVec_validSink_15_bits_data;
  wire         sinkVec_validSink_15_bits_last;
  wire [2:0]   sinkVec_validSink_15_bits_instructionIndex;
  assign sinkVec_sinkWire_15_valid = sinkVec_queue_15_deq_valid;
  assign sinkVec_sinkWire_15_bits_vd = sinkVec_queue_15_deq_bits_vd;
  assign sinkVec_sinkWire_15_bits_offset = sinkVec_queue_15_deq_bits_offset;
  assign sinkVec_sinkWire_15_bits_mask = sinkVec_queue_15_deq_bits_mask;
  assign sinkVec_sinkWire_15_bits_data = sinkVec_queue_15_deq_bits_data;
  assign sinkVec_sinkWire_15_bits_last = sinkVec_queue_15_deq_bits_last;
  assign sinkVec_sinkWire_15_bits_instructionIndex = sinkVec_queue_15_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_15_enq_bits_data;
  wire         sinkVec_queue_15_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_7 = {sinkVec_queue_15_enq_bits_data, sinkVec_queue_15_enq_bits_last};
  wire [2:0]   sinkVec_queue_15_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_15 = {sinkVec_queue_dataIn_lo_hi_7, sinkVec_queue_15_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_15_enq_bits_vd;
  wire [1:0]   sinkVec_queue_15_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_7 = {sinkVec_queue_15_enq_bits_vd, sinkVec_queue_15_enq_bits_offset};
  wire [3:0]   sinkVec_queue_15_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_15 = {sinkVec_queue_dataIn_hi_hi_7, sinkVec_queue_15_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_15 = {sinkVec_queue_dataIn_hi_15, sinkVec_queue_dataIn_lo_15};
  wire [2:0]   sinkVec_queue_dataOut_15_instructionIndex = _sinkVec_queue_fifo_15_data_out[2:0];
  wire         sinkVec_queue_dataOut_15_last = _sinkVec_queue_fifo_15_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_15_data = _sinkVec_queue_fifo_15_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_15_mask = _sinkVec_queue_fifo_15_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_15_offset = _sinkVec_queue_fifo_15_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_15_vd = _sinkVec_queue_fifo_15_data_out[46:42];
  wire         sinkVec_queue_15_enq_ready = ~_sinkVec_queue_fifo_15_full;
  wire         sinkVec_queue_15_enq_valid;
  assign sinkVec_queue_15_deq_valid = ~_sinkVec_queue_fifo_15_empty | sinkVec_queue_15_enq_valid;
  assign sinkVec_queue_15_deq_bits_vd = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_vd : sinkVec_queue_dataOut_15_vd;
  assign sinkVec_queue_15_deq_bits_offset = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_offset : sinkVec_queue_dataOut_15_offset;
  assign sinkVec_queue_15_deq_bits_mask = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_mask : sinkVec_queue_dataOut_15_mask;
  assign sinkVec_queue_15_deq_bits_data = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_data : sinkVec_queue_dataOut_15_data;
  assign sinkVec_queue_15_deq_bits_last = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_last : sinkVec_queue_dataOut_15_last;
  assign sinkVec_queue_15_deq_bits_instructionIndex = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_instructionIndex : sinkVec_queue_dataOut_15_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_15;
  wire         sinkVec_releasePipe_pipe_out_15_valid = sinkVec_releasePipe_pipe_v_15;
  wire         x22_3_1_ready;
  wire         x22_3_1_valid;
  wire         sinkVec_validSource_15_valid = x22_3_1_ready & x22_3_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_15;
  wire [2:0]   sinkVec_tokenCheck_counterChange_15 = sinkVec_validSource_15_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_15 = ~(sinkVec_tokenCheck_counter_15[2]);
  assign x22_3_1_ready = sinkVec_tokenCheck_15;
  assign sinkVec_queue_15_enq_valid = sinkVec_validSink_15_valid;
  assign sinkVec_queue_15_enq_bits_vd = sinkVec_validSink_15_bits_vd;
  assign sinkVec_queue_15_enq_bits_offset = sinkVec_validSink_15_bits_offset;
  assign sinkVec_queue_15_enq_bits_mask = sinkVec_validSink_15_bits_mask;
  assign sinkVec_queue_15_enq_bits_data = sinkVec_validSink_15_bits_data;
  assign sinkVec_queue_15_enq_bits_last = sinkVec_validSink_15_bits_last;
  assign sinkVec_queue_15_enq_bits_instructionIndex = sinkVec_validSink_15_bits_instructionIndex;
  reg          sinkVec_shifterReg_15_0_valid;
  assign sinkVec_validSink_15_valid = sinkVec_shifterReg_15_0_valid;
  reg  [4:0]   sinkVec_shifterReg_15_0_bits_vd;
  assign sinkVec_validSink_15_bits_vd = sinkVec_shifterReg_15_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_15_0_bits_offset;
  assign sinkVec_validSink_15_bits_offset = sinkVec_shifterReg_15_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_15_0_bits_mask;
  assign sinkVec_validSink_15_bits_mask = sinkVec_shifterReg_15_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_15_0_bits_data;
  assign sinkVec_validSink_15_bits_data = sinkVec_shifterReg_15_0_bits_data;
  reg          sinkVec_shifterReg_15_0_bits_last;
  assign sinkVec_validSink_15_bits_last = sinkVec_shifterReg_15_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_15_0_bits_instructionIndex;
  assign sinkVec_validSink_15_bits_instructionIndex = sinkVec_shifterReg_15_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_15 = sinkVec_shifterReg_15_0_valid | sinkVec_validSource_15_valid;
  assign sinkVec_sinkWire_14_ready = sinkVec_7_0_ready;
  assign sinkVec_sinkWire_15_ready = sinkVec_7_1_ready;
  reg          maskUnitFirst_7;
  wire         tryToRead_7 = sinkVec_7_0_valid | sinkVec_7_1_valid;
  wire         sinkWire_7_valid = maskUnitFirst_7 ? sinkVec_7_0_valid : sinkVec_7_1_valid;
  wire [4:0]   sinkWire_7_bits_vd = maskUnitFirst_7 ? sinkVec_7_0_bits_vd : sinkVec_7_1_bits_vd;
  wire [1:0]   sinkWire_7_bits_offset = maskUnitFirst_7 ? sinkVec_7_0_bits_offset : sinkVec_7_1_bits_offset;
  wire [3:0]   sinkWire_7_bits_mask = maskUnitFirst_7 ? sinkVec_7_0_bits_mask : sinkVec_7_1_bits_mask;
  wire [31:0]  sinkWire_7_bits_data = maskUnitFirst_7 ? sinkVec_7_0_bits_data : sinkVec_7_1_bits_data;
  wire         sinkWire_7_bits_last = maskUnitFirst_7 ? sinkVec_7_0_bits_last : sinkVec_7_1_bits_last;
  wire [2:0]   sinkWire_7_bits_instructionIndex = maskUnitFirst_7 ? sinkVec_7_0_bits_instructionIndex : sinkVec_7_1_bits_instructionIndex;
  wire         sinkWire_7_ready;
  assign sinkVec_7_1_ready = sinkWire_7_ready & ~maskUnitFirst_7;
  assign sinkVec_7_0_ready = sinkWire_7_ready & maskUnitFirst_7;
  reg          view__writeRelease_3_pipe_v;
  wire         view__writeRelease_3_pipe_out_valid = view__writeRelease_3_pipe_v;
  reg          pipe_v_9;
  wire         pipe_out_6_valid = pipe_v_9;
  wire         _probeWire_writeQueueEnqVec_3_valid_T = x22_3_0_ready & _maskUnit_exeResp_3_valid;
  reg          instructionFinishedPipe_pipe_v_3;
  wire         instructionFinishedPipe_pipe_out_3_valid = instructionFinishedPipe_pipe_v_3;
  reg  [7:0]   instructionFinishedPipe_pipe_b_3;
  wire [7:0]   instructionFinishedPipe_pipe_out_3_bits = instructionFinishedPipe_pipe_b_3;
  wire         instructionFinished_3_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_3_bits);
  assign vxsatReportVec_3 = _laneVec_3_vxsatReport[3:0];
  reg          pipe_v_10;
  reg  [31:0]  pipe_b_10;
  reg          pipe_pipe_v_3;
  wire         pipe_pipe_out_3_valid = pipe_pipe_v_3;
  reg  [31:0]  pipe_pipe_b_3;
  wire [31:0]  pipe_pipe_out_3_bits = pipe_pipe_b_3;
  reg          view__laneMaskSelect_3_pipe_v;
  reg  [5:0]   view__laneMaskSelect_3_pipe_b;
  reg          view__laneMaskSelect_3_pipe_pipe_v;
  wire         view__laneMaskSelect_3_pipe_pipe_out_valid = view__laneMaskSelect_3_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_3_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_3_pipe_pipe_out_bits = view__laneMaskSelect_3_pipe_pipe_b;
  reg          view__laneMaskSewSelect_3_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_3_pipe_b;
  reg          view__laneMaskSewSelect_3_pipe_pipe_v;
  wire         view__laneMaskSewSelect_3_pipe_pipe_out_valid = view__laneMaskSewSelect_3_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_3_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_3_pipe_pipe_out_bits = view__laneMaskSewSelect_3_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_3;
  wire         lsuLastPipe_pipe_out_3_valid = lsuLastPipe_pipe_v_3;
  reg  [7:0]   lsuLastPipe_pipe_b_3;
  wire [7:0]   lsuLastPipe_pipe_out_3_bits = lsuLastPipe_pipe_b_3;
  reg          maskLastPipe_pipe_v_3;
  wire         maskLastPipe_pipe_out_3_valid = maskLastPipe_pipe_v_3;
  reg  [7:0]   maskLastPipe_pipe_b_3;
  wire [7:0]   maskLastPipe_pipe_out_3_bits = maskLastPipe_pipe_b_3;
  wire [5:0]   writeCounter_3 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'hC};
  reg          pipe_v_11;
  wire         pipe_out_7_valid = pipe_v_11;
  reg  [5:0]   pipe_b_11;
  wire [5:0]   pipe_out_7_bits = pipe_b_11;
  assign laneRequestSinkWire_4_ready = ~laneRequestSinkWire_4_bits_issueInst | _laneVec_4_laneRequest_ready;
  wire         sinkVec_tokenCheck_16;
  wire [4:0]   sinkVec_validSource_16_bits_vs = x13_4_0_bits_vs;
  wire [1:0]   sinkVec_validSource_16_bits_offset = x13_4_0_bits_offset;
  wire [2:0]   sinkVec_validSource_16_bits_instructionIndex = x13_4_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_17;
  wire [4:0]   sinkVec_validSource_17_bits_vs = x13_4_1_bits_vs;
  wire [1:0]   sinkVec_validSource_17_bits_offset = x13_4_1_bits_offset;
  wire [2:0]   sinkVec_validSource_17_bits_instructionIndex = x13_4_1_bits_instructionIndex;
  wire         sinkVec_8_0_ready;
  wire         sinkVec_queue_16_deq_ready = sinkVec_sinkWire_16_ready;
  wire         sinkVec_queue_16_deq_valid;
  wire [4:0]   sinkVec_queue_16_deq_bits_vs;
  wire         sinkVec_8_0_valid = sinkVec_sinkWire_16_valid;
  wire [1:0]   sinkVec_queue_16_deq_bits_readSource;
  wire [4:0]   sinkVec_8_0_bits_vs = sinkVec_sinkWire_16_bits_vs;
  wire [1:0]   sinkVec_queue_16_deq_bits_offset;
  wire [1:0]   sinkVec_8_0_bits_readSource = sinkVec_sinkWire_16_bits_readSource;
  wire [2:0]   sinkVec_queue_16_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_8_0_bits_offset = sinkVec_sinkWire_16_bits_offset;
  wire [2:0]   sinkVec_8_0_bits_instructionIndex = sinkVec_sinkWire_16_bits_instructionIndex;
  wire         sinkVec_validSink_16_valid;
  wire [4:0]   sinkVec_validSink_16_bits_vs;
  wire [1:0]   sinkVec_validSink_16_bits_readSource;
  wire [1:0]   sinkVec_validSink_16_bits_offset;
  wire [2:0]   sinkVec_validSink_16_bits_instructionIndex;
  assign sinkVec_sinkWire_16_valid = sinkVec_queue_16_deq_valid;
  assign sinkVec_sinkWire_16_bits_vs = sinkVec_queue_16_deq_bits_vs;
  assign sinkVec_sinkWire_16_bits_readSource = sinkVec_queue_16_deq_bits_readSource;
  assign sinkVec_sinkWire_16_bits_offset = sinkVec_queue_16_deq_bits_offset;
  assign sinkVec_sinkWire_16_bits_instructionIndex = sinkVec_queue_16_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_16_enq_bits_offset;
  wire [2:0]   sinkVec_queue_16_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_16 = {sinkVec_queue_16_enq_bits_offset, sinkVec_queue_16_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_16_enq_bits_vs;
  wire [1:0]   sinkVec_queue_16_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_16 = {sinkVec_queue_16_enq_bits_vs, sinkVec_queue_16_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_16 = {sinkVec_queue_dataIn_hi_16, sinkVec_queue_dataIn_lo_16};
  wire [2:0]   sinkVec_queue_dataOut_16_instructionIndex = _sinkVec_queue_fifo_16_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_16_offset = _sinkVec_queue_fifo_16_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_16_readSource = _sinkVec_queue_fifo_16_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_16_vs = _sinkVec_queue_fifo_16_data_out[11:7];
  wire         sinkVec_queue_16_enq_ready = ~_sinkVec_queue_fifo_16_full;
  wire         sinkVec_queue_16_enq_valid;
  assign sinkVec_queue_16_deq_valid = ~_sinkVec_queue_fifo_16_empty | sinkVec_queue_16_enq_valid;
  assign sinkVec_queue_16_deq_bits_vs = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_vs : sinkVec_queue_dataOut_16_vs;
  assign sinkVec_queue_16_deq_bits_readSource = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_readSource : sinkVec_queue_dataOut_16_readSource;
  assign sinkVec_queue_16_deq_bits_offset = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_offset : sinkVec_queue_dataOut_16_offset;
  assign sinkVec_queue_16_deq_bits_instructionIndex = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_instructionIndex : sinkVec_queue_dataOut_16_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_16;
  wire         sinkVec_releasePipe_pipe_out_16_valid = sinkVec_releasePipe_pipe_v_16;
  wire         x13_4_0_ready;
  wire         x13_4_0_valid;
  wire         sinkVec_validSource_16_valid = x13_4_0_ready & x13_4_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_16;
  wire [2:0]   sinkVec_tokenCheck_counterChange_16 = sinkVec_validSource_16_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_16 = ~(sinkVec_tokenCheck_counter_16[2]);
  assign x13_4_0_ready = sinkVec_tokenCheck_16;
  assign sinkVec_queue_16_enq_valid = sinkVec_validSink_16_valid;
  assign sinkVec_queue_16_enq_bits_vs = sinkVec_validSink_16_bits_vs;
  assign sinkVec_queue_16_enq_bits_readSource = sinkVec_validSink_16_bits_readSource;
  assign sinkVec_queue_16_enq_bits_offset = sinkVec_validSink_16_bits_offset;
  assign sinkVec_queue_16_enq_bits_instructionIndex = sinkVec_validSink_16_bits_instructionIndex;
  reg          sinkVec_shifterReg_16_0_valid;
  assign sinkVec_validSink_16_valid = sinkVec_shifterReg_16_0_valid;
  reg  [4:0]   sinkVec_shifterReg_16_0_bits_vs;
  assign sinkVec_validSink_16_bits_vs = sinkVec_shifterReg_16_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_16_0_bits_readSource;
  assign sinkVec_validSink_16_bits_readSource = sinkVec_shifterReg_16_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_16_0_bits_offset;
  assign sinkVec_validSink_16_bits_offset = sinkVec_shifterReg_16_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_16_0_bits_instructionIndex;
  assign sinkVec_validSink_16_bits_instructionIndex = sinkVec_shifterReg_16_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_16 = sinkVec_shifterReg_16_0_valid | sinkVec_validSource_16_valid;
  wire         sinkVec_8_1_ready;
  wire         sinkVec_queue_17_deq_ready = sinkVec_sinkWire_17_ready;
  wire         sinkVec_queue_17_deq_valid;
  wire [4:0]   sinkVec_queue_17_deq_bits_vs;
  wire         sinkVec_8_1_valid = sinkVec_sinkWire_17_valid;
  wire [1:0]   sinkVec_queue_17_deq_bits_readSource;
  wire [4:0]   sinkVec_8_1_bits_vs = sinkVec_sinkWire_17_bits_vs;
  wire [1:0]   sinkVec_queue_17_deq_bits_offset;
  wire [1:0]   sinkVec_8_1_bits_readSource = sinkVec_sinkWire_17_bits_readSource;
  wire [2:0]   sinkVec_queue_17_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_8_1_bits_offset = sinkVec_sinkWire_17_bits_offset;
  wire [2:0]   sinkVec_8_1_bits_instructionIndex = sinkVec_sinkWire_17_bits_instructionIndex;
  wire         sinkVec_validSink_17_valid;
  wire [4:0]   sinkVec_validSink_17_bits_vs;
  wire [1:0]   sinkVec_validSink_17_bits_readSource;
  wire [1:0]   sinkVec_validSink_17_bits_offset;
  wire [2:0]   sinkVec_validSink_17_bits_instructionIndex;
  assign sinkVec_sinkWire_17_valid = sinkVec_queue_17_deq_valid;
  assign sinkVec_sinkWire_17_bits_vs = sinkVec_queue_17_deq_bits_vs;
  assign sinkVec_sinkWire_17_bits_readSource = sinkVec_queue_17_deq_bits_readSource;
  assign sinkVec_sinkWire_17_bits_offset = sinkVec_queue_17_deq_bits_offset;
  assign sinkVec_sinkWire_17_bits_instructionIndex = sinkVec_queue_17_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_17_enq_bits_offset;
  wire [2:0]   sinkVec_queue_17_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_17 = {sinkVec_queue_17_enq_bits_offset, sinkVec_queue_17_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_17_enq_bits_vs;
  wire [1:0]   sinkVec_queue_17_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_17 = {sinkVec_queue_17_enq_bits_vs, sinkVec_queue_17_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_17 = {sinkVec_queue_dataIn_hi_17, sinkVec_queue_dataIn_lo_17};
  wire [2:0]   sinkVec_queue_dataOut_17_instructionIndex = _sinkVec_queue_fifo_17_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_17_offset = _sinkVec_queue_fifo_17_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_17_readSource = _sinkVec_queue_fifo_17_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_17_vs = _sinkVec_queue_fifo_17_data_out[11:7];
  wire         sinkVec_queue_17_enq_ready = ~_sinkVec_queue_fifo_17_full;
  wire         sinkVec_queue_17_enq_valid;
  assign sinkVec_queue_17_deq_valid = ~_sinkVec_queue_fifo_17_empty | sinkVec_queue_17_enq_valid;
  assign sinkVec_queue_17_deq_bits_vs = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_vs : sinkVec_queue_dataOut_17_vs;
  assign sinkVec_queue_17_deq_bits_readSource = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_readSource : sinkVec_queue_dataOut_17_readSource;
  assign sinkVec_queue_17_deq_bits_offset = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_offset : sinkVec_queue_dataOut_17_offset;
  assign sinkVec_queue_17_deq_bits_instructionIndex = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_instructionIndex : sinkVec_queue_dataOut_17_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_17;
  wire         sinkVec_releasePipe_pipe_out_17_valid = sinkVec_releasePipe_pipe_v_17;
  wire         x13_4_1_ready;
  wire         x13_4_1_valid;
  wire         sinkVec_validSource_17_valid = x13_4_1_ready & x13_4_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_17;
  wire [2:0]   sinkVec_tokenCheck_counterChange_17 = sinkVec_validSource_17_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_17 = ~(sinkVec_tokenCheck_counter_17[2]);
  assign x13_4_1_ready = sinkVec_tokenCheck_17;
  assign sinkVec_queue_17_enq_valid = sinkVec_validSink_17_valid;
  assign sinkVec_queue_17_enq_bits_vs = sinkVec_validSink_17_bits_vs;
  assign sinkVec_queue_17_enq_bits_readSource = sinkVec_validSink_17_bits_readSource;
  assign sinkVec_queue_17_enq_bits_offset = sinkVec_validSink_17_bits_offset;
  assign sinkVec_queue_17_enq_bits_instructionIndex = sinkVec_validSink_17_bits_instructionIndex;
  reg          sinkVec_shifterReg_17_0_valid;
  assign sinkVec_validSink_17_valid = sinkVec_shifterReg_17_0_valid;
  reg  [4:0]   sinkVec_shifterReg_17_0_bits_vs;
  assign sinkVec_validSink_17_bits_vs = sinkVec_shifterReg_17_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_17_0_bits_readSource;
  assign sinkVec_validSink_17_bits_readSource = sinkVec_shifterReg_17_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_17_0_bits_offset;
  assign sinkVec_validSink_17_bits_offset = sinkVec_shifterReg_17_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_17_0_bits_instructionIndex;
  assign sinkVec_validSink_17_bits_instructionIndex = sinkVec_shifterReg_17_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_17 = sinkVec_shifterReg_17_0_valid | sinkVec_validSource_17_valid;
  assign sinkVec_sinkWire_16_ready = sinkVec_8_0_ready;
  assign sinkVec_sinkWire_17_ready = sinkVec_8_1_ready;
  reg          maskUnitFirst_8;
  wire         tryToRead_8 = sinkVec_8_0_valid | sinkVec_8_1_valid;
  wire         sinkWire_8_valid = maskUnitFirst_8 ? sinkVec_8_0_valid : sinkVec_8_1_valid;
  wire [4:0]   sinkWire_8_bits_vs = maskUnitFirst_8 ? sinkVec_8_0_bits_vs : sinkVec_8_1_bits_vs;
  wire [1:0]   sinkWire_8_bits_readSource = maskUnitFirst_8 ? sinkVec_8_0_bits_readSource : sinkVec_8_1_bits_readSource;
  wire [1:0]   sinkWire_8_bits_offset = maskUnitFirst_8 ? sinkVec_8_0_bits_offset : sinkVec_8_1_bits_offset;
  wire [2:0]   sinkWire_8_bits_instructionIndex = maskUnitFirst_8 ? sinkVec_8_0_bits_instructionIndex : sinkVec_8_1_bits_instructionIndex;
  wire         sinkWire_8_ready;
  assign sinkVec_8_1_ready = sinkWire_8_ready & ~maskUnitFirst_8;
  assign sinkVec_8_0_ready = sinkWire_8_ready & maskUnitFirst_8;
  reg          accessDataValid_pipe_v_8;
  reg          accessDataValid_pipe_pipe_v_8;
  wire         accessDataValid_pipe_pipe_out_8_valid = accessDataValid_pipe_pipe_v_8;
  wire         accessDataSource_8_valid = accessDataValid_pipe_pipe_out_8_valid;
  reg          shifterReg_24_0_valid;
  reg  [31:0]  shifterReg_24_0_bits;
  wire         shifterValid_24 = shifterReg_24_0_valid | accessDataSource_8_valid;
  reg          accessDataValid_pipe_v_9;
  reg          accessDataValid_pipe_pipe_v_9;
  wire         accessDataValid_pipe_pipe_out_9_valid = accessDataValid_pipe_pipe_v_9;
  wire         accessDataSource_9_valid = accessDataValid_pipe_pipe_out_9_valid;
  reg          shifterReg_25_0_valid;
  reg  [31:0]  shifterReg_25_0_bits;
  wire         shifterValid_25 = shifterReg_25_0_valid | accessDataSource_9_valid;
  wire         sinkVec_tokenCheck_18;
  wire [4:0]   sinkVec_validSource_18_bits_vd = x22_4_0_bits_vd;
  wire [1:0]   sinkVec_validSource_18_bits_offset = x22_4_0_bits_offset;
  wire [3:0]   sinkVec_validSource_18_bits_mask = x22_4_0_bits_mask;
  wire [31:0]  sinkVec_validSource_18_bits_data = x22_4_0_bits_data;
  wire [2:0]   sinkVec_validSource_18_bits_instructionIndex = x22_4_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_19;
  wire [4:0]   sinkVec_validSource_19_bits_vd = x22_4_1_bits_vd;
  wire [1:0]   sinkVec_validSource_19_bits_offset = x22_4_1_bits_offset;
  wire [3:0]   sinkVec_validSource_19_bits_mask = x22_4_1_bits_mask;
  wire [31:0]  sinkVec_validSource_19_bits_data = x22_4_1_bits_data;
  wire         sinkVec_validSource_19_bits_last = x22_4_1_bits_last;
  wire [2:0]   sinkVec_validSource_19_bits_instructionIndex = x22_4_1_bits_instructionIndex;
  wire         sinkVec_9_0_ready;
  wire         sinkVec_queue_18_deq_ready = sinkVec_sinkWire_18_ready;
  wire         sinkVec_queue_18_deq_valid;
  wire [4:0]   sinkVec_queue_18_deq_bits_vd;
  wire         sinkVec_9_0_valid = sinkVec_sinkWire_18_valid;
  wire [1:0]   sinkVec_queue_18_deq_bits_offset;
  wire [4:0]   sinkVec_9_0_bits_vd = sinkVec_sinkWire_18_bits_vd;
  wire [3:0]   sinkVec_queue_18_deq_bits_mask;
  wire [1:0]   sinkVec_9_0_bits_offset = sinkVec_sinkWire_18_bits_offset;
  wire [31:0]  sinkVec_queue_18_deq_bits_data;
  wire [3:0]   sinkVec_9_0_bits_mask = sinkVec_sinkWire_18_bits_mask;
  wire         sinkVec_queue_18_deq_bits_last;
  wire [31:0]  sinkVec_9_0_bits_data = sinkVec_sinkWire_18_bits_data;
  wire [2:0]   sinkVec_queue_18_deq_bits_instructionIndex;
  wire         sinkVec_9_0_bits_last = sinkVec_sinkWire_18_bits_last;
  wire [2:0]   sinkVec_9_0_bits_instructionIndex = sinkVec_sinkWire_18_bits_instructionIndex;
  wire         sinkVec_validSink_18_valid;
  wire [4:0]   sinkVec_validSink_18_bits_vd;
  wire [1:0]   sinkVec_validSink_18_bits_offset;
  wire [3:0]   sinkVec_validSink_18_bits_mask;
  wire [31:0]  sinkVec_validSink_18_bits_data;
  wire [2:0]   sinkVec_validSink_18_bits_instructionIndex;
  assign sinkVec_sinkWire_18_valid = sinkVec_queue_18_deq_valid;
  assign sinkVec_sinkWire_18_bits_vd = sinkVec_queue_18_deq_bits_vd;
  assign sinkVec_sinkWire_18_bits_offset = sinkVec_queue_18_deq_bits_offset;
  assign sinkVec_sinkWire_18_bits_mask = sinkVec_queue_18_deq_bits_mask;
  assign sinkVec_sinkWire_18_bits_data = sinkVec_queue_18_deq_bits_data;
  assign sinkVec_sinkWire_18_bits_last = sinkVec_queue_18_deq_bits_last;
  assign sinkVec_sinkWire_18_bits_instructionIndex = sinkVec_queue_18_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_18_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_8 = {sinkVec_queue_18_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_18_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_18 = {sinkVec_queue_dataIn_lo_hi_8, sinkVec_queue_18_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_18_enq_bits_vd;
  wire [1:0]   sinkVec_queue_18_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_8 = {sinkVec_queue_18_enq_bits_vd, sinkVec_queue_18_enq_bits_offset};
  wire [3:0]   sinkVec_queue_18_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_18 = {sinkVec_queue_dataIn_hi_hi_8, sinkVec_queue_18_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_18 = {sinkVec_queue_dataIn_hi_18, sinkVec_queue_dataIn_lo_18};
  wire [2:0]   sinkVec_queue_dataOut_18_instructionIndex = _sinkVec_queue_fifo_18_data_out[2:0];
  wire         sinkVec_queue_dataOut_18_last = _sinkVec_queue_fifo_18_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_18_data = _sinkVec_queue_fifo_18_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_18_mask = _sinkVec_queue_fifo_18_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_18_offset = _sinkVec_queue_fifo_18_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_18_vd = _sinkVec_queue_fifo_18_data_out[46:42];
  wire         sinkVec_queue_18_enq_ready = ~_sinkVec_queue_fifo_18_full;
  wire         sinkVec_queue_18_enq_valid;
  assign sinkVec_queue_18_deq_valid = ~_sinkVec_queue_fifo_18_empty | sinkVec_queue_18_enq_valid;
  assign sinkVec_queue_18_deq_bits_vd = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_vd : sinkVec_queue_dataOut_18_vd;
  assign sinkVec_queue_18_deq_bits_offset = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_offset : sinkVec_queue_dataOut_18_offset;
  assign sinkVec_queue_18_deq_bits_mask = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_mask : sinkVec_queue_dataOut_18_mask;
  assign sinkVec_queue_18_deq_bits_data = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_data : sinkVec_queue_dataOut_18_data;
  assign sinkVec_queue_18_deq_bits_last = ~_sinkVec_queue_fifo_18_empty & sinkVec_queue_dataOut_18_last;
  assign sinkVec_queue_18_deq_bits_instructionIndex = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_instructionIndex : sinkVec_queue_dataOut_18_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_18;
  wire         sinkVec_releasePipe_pipe_out_18_valid = sinkVec_releasePipe_pipe_v_18;
  wire         x22_4_0_ready;
  wire         x22_4_0_valid;
  wire         sinkVec_validSource_18_valid = x22_4_0_ready & x22_4_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_18;
  wire [2:0]   sinkVec_tokenCheck_counterChange_18 = sinkVec_validSource_18_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_18 = ~(sinkVec_tokenCheck_counter_18[2]);
  assign x22_4_0_ready = sinkVec_tokenCheck_18;
  assign sinkVec_queue_18_enq_valid = sinkVec_validSink_18_valid;
  assign sinkVec_queue_18_enq_bits_vd = sinkVec_validSink_18_bits_vd;
  assign sinkVec_queue_18_enq_bits_offset = sinkVec_validSink_18_bits_offset;
  assign sinkVec_queue_18_enq_bits_mask = sinkVec_validSink_18_bits_mask;
  assign sinkVec_queue_18_enq_bits_data = sinkVec_validSink_18_bits_data;
  assign sinkVec_queue_18_enq_bits_instructionIndex = sinkVec_validSink_18_bits_instructionIndex;
  reg          sinkVec_shifterReg_18_0_valid;
  assign sinkVec_validSink_18_valid = sinkVec_shifterReg_18_0_valid;
  reg  [4:0]   sinkVec_shifterReg_18_0_bits_vd;
  assign sinkVec_validSink_18_bits_vd = sinkVec_shifterReg_18_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_18_0_bits_offset;
  assign sinkVec_validSink_18_bits_offset = sinkVec_shifterReg_18_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_18_0_bits_mask;
  assign sinkVec_validSink_18_bits_mask = sinkVec_shifterReg_18_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_18_0_bits_data;
  assign sinkVec_validSink_18_bits_data = sinkVec_shifterReg_18_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_18_0_bits_instructionIndex;
  assign sinkVec_validSink_18_bits_instructionIndex = sinkVec_shifterReg_18_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_18 = sinkVec_shifterReg_18_0_valid | sinkVec_validSource_18_valid;
  wire         sinkVec_9_1_ready;
  wire         sinkVec_queue_19_deq_ready = sinkVec_sinkWire_19_ready;
  wire         sinkVec_queue_19_deq_valid;
  wire [4:0]   sinkVec_queue_19_deq_bits_vd;
  wire         sinkVec_9_1_valid = sinkVec_sinkWire_19_valid;
  wire [1:0]   sinkVec_queue_19_deq_bits_offset;
  wire [4:0]   sinkVec_9_1_bits_vd = sinkVec_sinkWire_19_bits_vd;
  wire [3:0]   sinkVec_queue_19_deq_bits_mask;
  wire [1:0]   sinkVec_9_1_bits_offset = sinkVec_sinkWire_19_bits_offset;
  wire [31:0]  sinkVec_queue_19_deq_bits_data;
  wire [3:0]   sinkVec_9_1_bits_mask = sinkVec_sinkWire_19_bits_mask;
  wire         sinkVec_queue_19_deq_bits_last;
  wire [31:0]  sinkVec_9_1_bits_data = sinkVec_sinkWire_19_bits_data;
  wire [2:0]   sinkVec_queue_19_deq_bits_instructionIndex;
  wire         sinkVec_9_1_bits_last = sinkVec_sinkWire_19_bits_last;
  wire [2:0]   sinkVec_9_1_bits_instructionIndex = sinkVec_sinkWire_19_bits_instructionIndex;
  wire         sinkVec_validSink_19_valid;
  wire [4:0]   sinkVec_validSink_19_bits_vd;
  wire [1:0]   sinkVec_validSink_19_bits_offset;
  wire [3:0]   sinkVec_validSink_19_bits_mask;
  wire [31:0]  sinkVec_validSink_19_bits_data;
  wire         sinkVec_validSink_19_bits_last;
  wire [2:0]   sinkVec_validSink_19_bits_instructionIndex;
  assign sinkVec_sinkWire_19_valid = sinkVec_queue_19_deq_valid;
  assign sinkVec_sinkWire_19_bits_vd = sinkVec_queue_19_deq_bits_vd;
  assign sinkVec_sinkWire_19_bits_offset = sinkVec_queue_19_deq_bits_offset;
  assign sinkVec_sinkWire_19_bits_mask = sinkVec_queue_19_deq_bits_mask;
  assign sinkVec_sinkWire_19_bits_data = sinkVec_queue_19_deq_bits_data;
  assign sinkVec_sinkWire_19_bits_last = sinkVec_queue_19_deq_bits_last;
  assign sinkVec_sinkWire_19_bits_instructionIndex = sinkVec_queue_19_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_19_enq_bits_data;
  wire         sinkVec_queue_19_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_9 = {sinkVec_queue_19_enq_bits_data, sinkVec_queue_19_enq_bits_last};
  wire [2:0]   sinkVec_queue_19_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_19 = {sinkVec_queue_dataIn_lo_hi_9, sinkVec_queue_19_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_19_enq_bits_vd;
  wire [1:0]   sinkVec_queue_19_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_9 = {sinkVec_queue_19_enq_bits_vd, sinkVec_queue_19_enq_bits_offset};
  wire [3:0]   sinkVec_queue_19_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_19 = {sinkVec_queue_dataIn_hi_hi_9, sinkVec_queue_19_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_19 = {sinkVec_queue_dataIn_hi_19, sinkVec_queue_dataIn_lo_19};
  wire [2:0]   sinkVec_queue_dataOut_19_instructionIndex = _sinkVec_queue_fifo_19_data_out[2:0];
  wire         sinkVec_queue_dataOut_19_last = _sinkVec_queue_fifo_19_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_19_data = _sinkVec_queue_fifo_19_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_19_mask = _sinkVec_queue_fifo_19_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_19_offset = _sinkVec_queue_fifo_19_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_19_vd = _sinkVec_queue_fifo_19_data_out[46:42];
  wire         sinkVec_queue_19_enq_ready = ~_sinkVec_queue_fifo_19_full;
  wire         sinkVec_queue_19_enq_valid;
  assign sinkVec_queue_19_deq_valid = ~_sinkVec_queue_fifo_19_empty | sinkVec_queue_19_enq_valid;
  assign sinkVec_queue_19_deq_bits_vd = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_vd : sinkVec_queue_dataOut_19_vd;
  assign sinkVec_queue_19_deq_bits_offset = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_offset : sinkVec_queue_dataOut_19_offset;
  assign sinkVec_queue_19_deq_bits_mask = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_mask : sinkVec_queue_dataOut_19_mask;
  assign sinkVec_queue_19_deq_bits_data = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_data : sinkVec_queue_dataOut_19_data;
  assign sinkVec_queue_19_deq_bits_last = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_last : sinkVec_queue_dataOut_19_last;
  assign sinkVec_queue_19_deq_bits_instructionIndex = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_instructionIndex : sinkVec_queue_dataOut_19_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_19;
  wire         sinkVec_releasePipe_pipe_out_19_valid = sinkVec_releasePipe_pipe_v_19;
  wire         x22_4_1_ready;
  wire         x22_4_1_valid;
  wire         sinkVec_validSource_19_valid = x22_4_1_ready & x22_4_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_19;
  wire [2:0]   sinkVec_tokenCheck_counterChange_19 = sinkVec_validSource_19_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_19 = ~(sinkVec_tokenCheck_counter_19[2]);
  assign x22_4_1_ready = sinkVec_tokenCheck_19;
  assign sinkVec_queue_19_enq_valid = sinkVec_validSink_19_valid;
  assign sinkVec_queue_19_enq_bits_vd = sinkVec_validSink_19_bits_vd;
  assign sinkVec_queue_19_enq_bits_offset = sinkVec_validSink_19_bits_offset;
  assign sinkVec_queue_19_enq_bits_mask = sinkVec_validSink_19_bits_mask;
  assign sinkVec_queue_19_enq_bits_data = sinkVec_validSink_19_bits_data;
  assign sinkVec_queue_19_enq_bits_last = sinkVec_validSink_19_bits_last;
  assign sinkVec_queue_19_enq_bits_instructionIndex = sinkVec_validSink_19_bits_instructionIndex;
  reg          sinkVec_shifterReg_19_0_valid;
  assign sinkVec_validSink_19_valid = sinkVec_shifterReg_19_0_valid;
  reg  [4:0]   sinkVec_shifterReg_19_0_bits_vd;
  assign sinkVec_validSink_19_bits_vd = sinkVec_shifterReg_19_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_19_0_bits_offset;
  assign sinkVec_validSink_19_bits_offset = sinkVec_shifterReg_19_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_19_0_bits_mask;
  assign sinkVec_validSink_19_bits_mask = sinkVec_shifterReg_19_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_19_0_bits_data;
  assign sinkVec_validSink_19_bits_data = sinkVec_shifterReg_19_0_bits_data;
  reg          sinkVec_shifterReg_19_0_bits_last;
  assign sinkVec_validSink_19_bits_last = sinkVec_shifterReg_19_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_19_0_bits_instructionIndex;
  assign sinkVec_validSink_19_bits_instructionIndex = sinkVec_shifterReg_19_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_19 = sinkVec_shifterReg_19_0_valid | sinkVec_validSource_19_valid;
  assign sinkVec_sinkWire_18_ready = sinkVec_9_0_ready;
  assign sinkVec_sinkWire_19_ready = sinkVec_9_1_ready;
  reg          maskUnitFirst_9;
  wire         tryToRead_9 = sinkVec_9_0_valid | sinkVec_9_1_valid;
  wire         sinkWire_9_valid = maskUnitFirst_9 ? sinkVec_9_0_valid : sinkVec_9_1_valid;
  wire [4:0]   sinkWire_9_bits_vd = maskUnitFirst_9 ? sinkVec_9_0_bits_vd : sinkVec_9_1_bits_vd;
  wire [1:0]   sinkWire_9_bits_offset = maskUnitFirst_9 ? sinkVec_9_0_bits_offset : sinkVec_9_1_bits_offset;
  wire [3:0]   sinkWire_9_bits_mask = maskUnitFirst_9 ? sinkVec_9_0_bits_mask : sinkVec_9_1_bits_mask;
  wire [31:0]  sinkWire_9_bits_data = maskUnitFirst_9 ? sinkVec_9_0_bits_data : sinkVec_9_1_bits_data;
  wire         sinkWire_9_bits_last = maskUnitFirst_9 ? sinkVec_9_0_bits_last : sinkVec_9_1_bits_last;
  wire [2:0]   sinkWire_9_bits_instructionIndex = maskUnitFirst_9 ? sinkVec_9_0_bits_instructionIndex : sinkVec_9_1_bits_instructionIndex;
  wire         sinkWire_9_ready;
  assign sinkVec_9_1_ready = sinkWire_9_ready & ~maskUnitFirst_9;
  assign sinkVec_9_0_ready = sinkWire_9_ready & maskUnitFirst_9;
  reg          view__writeRelease_4_pipe_v;
  wire         view__writeRelease_4_pipe_out_valid = view__writeRelease_4_pipe_v;
  reg          pipe_v_12;
  wire         pipe_out_8_valid = pipe_v_12;
  wire         _probeWire_writeQueueEnqVec_4_valid_T = x22_4_0_ready & _maskUnit_exeResp_4_valid;
  reg          instructionFinishedPipe_pipe_v_4;
  wire         instructionFinishedPipe_pipe_out_4_valid = instructionFinishedPipe_pipe_v_4;
  reg  [7:0]   instructionFinishedPipe_pipe_b_4;
  wire [7:0]   instructionFinishedPipe_pipe_out_4_bits = instructionFinishedPipe_pipe_b_4;
  wire         instructionFinished_4_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_4_bits);
  assign vxsatReportVec_4 = _laneVec_4_vxsatReport[3:0];
  reg          pipe_v_13;
  reg  [31:0]  pipe_b_13;
  reg          pipe_pipe_v_4;
  wire         pipe_pipe_out_4_valid = pipe_pipe_v_4;
  reg  [31:0]  pipe_pipe_b_4;
  wire [31:0]  pipe_pipe_out_4_bits = pipe_pipe_b_4;
  reg          view__laneMaskSelect_4_pipe_v;
  reg  [5:0]   view__laneMaskSelect_4_pipe_b;
  reg          view__laneMaskSelect_4_pipe_pipe_v;
  wire         view__laneMaskSelect_4_pipe_pipe_out_valid = view__laneMaskSelect_4_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_4_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_4_pipe_pipe_out_bits = view__laneMaskSelect_4_pipe_pipe_b;
  reg          view__laneMaskSewSelect_4_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_4_pipe_b;
  reg          view__laneMaskSewSelect_4_pipe_pipe_v;
  wire         view__laneMaskSewSelect_4_pipe_pipe_out_valid = view__laneMaskSewSelect_4_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_4_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_4_pipe_pipe_out_bits = view__laneMaskSewSelect_4_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_4;
  wire         lsuLastPipe_pipe_out_4_valid = lsuLastPipe_pipe_v_4;
  reg  [7:0]   lsuLastPipe_pipe_b_4;
  wire [7:0]   lsuLastPipe_pipe_out_4_bits = lsuLastPipe_pipe_b_4;
  reg          maskLastPipe_pipe_v_4;
  wire         maskLastPipe_pipe_out_4_valid = maskLastPipe_pipe_v_4;
  reg  [7:0]   maskLastPipe_pipe_b_4;
  wire [7:0]   maskLastPipe_pipe_out_4_bits = maskLastPipe_pipe_b_4;
  wire [5:0]   writeCounter_4 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h10};
  reg          pipe_v_14;
  wire         pipe_out_9_valid = pipe_v_14;
  reg  [5:0]   pipe_b_14;
  wire [5:0]   pipe_out_9_bits = pipe_b_14;
  assign laneRequestSinkWire_5_ready = ~laneRequestSinkWire_5_bits_issueInst | _laneVec_5_laneRequest_ready;
  wire         sinkVec_tokenCheck_20;
  wire [4:0]   sinkVec_validSource_20_bits_vs = x13_5_0_bits_vs;
  wire [1:0]   sinkVec_validSource_20_bits_offset = x13_5_0_bits_offset;
  wire [2:0]   sinkVec_validSource_20_bits_instructionIndex = x13_5_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_21;
  wire [4:0]   sinkVec_validSource_21_bits_vs = x13_5_1_bits_vs;
  wire [1:0]   sinkVec_validSource_21_bits_offset = x13_5_1_bits_offset;
  wire [2:0]   sinkVec_validSource_21_bits_instructionIndex = x13_5_1_bits_instructionIndex;
  wire         sinkVec_10_0_ready;
  wire         sinkVec_queue_20_deq_ready = sinkVec_sinkWire_20_ready;
  wire         sinkVec_queue_20_deq_valid;
  wire [4:0]   sinkVec_queue_20_deq_bits_vs;
  wire         sinkVec_10_0_valid = sinkVec_sinkWire_20_valid;
  wire [1:0]   sinkVec_queue_20_deq_bits_readSource;
  wire [4:0]   sinkVec_10_0_bits_vs = sinkVec_sinkWire_20_bits_vs;
  wire [1:0]   sinkVec_queue_20_deq_bits_offset;
  wire [1:0]   sinkVec_10_0_bits_readSource = sinkVec_sinkWire_20_bits_readSource;
  wire [2:0]   sinkVec_queue_20_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_10_0_bits_offset = sinkVec_sinkWire_20_bits_offset;
  wire [2:0]   sinkVec_10_0_bits_instructionIndex = sinkVec_sinkWire_20_bits_instructionIndex;
  wire         sinkVec_validSink_20_valid;
  wire [4:0]   sinkVec_validSink_20_bits_vs;
  wire [1:0]   sinkVec_validSink_20_bits_readSource;
  wire [1:0]   sinkVec_validSink_20_bits_offset;
  wire [2:0]   sinkVec_validSink_20_bits_instructionIndex;
  assign sinkVec_sinkWire_20_valid = sinkVec_queue_20_deq_valid;
  assign sinkVec_sinkWire_20_bits_vs = sinkVec_queue_20_deq_bits_vs;
  assign sinkVec_sinkWire_20_bits_readSource = sinkVec_queue_20_deq_bits_readSource;
  assign sinkVec_sinkWire_20_bits_offset = sinkVec_queue_20_deq_bits_offset;
  assign sinkVec_sinkWire_20_bits_instructionIndex = sinkVec_queue_20_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_20_enq_bits_offset;
  wire [2:0]   sinkVec_queue_20_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_20 = {sinkVec_queue_20_enq_bits_offset, sinkVec_queue_20_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_20_enq_bits_vs;
  wire [1:0]   sinkVec_queue_20_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_20 = {sinkVec_queue_20_enq_bits_vs, sinkVec_queue_20_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_20 = {sinkVec_queue_dataIn_hi_20, sinkVec_queue_dataIn_lo_20};
  wire [2:0]   sinkVec_queue_dataOut_20_instructionIndex = _sinkVec_queue_fifo_20_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_20_offset = _sinkVec_queue_fifo_20_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_20_readSource = _sinkVec_queue_fifo_20_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_20_vs = _sinkVec_queue_fifo_20_data_out[11:7];
  wire         sinkVec_queue_20_enq_ready = ~_sinkVec_queue_fifo_20_full;
  wire         sinkVec_queue_20_enq_valid;
  assign sinkVec_queue_20_deq_valid = ~_sinkVec_queue_fifo_20_empty | sinkVec_queue_20_enq_valid;
  assign sinkVec_queue_20_deq_bits_vs = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_vs : sinkVec_queue_dataOut_20_vs;
  assign sinkVec_queue_20_deq_bits_readSource = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_readSource : sinkVec_queue_dataOut_20_readSource;
  assign sinkVec_queue_20_deq_bits_offset = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_offset : sinkVec_queue_dataOut_20_offset;
  assign sinkVec_queue_20_deq_bits_instructionIndex = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_instructionIndex : sinkVec_queue_dataOut_20_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_20;
  wire         sinkVec_releasePipe_pipe_out_20_valid = sinkVec_releasePipe_pipe_v_20;
  wire         x13_5_0_ready;
  wire         x13_5_0_valid;
  wire         sinkVec_validSource_20_valid = x13_5_0_ready & x13_5_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_20;
  wire [2:0]   sinkVec_tokenCheck_counterChange_20 = sinkVec_validSource_20_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_20 = ~(sinkVec_tokenCheck_counter_20[2]);
  assign x13_5_0_ready = sinkVec_tokenCheck_20;
  assign sinkVec_queue_20_enq_valid = sinkVec_validSink_20_valid;
  assign sinkVec_queue_20_enq_bits_vs = sinkVec_validSink_20_bits_vs;
  assign sinkVec_queue_20_enq_bits_readSource = sinkVec_validSink_20_bits_readSource;
  assign sinkVec_queue_20_enq_bits_offset = sinkVec_validSink_20_bits_offset;
  assign sinkVec_queue_20_enq_bits_instructionIndex = sinkVec_validSink_20_bits_instructionIndex;
  reg          sinkVec_shifterReg_20_0_valid;
  assign sinkVec_validSink_20_valid = sinkVec_shifterReg_20_0_valid;
  reg  [4:0]   sinkVec_shifterReg_20_0_bits_vs;
  assign sinkVec_validSink_20_bits_vs = sinkVec_shifterReg_20_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_20_0_bits_readSource;
  assign sinkVec_validSink_20_bits_readSource = sinkVec_shifterReg_20_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_20_0_bits_offset;
  assign sinkVec_validSink_20_bits_offset = sinkVec_shifterReg_20_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_20_0_bits_instructionIndex;
  assign sinkVec_validSink_20_bits_instructionIndex = sinkVec_shifterReg_20_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_20 = sinkVec_shifterReg_20_0_valid | sinkVec_validSource_20_valid;
  wire         sinkVec_10_1_ready;
  wire         sinkVec_queue_21_deq_ready = sinkVec_sinkWire_21_ready;
  wire         sinkVec_queue_21_deq_valid;
  wire [4:0]   sinkVec_queue_21_deq_bits_vs;
  wire         sinkVec_10_1_valid = sinkVec_sinkWire_21_valid;
  wire [1:0]   sinkVec_queue_21_deq_bits_readSource;
  wire [4:0]   sinkVec_10_1_bits_vs = sinkVec_sinkWire_21_bits_vs;
  wire [1:0]   sinkVec_queue_21_deq_bits_offset;
  wire [1:0]   sinkVec_10_1_bits_readSource = sinkVec_sinkWire_21_bits_readSource;
  wire [2:0]   sinkVec_queue_21_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_10_1_bits_offset = sinkVec_sinkWire_21_bits_offset;
  wire [2:0]   sinkVec_10_1_bits_instructionIndex = sinkVec_sinkWire_21_bits_instructionIndex;
  wire         sinkVec_validSink_21_valid;
  wire [4:0]   sinkVec_validSink_21_bits_vs;
  wire [1:0]   sinkVec_validSink_21_bits_readSource;
  wire [1:0]   sinkVec_validSink_21_bits_offset;
  wire [2:0]   sinkVec_validSink_21_bits_instructionIndex;
  assign sinkVec_sinkWire_21_valid = sinkVec_queue_21_deq_valid;
  assign sinkVec_sinkWire_21_bits_vs = sinkVec_queue_21_deq_bits_vs;
  assign sinkVec_sinkWire_21_bits_readSource = sinkVec_queue_21_deq_bits_readSource;
  assign sinkVec_sinkWire_21_bits_offset = sinkVec_queue_21_deq_bits_offset;
  assign sinkVec_sinkWire_21_bits_instructionIndex = sinkVec_queue_21_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_21_enq_bits_offset;
  wire [2:0]   sinkVec_queue_21_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_21 = {sinkVec_queue_21_enq_bits_offset, sinkVec_queue_21_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_21_enq_bits_vs;
  wire [1:0]   sinkVec_queue_21_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_21 = {sinkVec_queue_21_enq_bits_vs, sinkVec_queue_21_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_21 = {sinkVec_queue_dataIn_hi_21, sinkVec_queue_dataIn_lo_21};
  wire [2:0]   sinkVec_queue_dataOut_21_instructionIndex = _sinkVec_queue_fifo_21_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_21_offset = _sinkVec_queue_fifo_21_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_21_readSource = _sinkVec_queue_fifo_21_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_21_vs = _sinkVec_queue_fifo_21_data_out[11:7];
  wire         sinkVec_queue_21_enq_ready = ~_sinkVec_queue_fifo_21_full;
  wire         sinkVec_queue_21_enq_valid;
  assign sinkVec_queue_21_deq_valid = ~_sinkVec_queue_fifo_21_empty | sinkVec_queue_21_enq_valid;
  assign sinkVec_queue_21_deq_bits_vs = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_vs : sinkVec_queue_dataOut_21_vs;
  assign sinkVec_queue_21_deq_bits_readSource = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_readSource : sinkVec_queue_dataOut_21_readSource;
  assign sinkVec_queue_21_deq_bits_offset = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_offset : sinkVec_queue_dataOut_21_offset;
  assign sinkVec_queue_21_deq_bits_instructionIndex = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_instructionIndex : sinkVec_queue_dataOut_21_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_21;
  wire         sinkVec_releasePipe_pipe_out_21_valid = sinkVec_releasePipe_pipe_v_21;
  wire         x13_5_1_ready;
  wire         x13_5_1_valid;
  wire         sinkVec_validSource_21_valid = x13_5_1_ready & x13_5_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_21;
  wire [2:0]   sinkVec_tokenCheck_counterChange_21 = sinkVec_validSource_21_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_21 = ~(sinkVec_tokenCheck_counter_21[2]);
  assign x13_5_1_ready = sinkVec_tokenCheck_21;
  assign sinkVec_queue_21_enq_valid = sinkVec_validSink_21_valid;
  assign sinkVec_queue_21_enq_bits_vs = sinkVec_validSink_21_bits_vs;
  assign sinkVec_queue_21_enq_bits_readSource = sinkVec_validSink_21_bits_readSource;
  assign sinkVec_queue_21_enq_bits_offset = sinkVec_validSink_21_bits_offset;
  assign sinkVec_queue_21_enq_bits_instructionIndex = sinkVec_validSink_21_bits_instructionIndex;
  reg          sinkVec_shifterReg_21_0_valid;
  assign sinkVec_validSink_21_valid = sinkVec_shifterReg_21_0_valid;
  reg  [4:0]   sinkVec_shifterReg_21_0_bits_vs;
  assign sinkVec_validSink_21_bits_vs = sinkVec_shifterReg_21_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_21_0_bits_readSource;
  assign sinkVec_validSink_21_bits_readSource = sinkVec_shifterReg_21_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_21_0_bits_offset;
  assign sinkVec_validSink_21_bits_offset = sinkVec_shifterReg_21_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_21_0_bits_instructionIndex;
  assign sinkVec_validSink_21_bits_instructionIndex = sinkVec_shifterReg_21_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_21 = sinkVec_shifterReg_21_0_valid | sinkVec_validSource_21_valid;
  assign sinkVec_sinkWire_20_ready = sinkVec_10_0_ready;
  assign sinkVec_sinkWire_21_ready = sinkVec_10_1_ready;
  reg          maskUnitFirst_10;
  wire         tryToRead_10 = sinkVec_10_0_valid | sinkVec_10_1_valid;
  wire         sinkWire_10_valid = maskUnitFirst_10 ? sinkVec_10_0_valid : sinkVec_10_1_valid;
  wire [4:0]   sinkWire_10_bits_vs = maskUnitFirst_10 ? sinkVec_10_0_bits_vs : sinkVec_10_1_bits_vs;
  wire [1:0]   sinkWire_10_bits_readSource = maskUnitFirst_10 ? sinkVec_10_0_bits_readSource : sinkVec_10_1_bits_readSource;
  wire [1:0]   sinkWire_10_bits_offset = maskUnitFirst_10 ? sinkVec_10_0_bits_offset : sinkVec_10_1_bits_offset;
  wire [2:0]   sinkWire_10_bits_instructionIndex = maskUnitFirst_10 ? sinkVec_10_0_bits_instructionIndex : sinkVec_10_1_bits_instructionIndex;
  wire         sinkWire_10_ready;
  assign sinkVec_10_1_ready = sinkWire_10_ready & ~maskUnitFirst_10;
  assign sinkVec_10_0_ready = sinkWire_10_ready & maskUnitFirst_10;
  reg          accessDataValid_pipe_v_10;
  reg          accessDataValid_pipe_pipe_v_10;
  wire         accessDataValid_pipe_pipe_out_10_valid = accessDataValid_pipe_pipe_v_10;
  wire         accessDataSource_10_valid = accessDataValid_pipe_pipe_out_10_valid;
  reg          shifterReg_26_0_valid;
  reg  [31:0]  shifterReg_26_0_bits;
  wire         shifterValid_26 = shifterReg_26_0_valid | accessDataSource_10_valid;
  reg          accessDataValid_pipe_v_11;
  reg          accessDataValid_pipe_pipe_v_11;
  wire         accessDataValid_pipe_pipe_out_11_valid = accessDataValid_pipe_pipe_v_11;
  wire         accessDataSource_11_valid = accessDataValid_pipe_pipe_out_11_valid;
  reg          shifterReg_27_0_valid;
  reg  [31:0]  shifterReg_27_0_bits;
  wire         shifterValid_27 = shifterReg_27_0_valid | accessDataSource_11_valid;
  wire         sinkVec_tokenCheck_22;
  wire [4:0]   sinkVec_validSource_22_bits_vd = x22_5_0_bits_vd;
  wire [1:0]   sinkVec_validSource_22_bits_offset = x22_5_0_bits_offset;
  wire [3:0]   sinkVec_validSource_22_bits_mask = x22_5_0_bits_mask;
  wire [31:0]  sinkVec_validSource_22_bits_data = x22_5_0_bits_data;
  wire [2:0]   sinkVec_validSource_22_bits_instructionIndex = x22_5_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_23;
  wire [4:0]   sinkVec_validSource_23_bits_vd = x22_5_1_bits_vd;
  wire [1:0]   sinkVec_validSource_23_bits_offset = x22_5_1_bits_offset;
  wire [3:0]   sinkVec_validSource_23_bits_mask = x22_5_1_bits_mask;
  wire [31:0]  sinkVec_validSource_23_bits_data = x22_5_1_bits_data;
  wire         sinkVec_validSource_23_bits_last = x22_5_1_bits_last;
  wire [2:0]   sinkVec_validSource_23_bits_instructionIndex = x22_5_1_bits_instructionIndex;
  wire         sinkVec_11_0_ready;
  wire         sinkVec_queue_22_deq_ready = sinkVec_sinkWire_22_ready;
  wire         sinkVec_queue_22_deq_valid;
  wire [4:0]   sinkVec_queue_22_deq_bits_vd;
  wire         sinkVec_11_0_valid = sinkVec_sinkWire_22_valid;
  wire [1:0]   sinkVec_queue_22_deq_bits_offset;
  wire [4:0]   sinkVec_11_0_bits_vd = sinkVec_sinkWire_22_bits_vd;
  wire [3:0]   sinkVec_queue_22_deq_bits_mask;
  wire [1:0]   sinkVec_11_0_bits_offset = sinkVec_sinkWire_22_bits_offset;
  wire [31:0]  sinkVec_queue_22_deq_bits_data;
  wire [3:0]   sinkVec_11_0_bits_mask = sinkVec_sinkWire_22_bits_mask;
  wire         sinkVec_queue_22_deq_bits_last;
  wire [31:0]  sinkVec_11_0_bits_data = sinkVec_sinkWire_22_bits_data;
  wire [2:0]   sinkVec_queue_22_deq_bits_instructionIndex;
  wire         sinkVec_11_0_bits_last = sinkVec_sinkWire_22_bits_last;
  wire [2:0]   sinkVec_11_0_bits_instructionIndex = sinkVec_sinkWire_22_bits_instructionIndex;
  wire         sinkVec_validSink_22_valid;
  wire [4:0]   sinkVec_validSink_22_bits_vd;
  wire [1:0]   sinkVec_validSink_22_bits_offset;
  wire [3:0]   sinkVec_validSink_22_bits_mask;
  wire [31:0]  sinkVec_validSink_22_bits_data;
  wire [2:0]   sinkVec_validSink_22_bits_instructionIndex;
  assign sinkVec_sinkWire_22_valid = sinkVec_queue_22_deq_valid;
  assign sinkVec_sinkWire_22_bits_vd = sinkVec_queue_22_deq_bits_vd;
  assign sinkVec_sinkWire_22_bits_offset = sinkVec_queue_22_deq_bits_offset;
  assign sinkVec_sinkWire_22_bits_mask = sinkVec_queue_22_deq_bits_mask;
  assign sinkVec_sinkWire_22_bits_data = sinkVec_queue_22_deq_bits_data;
  assign sinkVec_sinkWire_22_bits_last = sinkVec_queue_22_deq_bits_last;
  assign sinkVec_sinkWire_22_bits_instructionIndex = sinkVec_queue_22_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_22_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_10 = {sinkVec_queue_22_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_22_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_22 = {sinkVec_queue_dataIn_lo_hi_10, sinkVec_queue_22_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_22_enq_bits_vd;
  wire [1:0]   sinkVec_queue_22_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_10 = {sinkVec_queue_22_enq_bits_vd, sinkVec_queue_22_enq_bits_offset};
  wire [3:0]   sinkVec_queue_22_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_22 = {sinkVec_queue_dataIn_hi_hi_10, sinkVec_queue_22_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_22 = {sinkVec_queue_dataIn_hi_22, sinkVec_queue_dataIn_lo_22};
  wire [2:0]   sinkVec_queue_dataOut_22_instructionIndex = _sinkVec_queue_fifo_22_data_out[2:0];
  wire         sinkVec_queue_dataOut_22_last = _sinkVec_queue_fifo_22_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_22_data = _sinkVec_queue_fifo_22_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_22_mask = _sinkVec_queue_fifo_22_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_22_offset = _sinkVec_queue_fifo_22_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_22_vd = _sinkVec_queue_fifo_22_data_out[46:42];
  wire         sinkVec_queue_22_enq_ready = ~_sinkVec_queue_fifo_22_full;
  wire         sinkVec_queue_22_enq_valid;
  assign sinkVec_queue_22_deq_valid = ~_sinkVec_queue_fifo_22_empty | sinkVec_queue_22_enq_valid;
  assign sinkVec_queue_22_deq_bits_vd = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_vd : sinkVec_queue_dataOut_22_vd;
  assign sinkVec_queue_22_deq_bits_offset = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_offset : sinkVec_queue_dataOut_22_offset;
  assign sinkVec_queue_22_deq_bits_mask = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_mask : sinkVec_queue_dataOut_22_mask;
  assign sinkVec_queue_22_deq_bits_data = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_data : sinkVec_queue_dataOut_22_data;
  assign sinkVec_queue_22_deq_bits_last = ~_sinkVec_queue_fifo_22_empty & sinkVec_queue_dataOut_22_last;
  assign sinkVec_queue_22_deq_bits_instructionIndex = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_instructionIndex : sinkVec_queue_dataOut_22_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_22;
  wire         sinkVec_releasePipe_pipe_out_22_valid = sinkVec_releasePipe_pipe_v_22;
  wire         x22_5_0_ready;
  wire         x22_5_0_valid;
  wire         sinkVec_validSource_22_valid = x22_5_0_ready & x22_5_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_22;
  wire [2:0]   sinkVec_tokenCheck_counterChange_22 = sinkVec_validSource_22_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_22 = ~(sinkVec_tokenCheck_counter_22[2]);
  assign x22_5_0_ready = sinkVec_tokenCheck_22;
  assign sinkVec_queue_22_enq_valid = sinkVec_validSink_22_valid;
  assign sinkVec_queue_22_enq_bits_vd = sinkVec_validSink_22_bits_vd;
  assign sinkVec_queue_22_enq_bits_offset = sinkVec_validSink_22_bits_offset;
  assign sinkVec_queue_22_enq_bits_mask = sinkVec_validSink_22_bits_mask;
  assign sinkVec_queue_22_enq_bits_data = sinkVec_validSink_22_bits_data;
  assign sinkVec_queue_22_enq_bits_instructionIndex = sinkVec_validSink_22_bits_instructionIndex;
  reg          sinkVec_shifterReg_22_0_valid;
  assign sinkVec_validSink_22_valid = sinkVec_shifterReg_22_0_valid;
  reg  [4:0]   sinkVec_shifterReg_22_0_bits_vd;
  assign sinkVec_validSink_22_bits_vd = sinkVec_shifterReg_22_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_22_0_bits_offset;
  assign sinkVec_validSink_22_bits_offset = sinkVec_shifterReg_22_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_22_0_bits_mask;
  assign sinkVec_validSink_22_bits_mask = sinkVec_shifterReg_22_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_22_0_bits_data;
  assign sinkVec_validSink_22_bits_data = sinkVec_shifterReg_22_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_22_0_bits_instructionIndex;
  assign sinkVec_validSink_22_bits_instructionIndex = sinkVec_shifterReg_22_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_22 = sinkVec_shifterReg_22_0_valid | sinkVec_validSource_22_valid;
  wire         sinkVec_11_1_ready;
  wire         sinkVec_queue_23_deq_ready = sinkVec_sinkWire_23_ready;
  wire         sinkVec_queue_23_deq_valid;
  wire [4:0]   sinkVec_queue_23_deq_bits_vd;
  wire         sinkVec_11_1_valid = sinkVec_sinkWire_23_valid;
  wire [1:0]   sinkVec_queue_23_deq_bits_offset;
  wire [4:0]   sinkVec_11_1_bits_vd = sinkVec_sinkWire_23_bits_vd;
  wire [3:0]   sinkVec_queue_23_deq_bits_mask;
  wire [1:0]   sinkVec_11_1_bits_offset = sinkVec_sinkWire_23_bits_offset;
  wire [31:0]  sinkVec_queue_23_deq_bits_data;
  wire [3:0]   sinkVec_11_1_bits_mask = sinkVec_sinkWire_23_bits_mask;
  wire         sinkVec_queue_23_deq_bits_last;
  wire [31:0]  sinkVec_11_1_bits_data = sinkVec_sinkWire_23_bits_data;
  wire [2:0]   sinkVec_queue_23_deq_bits_instructionIndex;
  wire         sinkVec_11_1_bits_last = sinkVec_sinkWire_23_bits_last;
  wire [2:0]   sinkVec_11_1_bits_instructionIndex = sinkVec_sinkWire_23_bits_instructionIndex;
  wire         sinkVec_validSink_23_valid;
  wire [4:0]   sinkVec_validSink_23_bits_vd;
  wire [1:0]   sinkVec_validSink_23_bits_offset;
  wire [3:0]   sinkVec_validSink_23_bits_mask;
  wire [31:0]  sinkVec_validSink_23_bits_data;
  wire         sinkVec_validSink_23_bits_last;
  wire [2:0]   sinkVec_validSink_23_bits_instructionIndex;
  assign sinkVec_sinkWire_23_valid = sinkVec_queue_23_deq_valid;
  assign sinkVec_sinkWire_23_bits_vd = sinkVec_queue_23_deq_bits_vd;
  assign sinkVec_sinkWire_23_bits_offset = sinkVec_queue_23_deq_bits_offset;
  assign sinkVec_sinkWire_23_bits_mask = sinkVec_queue_23_deq_bits_mask;
  assign sinkVec_sinkWire_23_bits_data = sinkVec_queue_23_deq_bits_data;
  assign sinkVec_sinkWire_23_bits_last = sinkVec_queue_23_deq_bits_last;
  assign sinkVec_sinkWire_23_bits_instructionIndex = sinkVec_queue_23_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_23_enq_bits_data;
  wire         sinkVec_queue_23_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_11 = {sinkVec_queue_23_enq_bits_data, sinkVec_queue_23_enq_bits_last};
  wire [2:0]   sinkVec_queue_23_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_23 = {sinkVec_queue_dataIn_lo_hi_11, sinkVec_queue_23_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_23_enq_bits_vd;
  wire [1:0]   sinkVec_queue_23_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_11 = {sinkVec_queue_23_enq_bits_vd, sinkVec_queue_23_enq_bits_offset};
  wire [3:0]   sinkVec_queue_23_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_23 = {sinkVec_queue_dataIn_hi_hi_11, sinkVec_queue_23_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_23 = {sinkVec_queue_dataIn_hi_23, sinkVec_queue_dataIn_lo_23};
  wire [2:0]   sinkVec_queue_dataOut_23_instructionIndex = _sinkVec_queue_fifo_23_data_out[2:0];
  wire         sinkVec_queue_dataOut_23_last = _sinkVec_queue_fifo_23_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_23_data = _sinkVec_queue_fifo_23_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_23_mask = _sinkVec_queue_fifo_23_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_23_offset = _sinkVec_queue_fifo_23_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_23_vd = _sinkVec_queue_fifo_23_data_out[46:42];
  wire         sinkVec_queue_23_enq_ready = ~_sinkVec_queue_fifo_23_full;
  wire         sinkVec_queue_23_enq_valid;
  assign sinkVec_queue_23_deq_valid = ~_sinkVec_queue_fifo_23_empty | sinkVec_queue_23_enq_valid;
  assign sinkVec_queue_23_deq_bits_vd = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_vd : sinkVec_queue_dataOut_23_vd;
  assign sinkVec_queue_23_deq_bits_offset = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_offset : sinkVec_queue_dataOut_23_offset;
  assign sinkVec_queue_23_deq_bits_mask = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_mask : sinkVec_queue_dataOut_23_mask;
  assign sinkVec_queue_23_deq_bits_data = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_data : sinkVec_queue_dataOut_23_data;
  assign sinkVec_queue_23_deq_bits_last = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_last : sinkVec_queue_dataOut_23_last;
  assign sinkVec_queue_23_deq_bits_instructionIndex = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_instructionIndex : sinkVec_queue_dataOut_23_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_23;
  wire         sinkVec_releasePipe_pipe_out_23_valid = sinkVec_releasePipe_pipe_v_23;
  wire         x22_5_1_ready;
  wire         x22_5_1_valid;
  wire         sinkVec_validSource_23_valid = x22_5_1_ready & x22_5_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_23;
  wire [2:0]   sinkVec_tokenCheck_counterChange_23 = sinkVec_validSource_23_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_23 = ~(sinkVec_tokenCheck_counter_23[2]);
  assign x22_5_1_ready = sinkVec_tokenCheck_23;
  assign sinkVec_queue_23_enq_valid = sinkVec_validSink_23_valid;
  assign sinkVec_queue_23_enq_bits_vd = sinkVec_validSink_23_bits_vd;
  assign sinkVec_queue_23_enq_bits_offset = sinkVec_validSink_23_bits_offset;
  assign sinkVec_queue_23_enq_bits_mask = sinkVec_validSink_23_bits_mask;
  assign sinkVec_queue_23_enq_bits_data = sinkVec_validSink_23_bits_data;
  assign sinkVec_queue_23_enq_bits_last = sinkVec_validSink_23_bits_last;
  assign sinkVec_queue_23_enq_bits_instructionIndex = sinkVec_validSink_23_bits_instructionIndex;
  reg          sinkVec_shifterReg_23_0_valid;
  assign sinkVec_validSink_23_valid = sinkVec_shifterReg_23_0_valid;
  reg  [4:0]   sinkVec_shifterReg_23_0_bits_vd;
  assign sinkVec_validSink_23_bits_vd = sinkVec_shifterReg_23_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_23_0_bits_offset;
  assign sinkVec_validSink_23_bits_offset = sinkVec_shifterReg_23_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_23_0_bits_mask;
  assign sinkVec_validSink_23_bits_mask = sinkVec_shifterReg_23_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_23_0_bits_data;
  assign sinkVec_validSink_23_bits_data = sinkVec_shifterReg_23_0_bits_data;
  reg          sinkVec_shifterReg_23_0_bits_last;
  assign sinkVec_validSink_23_bits_last = sinkVec_shifterReg_23_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_23_0_bits_instructionIndex;
  assign sinkVec_validSink_23_bits_instructionIndex = sinkVec_shifterReg_23_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_23 = sinkVec_shifterReg_23_0_valid | sinkVec_validSource_23_valid;
  assign sinkVec_sinkWire_22_ready = sinkVec_11_0_ready;
  assign sinkVec_sinkWire_23_ready = sinkVec_11_1_ready;
  reg          maskUnitFirst_11;
  wire         tryToRead_11 = sinkVec_11_0_valid | sinkVec_11_1_valid;
  wire         sinkWire_11_valid = maskUnitFirst_11 ? sinkVec_11_0_valid : sinkVec_11_1_valid;
  wire [4:0]   sinkWire_11_bits_vd = maskUnitFirst_11 ? sinkVec_11_0_bits_vd : sinkVec_11_1_bits_vd;
  wire [1:0]   sinkWire_11_bits_offset = maskUnitFirst_11 ? sinkVec_11_0_bits_offset : sinkVec_11_1_bits_offset;
  wire [3:0]   sinkWire_11_bits_mask = maskUnitFirst_11 ? sinkVec_11_0_bits_mask : sinkVec_11_1_bits_mask;
  wire [31:0]  sinkWire_11_bits_data = maskUnitFirst_11 ? sinkVec_11_0_bits_data : sinkVec_11_1_bits_data;
  wire         sinkWire_11_bits_last = maskUnitFirst_11 ? sinkVec_11_0_bits_last : sinkVec_11_1_bits_last;
  wire [2:0]   sinkWire_11_bits_instructionIndex = maskUnitFirst_11 ? sinkVec_11_0_bits_instructionIndex : sinkVec_11_1_bits_instructionIndex;
  wire         sinkWire_11_ready;
  assign sinkVec_11_1_ready = sinkWire_11_ready & ~maskUnitFirst_11;
  assign sinkVec_11_0_ready = sinkWire_11_ready & maskUnitFirst_11;
  reg          view__writeRelease_5_pipe_v;
  wire         view__writeRelease_5_pipe_out_valid = view__writeRelease_5_pipe_v;
  reg          pipe_v_15;
  wire         pipe_out_10_valid = pipe_v_15;
  wire         _probeWire_writeQueueEnqVec_5_valid_T = x22_5_0_ready & _maskUnit_exeResp_5_valid;
  reg          instructionFinishedPipe_pipe_v_5;
  wire         instructionFinishedPipe_pipe_out_5_valid = instructionFinishedPipe_pipe_v_5;
  reg  [7:0]   instructionFinishedPipe_pipe_b_5;
  wire [7:0]   instructionFinishedPipe_pipe_out_5_bits = instructionFinishedPipe_pipe_b_5;
  wire         instructionFinished_5_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_5_bits);
  assign vxsatReportVec_5 = _laneVec_5_vxsatReport[3:0];
  reg          pipe_v_16;
  reg  [31:0]  pipe_b_16;
  reg          pipe_pipe_v_5;
  wire         pipe_pipe_out_5_valid = pipe_pipe_v_5;
  reg  [31:0]  pipe_pipe_b_5;
  wire [31:0]  pipe_pipe_out_5_bits = pipe_pipe_b_5;
  reg          view__laneMaskSelect_5_pipe_v;
  reg  [5:0]   view__laneMaskSelect_5_pipe_b;
  reg          view__laneMaskSelect_5_pipe_pipe_v;
  wire         view__laneMaskSelect_5_pipe_pipe_out_valid = view__laneMaskSelect_5_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_5_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_5_pipe_pipe_out_bits = view__laneMaskSelect_5_pipe_pipe_b;
  reg          view__laneMaskSewSelect_5_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_5_pipe_b;
  reg          view__laneMaskSewSelect_5_pipe_pipe_v;
  wire         view__laneMaskSewSelect_5_pipe_pipe_out_valid = view__laneMaskSewSelect_5_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_5_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_5_pipe_pipe_out_bits = view__laneMaskSewSelect_5_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_5;
  wire         lsuLastPipe_pipe_out_5_valid = lsuLastPipe_pipe_v_5;
  reg  [7:0]   lsuLastPipe_pipe_b_5;
  wire [7:0]   lsuLastPipe_pipe_out_5_bits = lsuLastPipe_pipe_b_5;
  reg          maskLastPipe_pipe_v_5;
  wire         maskLastPipe_pipe_out_5_valid = maskLastPipe_pipe_v_5;
  reg  [7:0]   maskLastPipe_pipe_b_5;
  wire [7:0]   maskLastPipe_pipe_out_5_bits = maskLastPipe_pipe_b_5;
  wire [5:0]   writeCounter_5 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h14};
  reg          pipe_v_17;
  wire         pipe_out_11_valid = pipe_v_17;
  reg  [5:0]   pipe_b_17;
  wire [5:0]   pipe_out_11_bits = pipe_b_17;
  assign laneRequestSinkWire_6_ready = ~laneRequestSinkWire_6_bits_issueInst | _laneVec_6_laneRequest_ready;
  wire         sinkVec_tokenCheck_24;
  wire [4:0]   sinkVec_validSource_24_bits_vs = x13_6_0_bits_vs;
  wire [1:0]   sinkVec_validSource_24_bits_offset = x13_6_0_bits_offset;
  wire [2:0]   sinkVec_validSource_24_bits_instructionIndex = x13_6_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_25;
  wire [4:0]   sinkVec_validSource_25_bits_vs = x13_6_1_bits_vs;
  wire [1:0]   sinkVec_validSource_25_bits_offset = x13_6_1_bits_offset;
  wire [2:0]   sinkVec_validSource_25_bits_instructionIndex = x13_6_1_bits_instructionIndex;
  wire         sinkVec_12_0_ready;
  wire         sinkVec_queue_24_deq_ready = sinkVec_sinkWire_24_ready;
  wire         sinkVec_queue_24_deq_valid;
  wire [4:0]   sinkVec_queue_24_deq_bits_vs;
  wire         sinkVec_12_0_valid = sinkVec_sinkWire_24_valid;
  wire [1:0]   sinkVec_queue_24_deq_bits_readSource;
  wire [4:0]   sinkVec_12_0_bits_vs = sinkVec_sinkWire_24_bits_vs;
  wire [1:0]   sinkVec_queue_24_deq_bits_offset;
  wire [1:0]   sinkVec_12_0_bits_readSource = sinkVec_sinkWire_24_bits_readSource;
  wire [2:0]   sinkVec_queue_24_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_12_0_bits_offset = sinkVec_sinkWire_24_bits_offset;
  wire [2:0]   sinkVec_12_0_bits_instructionIndex = sinkVec_sinkWire_24_bits_instructionIndex;
  wire         sinkVec_validSink_24_valid;
  wire [4:0]   sinkVec_validSink_24_bits_vs;
  wire [1:0]   sinkVec_validSink_24_bits_readSource;
  wire [1:0]   sinkVec_validSink_24_bits_offset;
  wire [2:0]   sinkVec_validSink_24_bits_instructionIndex;
  assign sinkVec_sinkWire_24_valid = sinkVec_queue_24_deq_valid;
  assign sinkVec_sinkWire_24_bits_vs = sinkVec_queue_24_deq_bits_vs;
  assign sinkVec_sinkWire_24_bits_readSource = sinkVec_queue_24_deq_bits_readSource;
  assign sinkVec_sinkWire_24_bits_offset = sinkVec_queue_24_deq_bits_offset;
  assign sinkVec_sinkWire_24_bits_instructionIndex = sinkVec_queue_24_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_24_enq_bits_offset;
  wire [2:0]   sinkVec_queue_24_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_24 = {sinkVec_queue_24_enq_bits_offset, sinkVec_queue_24_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_24_enq_bits_vs;
  wire [1:0]   sinkVec_queue_24_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_24 = {sinkVec_queue_24_enq_bits_vs, sinkVec_queue_24_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_24 = {sinkVec_queue_dataIn_hi_24, sinkVec_queue_dataIn_lo_24};
  wire [2:0]   sinkVec_queue_dataOut_24_instructionIndex = _sinkVec_queue_fifo_24_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_24_offset = _sinkVec_queue_fifo_24_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_24_readSource = _sinkVec_queue_fifo_24_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_24_vs = _sinkVec_queue_fifo_24_data_out[11:7];
  wire         sinkVec_queue_24_enq_ready = ~_sinkVec_queue_fifo_24_full;
  wire         sinkVec_queue_24_enq_valid;
  assign sinkVec_queue_24_deq_valid = ~_sinkVec_queue_fifo_24_empty | sinkVec_queue_24_enq_valid;
  assign sinkVec_queue_24_deq_bits_vs = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_vs : sinkVec_queue_dataOut_24_vs;
  assign sinkVec_queue_24_deq_bits_readSource = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_readSource : sinkVec_queue_dataOut_24_readSource;
  assign sinkVec_queue_24_deq_bits_offset = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_offset : sinkVec_queue_dataOut_24_offset;
  assign sinkVec_queue_24_deq_bits_instructionIndex = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_instructionIndex : sinkVec_queue_dataOut_24_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_24;
  wire         sinkVec_releasePipe_pipe_out_24_valid = sinkVec_releasePipe_pipe_v_24;
  wire         x13_6_0_ready;
  wire         x13_6_0_valid;
  wire         sinkVec_validSource_24_valid = x13_6_0_ready & x13_6_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_24;
  wire [2:0]   sinkVec_tokenCheck_counterChange_24 = sinkVec_validSource_24_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_24 = ~(sinkVec_tokenCheck_counter_24[2]);
  assign x13_6_0_ready = sinkVec_tokenCheck_24;
  assign sinkVec_queue_24_enq_valid = sinkVec_validSink_24_valid;
  assign sinkVec_queue_24_enq_bits_vs = sinkVec_validSink_24_bits_vs;
  assign sinkVec_queue_24_enq_bits_readSource = sinkVec_validSink_24_bits_readSource;
  assign sinkVec_queue_24_enq_bits_offset = sinkVec_validSink_24_bits_offset;
  assign sinkVec_queue_24_enq_bits_instructionIndex = sinkVec_validSink_24_bits_instructionIndex;
  reg          sinkVec_shifterReg_24_0_valid;
  assign sinkVec_validSink_24_valid = sinkVec_shifterReg_24_0_valid;
  reg  [4:0]   sinkVec_shifterReg_24_0_bits_vs;
  assign sinkVec_validSink_24_bits_vs = sinkVec_shifterReg_24_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_24_0_bits_readSource;
  assign sinkVec_validSink_24_bits_readSource = sinkVec_shifterReg_24_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_24_0_bits_offset;
  assign sinkVec_validSink_24_bits_offset = sinkVec_shifterReg_24_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_24_0_bits_instructionIndex;
  assign sinkVec_validSink_24_bits_instructionIndex = sinkVec_shifterReg_24_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_24 = sinkVec_shifterReg_24_0_valid | sinkVec_validSource_24_valid;
  wire         sinkVec_12_1_ready;
  wire         sinkVec_queue_25_deq_ready = sinkVec_sinkWire_25_ready;
  wire         sinkVec_queue_25_deq_valid;
  wire [4:0]   sinkVec_queue_25_deq_bits_vs;
  wire         sinkVec_12_1_valid = sinkVec_sinkWire_25_valid;
  wire [1:0]   sinkVec_queue_25_deq_bits_readSource;
  wire [4:0]   sinkVec_12_1_bits_vs = sinkVec_sinkWire_25_bits_vs;
  wire [1:0]   sinkVec_queue_25_deq_bits_offset;
  wire [1:0]   sinkVec_12_1_bits_readSource = sinkVec_sinkWire_25_bits_readSource;
  wire [2:0]   sinkVec_queue_25_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_12_1_bits_offset = sinkVec_sinkWire_25_bits_offset;
  wire [2:0]   sinkVec_12_1_bits_instructionIndex = sinkVec_sinkWire_25_bits_instructionIndex;
  wire         sinkVec_validSink_25_valid;
  wire [4:0]   sinkVec_validSink_25_bits_vs;
  wire [1:0]   sinkVec_validSink_25_bits_readSource;
  wire [1:0]   sinkVec_validSink_25_bits_offset;
  wire [2:0]   sinkVec_validSink_25_bits_instructionIndex;
  assign sinkVec_sinkWire_25_valid = sinkVec_queue_25_deq_valid;
  assign sinkVec_sinkWire_25_bits_vs = sinkVec_queue_25_deq_bits_vs;
  assign sinkVec_sinkWire_25_bits_readSource = sinkVec_queue_25_deq_bits_readSource;
  assign sinkVec_sinkWire_25_bits_offset = sinkVec_queue_25_deq_bits_offset;
  assign sinkVec_sinkWire_25_bits_instructionIndex = sinkVec_queue_25_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_25_enq_bits_offset;
  wire [2:0]   sinkVec_queue_25_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_25 = {sinkVec_queue_25_enq_bits_offset, sinkVec_queue_25_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_25_enq_bits_vs;
  wire [1:0]   sinkVec_queue_25_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_25 = {sinkVec_queue_25_enq_bits_vs, sinkVec_queue_25_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_25 = {sinkVec_queue_dataIn_hi_25, sinkVec_queue_dataIn_lo_25};
  wire [2:0]   sinkVec_queue_dataOut_25_instructionIndex = _sinkVec_queue_fifo_25_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_25_offset = _sinkVec_queue_fifo_25_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_25_readSource = _sinkVec_queue_fifo_25_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_25_vs = _sinkVec_queue_fifo_25_data_out[11:7];
  wire         sinkVec_queue_25_enq_ready = ~_sinkVec_queue_fifo_25_full;
  wire         sinkVec_queue_25_enq_valid;
  assign sinkVec_queue_25_deq_valid = ~_sinkVec_queue_fifo_25_empty | sinkVec_queue_25_enq_valid;
  assign sinkVec_queue_25_deq_bits_vs = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_vs : sinkVec_queue_dataOut_25_vs;
  assign sinkVec_queue_25_deq_bits_readSource = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_readSource : sinkVec_queue_dataOut_25_readSource;
  assign sinkVec_queue_25_deq_bits_offset = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_offset : sinkVec_queue_dataOut_25_offset;
  assign sinkVec_queue_25_deq_bits_instructionIndex = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_instructionIndex : sinkVec_queue_dataOut_25_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_25;
  wire         sinkVec_releasePipe_pipe_out_25_valid = sinkVec_releasePipe_pipe_v_25;
  wire         x13_6_1_ready;
  wire         x13_6_1_valid;
  wire         sinkVec_validSource_25_valid = x13_6_1_ready & x13_6_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_25;
  wire [2:0]   sinkVec_tokenCheck_counterChange_25 = sinkVec_validSource_25_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_25 = ~(sinkVec_tokenCheck_counter_25[2]);
  assign x13_6_1_ready = sinkVec_tokenCheck_25;
  assign sinkVec_queue_25_enq_valid = sinkVec_validSink_25_valid;
  assign sinkVec_queue_25_enq_bits_vs = sinkVec_validSink_25_bits_vs;
  assign sinkVec_queue_25_enq_bits_readSource = sinkVec_validSink_25_bits_readSource;
  assign sinkVec_queue_25_enq_bits_offset = sinkVec_validSink_25_bits_offset;
  assign sinkVec_queue_25_enq_bits_instructionIndex = sinkVec_validSink_25_bits_instructionIndex;
  reg          sinkVec_shifterReg_25_0_valid;
  assign sinkVec_validSink_25_valid = sinkVec_shifterReg_25_0_valid;
  reg  [4:0]   sinkVec_shifterReg_25_0_bits_vs;
  assign sinkVec_validSink_25_bits_vs = sinkVec_shifterReg_25_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_25_0_bits_readSource;
  assign sinkVec_validSink_25_bits_readSource = sinkVec_shifterReg_25_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_25_0_bits_offset;
  assign sinkVec_validSink_25_bits_offset = sinkVec_shifterReg_25_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_25_0_bits_instructionIndex;
  assign sinkVec_validSink_25_bits_instructionIndex = sinkVec_shifterReg_25_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_25 = sinkVec_shifterReg_25_0_valid | sinkVec_validSource_25_valid;
  assign sinkVec_sinkWire_24_ready = sinkVec_12_0_ready;
  assign sinkVec_sinkWire_25_ready = sinkVec_12_1_ready;
  reg          maskUnitFirst_12;
  wire         tryToRead_12 = sinkVec_12_0_valid | sinkVec_12_1_valid;
  wire         sinkWire_12_valid = maskUnitFirst_12 ? sinkVec_12_0_valid : sinkVec_12_1_valid;
  wire [4:0]   sinkWire_12_bits_vs = maskUnitFirst_12 ? sinkVec_12_0_bits_vs : sinkVec_12_1_bits_vs;
  wire [1:0]   sinkWire_12_bits_readSource = maskUnitFirst_12 ? sinkVec_12_0_bits_readSource : sinkVec_12_1_bits_readSource;
  wire [1:0]   sinkWire_12_bits_offset = maskUnitFirst_12 ? sinkVec_12_0_bits_offset : sinkVec_12_1_bits_offset;
  wire [2:0]   sinkWire_12_bits_instructionIndex = maskUnitFirst_12 ? sinkVec_12_0_bits_instructionIndex : sinkVec_12_1_bits_instructionIndex;
  wire         sinkWire_12_ready;
  assign sinkVec_12_1_ready = sinkWire_12_ready & ~maskUnitFirst_12;
  assign sinkVec_12_0_ready = sinkWire_12_ready & maskUnitFirst_12;
  reg          accessDataValid_pipe_v_12;
  reg          accessDataValid_pipe_pipe_v_12;
  wire         accessDataValid_pipe_pipe_out_12_valid = accessDataValid_pipe_pipe_v_12;
  wire         accessDataSource_12_valid = accessDataValid_pipe_pipe_out_12_valid;
  reg          shifterReg_28_0_valid;
  reg  [31:0]  shifterReg_28_0_bits;
  wire         shifterValid_28 = shifterReg_28_0_valid | accessDataSource_12_valid;
  reg          accessDataValid_pipe_v_13;
  reg          accessDataValid_pipe_pipe_v_13;
  wire         accessDataValid_pipe_pipe_out_13_valid = accessDataValid_pipe_pipe_v_13;
  wire         accessDataSource_13_valid = accessDataValid_pipe_pipe_out_13_valid;
  reg          shifterReg_29_0_valid;
  reg  [31:0]  shifterReg_29_0_bits;
  wire         shifterValid_29 = shifterReg_29_0_valid | accessDataSource_13_valid;
  wire         sinkVec_tokenCheck_26;
  wire [4:0]   sinkVec_validSource_26_bits_vd = x22_6_0_bits_vd;
  wire [1:0]   sinkVec_validSource_26_bits_offset = x22_6_0_bits_offset;
  wire [3:0]   sinkVec_validSource_26_bits_mask = x22_6_0_bits_mask;
  wire [31:0]  sinkVec_validSource_26_bits_data = x22_6_0_bits_data;
  wire [2:0]   sinkVec_validSource_26_bits_instructionIndex = x22_6_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_27;
  wire [4:0]   sinkVec_validSource_27_bits_vd = x22_6_1_bits_vd;
  wire [1:0]   sinkVec_validSource_27_bits_offset = x22_6_1_bits_offset;
  wire [3:0]   sinkVec_validSource_27_bits_mask = x22_6_1_bits_mask;
  wire [31:0]  sinkVec_validSource_27_bits_data = x22_6_1_bits_data;
  wire         sinkVec_validSource_27_bits_last = x22_6_1_bits_last;
  wire [2:0]   sinkVec_validSource_27_bits_instructionIndex = x22_6_1_bits_instructionIndex;
  wire         sinkVec_13_0_ready;
  wire         sinkVec_queue_26_deq_ready = sinkVec_sinkWire_26_ready;
  wire         sinkVec_queue_26_deq_valid;
  wire [4:0]   sinkVec_queue_26_deq_bits_vd;
  wire         sinkVec_13_0_valid = sinkVec_sinkWire_26_valid;
  wire [1:0]   sinkVec_queue_26_deq_bits_offset;
  wire [4:0]   sinkVec_13_0_bits_vd = sinkVec_sinkWire_26_bits_vd;
  wire [3:0]   sinkVec_queue_26_deq_bits_mask;
  wire [1:0]   sinkVec_13_0_bits_offset = sinkVec_sinkWire_26_bits_offset;
  wire [31:0]  sinkVec_queue_26_deq_bits_data;
  wire [3:0]   sinkVec_13_0_bits_mask = sinkVec_sinkWire_26_bits_mask;
  wire         sinkVec_queue_26_deq_bits_last;
  wire [31:0]  sinkVec_13_0_bits_data = sinkVec_sinkWire_26_bits_data;
  wire [2:0]   sinkVec_queue_26_deq_bits_instructionIndex;
  wire         sinkVec_13_0_bits_last = sinkVec_sinkWire_26_bits_last;
  wire [2:0]   sinkVec_13_0_bits_instructionIndex = sinkVec_sinkWire_26_bits_instructionIndex;
  wire         sinkVec_validSink_26_valid;
  wire [4:0]   sinkVec_validSink_26_bits_vd;
  wire [1:0]   sinkVec_validSink_26_bits_offset;
  wire [3:0]   sinkVec_validSink_26_bits_mask;
  wire [31:0]  sinkVec_validSink_26_bits_data;
  wire [2:0]   sinkVec_validSink_26_bits_instructionIndex;
  assign sinkVec_sinkWire_26_valid = sinkVec_queue_26_deq_valid;
  assign sinkVec_sinkWire_26_bits_vd = sinkVec_queue_26_deq_bits_vd;
  assign sinkVec_sinkWire_26_bits_offset = sinkVec_queue_26_deq_bits_offset;
  assign sinkVec_sinkWire_26_bits_mask = sinkVec_queue_26_deq_bits_mask;
  assign sinkVec_sinkWire_26_bits_data = sinkVec_queue_26_deq_bits_data;
  assign sinkVec_sinkWire_26_bits_last = sinkVec_queue_26_deq_bits_last;
  assign sinkVec_sinkWire_26_bits_instructionIndex = sinkVec_queue_26_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_26_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_12 = {sinkVec_queue_26_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_26_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_26 = {sinkVec_queue_dataIn_lo_hi_12, sinkVec_queue_26_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_26_enq_bits_vd;
  wire [1:0]   sinkVec_queue_26_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_12 = {sinkVec_queue_26_enq_bits_vd, sinkVec_queue_26_enq_bits_offset};
  wire [3:0]   sinkVec_queue_26_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_26 = {sinkVec_queue_dataIn_hi_hi_12, sinkVec_queue_26_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_26 = {sinkVec_queue_dataIn_hi_26, sinkVec_queue_dataIn_lo_26};
  wire [2:0]   sinkVec_queue_dataOut_26_instructionIndex = _sinkVec_queue_fifo_26_data_out[2:0];
  wire         sinkVec_queue_dataOut_26_last = _sinkVec_queue_fifo_26_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_26_data = _sinkVec_queue_fifo_26_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_26_mask = _sinkVec_queue_fifo_26_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_26_offset = _sinkVec_queue_fifo_26_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_26_vd = _sinkVec_queue_fifo_26_data_out[46:42];
  wire         sinkVec_queue_26_enq_ready = ~_sinkVec_queue_fifo_26_full;
  wire         sinkVec_queue_26_enq_valid;
  assign sinkVec_queue_26_deq_valid = ~_sinkVec_queue_fifo_26_empty | sinkVec_queue_26_enq_valid;
  assign sinkVec_queue_26_deq_bits_vd = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_vd : sinkVec_queue_dataOut_26_vd;
  assign sinkVec_queue_26_deq_bits_offset = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_offset : sinkVec_queue_dataOut_26_offset;
  assign sinkVec_queue_26_deq_bits_mask = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_mask : sinkVec_queue_dataOut_26_mask;
  assign sinkVec_queue_26_deq_bits_data = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_data : sinkVec_queue_dataOut_26_data;
  assign sinkVec_queue_26_deq_bits_last = ~_sinkVec_queue_fifo_26_empty & sinkVec_queue_dataOut_26_last;
  assign sinkVec_queue_26_deq_bits_instructionIndex = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_instructionIndex : sinkVec_queue_dataOut_26_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_26;
  wire         sinkVec_releasePipe_pipe_out_26_valid = sinkVec_releasePipe_pipe_v_26;
  wire         x22_6_0_ready;
  wire         x22_6_0_valid;
  wire         sinkVec_validSource_26_valid = x22_6_0_ready & x22_6_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_26;
  wire [2:0]   sinkVec_tokenCheck_counterChange_26 = sinkVec_validSource_26_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_26 = ~(sinkVec_tokenCheck_counter_26[2]);
  assign x22_6_0_ready = sinkVec_tokenCheck_26;
  assign sinkVec_queue_26_enq_valid = sinkVec_validSink_26_valid;
  assign sinkVec_queue_26_enq_bits_vd = sinkVec_validSink_26_bits_vd;
  assign sinkVec_queue_26_enq_bits_offset = sinkVec_validSink_26_bits_offset;
  assign sinkVec_queue_26_enq_bits_mask = sinkVec_validSink_26_bits_mask;
  assign sinkVec_queue_26_enq_bits_data = sinkVec_validSink_26_bits_data;
  assign sinkVec_queue_26_enq_bits_instructionIndex = sinkVec_validSink_26_bits_instructionIndex;
  reg          sinkVec_shifterReg_26_0_valid;
  assign sinkVec_validSink_26_valid = sinkVec_shifterReg_26_0_valid;
  reg  [4:0]   sinkVec_shifterReg_26_0_bits_vd;
  assign sinkVec_validSink_26_bits_vd = sinkVec_shifterReg_26_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_26_0_bits_offset;
  assign sinkVec_validSink_26_bits_offset = sinkVec_shifterReg_26_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_26_0_bits_mask;
  assign sinkVec_validSink_26_bits_mask = sinkVec_shifterReg_26_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_26_0_bits_data;
  assign sinkVec_validSink_26_bits_data = sinkVec_shifterReg_26_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_26_0_bits_instructionIndex;
  assign sinkVec_validSink_26_bits_instructionIndex = sinkVec_shifterReg_26_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_26 = sinkVec_shifterReg_26_0_valid | sinkVec_validSource_26_valid;
  wire         sinkVec_13_1_ready;
  wire         sinkVec_queue_27_deq_ready = sinkVec_sinkWire_27_ready;
  wire         sinkVec_queue_27_deq_valid;
  wire [4:0]   sinkVec_queue_27_deq_bits_vd;
  wire         sinkVec_13_1_valid = sinkVec_sinkWire_27_valid;
  wire [1:0]   sinkVec_queue_27_deq_bits_offset;
  wire [4:0]   sinkVec_13_1_bits_vd = sinkVec_sinkWire_27_bits_vd;
  wire [3:0]   sinkVec_queue_27_deq_bits_mask;
  wire [1:0]   sinkVec_13_1_bits_offset = sinkVec_sinkWire_27_bits_offset;
  wire [31:0]  sinkVec_queue_27_deq_bits_data;
  wire [3:0]   sinkVec_13_1_bits_mask = sinkVec_sinkWire_27_bits_mask;
  wire         sinkVec_queue_27_deq_bits_last;
  wire [31:0]  sinkVec_13_1_bits_data = sinkVec_sinkWire_27_bits_data;
  wire [2:0]   sinkVec_queue_27_deq_bits_instructionIndex;
  wire         sinkVec_13_1_bits_last = sinkVec_sinkWire_27_bits_last;
  wire [2:0]   sinkVec_13_1_bits_instructionIndex = sinkVec_sinkWire_27_bits_instructionIndex;
  wire         sinkVec_validSink_27_valid;
  wire [4:0]   sinkVec_validSink_27_bits_vd;
  wire [1:0]   sinkVec_validSink_27_bits_offset;
  wire [3:0]   sinkVec_validSink_27_bits_mask;
  wire [31:0]  sinkVec_validSink_27_bits_data;
  wire         sinkVec_validSink_27_bits_last;
  wire [2:0]   sinkVec_validSink_27_bits_instructionIndex;
  assign sinkVec_sinkWire_27_valid = sinkVec_queue_27_deq_valid;
  assign sinkVec_sinkWire_27_bits_vd = sinkVec_queue_27_deq_bits_vd;
  assign sinkVec_sinkWire_27_bits_offset = sinkVec_queue_27_deq_bits_offset;
  assign sinkVec_sinkWire_27_bits_mask = sinkVec_queue_27_deq_bits_mask;
  assign sinkVec_sinkWire_27_bits_data = sinkVec_queue_27_deq_bits_data;
  assign sinkVec_sinkWire_27_bits_last = sinkVec_queue_27_deq_bits_last;
  assign sinkVec_sinkWire_27_bits_instructionIndex = sinkVec_queue_27_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_27_enq_bits_data;
  wire         sinkVec_queue_27_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_13 = {sinkVec_queue_27_enq_bits_data, sinkVec_queue_27_enq_bits_last};
  wire [2:0]   sinkVec_queue_27_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_27 = {sinkVec_queue_dataIn_lo_hi_13, sinkVec_queue_27_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_27_enq_bits_vd;
  wire [1:0]   sinkVec_queue_27_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_13 = {sinkVec_queue_27_enq_bits_vd, sinkVec_queue_27_enq_bits_offset};
  wire [3:0]   sinkVec_queue_27_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_27 = {sinkVec_queue_dataIn_hi_hi_13, sinkVec_queue_27_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_27 = {sinkVec_queue_dataIn_hi_27, sinkVec_queue_dataIn_lo_27};
  wire [2:0]   sinkVec_queue_dataOut_27_instructionIndex = _sinkVec_queue_fifo_27_data_out[2:0];
  wire         sinkVec_queue_dataOut_27_last = _sinkVec_queue_fifo_27_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_27_data = _sinkVec_queue_fifo_27_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_27_mask = _sinkVec_queue_fifo_27_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_27_offset = _sinkVec_queue_fifo_27_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_27_vd = _sinkVec_queue_fifo_27_data_out[46:42];
  wire         sinkVec_queue_27_enq_ready = ~_sinkVec_queue_fifo_27_full;
  wire         sinkVec_queue_27_enq_valid;
  assign sinkVec_queue_27_deq_valid = ~_sinkVec_queue_fifo_27_empty | sinkVec_queue_27_enq_valid;
  assign sinkVec_queue_27_deq_bits_vd = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_vd : sinkVec_queue_dataOut_27_vd;
  assign sinkVec_queue_27_deq_bits_offset = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_offset : sinkVec_queue_dataOut_27_offset;
  assign sinkVec_queue_27_deq_bits_mask = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_mask : sinkVec_queue_dataOut_27_mask;
  assign sinkVec_queue_27_deq_bits_data = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_data : sinkVec_queue_dataOut_27_data;
  assign sinkVec_queue_27_deq_bits_last = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_last : sinkVec_queue_dataOut_27_last;
  assign sinkVec_queue_27_deq_bits_instructionIndex = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_instructionIndex : sinkVec_queue_dataOut_27_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_27;
  wire         sinkVec_releasePipe_pipe_out_27_valid = sinkVec_releasePipe_pipe_v_27;
  wire         x22_6_1_ready;
  wire         x22_6_1_valid;
  wire         sinkVec_validSource_27_valid = x22_6_1_ready & x22_6_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_27;
  wire [2:0]   sinkVec_tokenCheck_counterChange_27 = sinkVec_validSource_27_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_27 = ~(sinkVec_tokenCheck_counter_27[2]);
  assign x22_6_1_ready = sinkVec_tokenCheck_27;
  assign sinkVec_queue_27_enq_valid = sinkVec_validSink_27_valid;
  assign sinkVec_queue_27_enq_bits_vd = sinkVec_validSink_27_bits_vd;
  assign sinkVec_queue_27_enq_bits_offset = sinkVec_validSink_27_bits_offset;
  assign sinkVec_queue_27_enq_bits_mask = sinkVec_validSink_27_bits_mask;
  assign sinkVec_queue_27_enq_bits_data = sinkVec_validSink_27_bits_data;
  assign sinkVec_queue_27_enq_bits_last = sinkVec_validSink_27_bits_last;
  assign sinkVec_queue_27_enq_bits_instructionIndex = sinkVec_validSink_27_bits_instructionIndex;
  reg          sinkVec_shifterReg_27_0_valid;
  assign sinkVec_validSink_27_valid = sinkVec_shifterReg_27_0_valid;
  reg  [4:0]   sinkVec_shifterReg_27_0_bits_vd;
  assign sinkVec_validSink_27_bits_vd = sinkVec_shifterReg_27_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_27_0_bits_offset;
  assign sinkVec_validSink_27_bits_offset = sinkVec_shifterReg_27_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_27_0_bits_mask;
  assign sinkVec_validSink_27_bits_mask = sinkVec_shifterReg_27_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_27_0_bits_data;
  assign sinkVec_validSink_27_bits_data = sinkVec_shifterReg_27_0_bits_data;
  reg          sinkVec_shifterReg_27_0_bits_last;
  assign sinkVec_validSink_27_bits_last = sinkVec_shifterReg_27_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_27_0_bits_instructionIndex;
  assign sinkVec_validSink_27_bits_instructionIndex = sinkVec_shifterReg_27_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_27 = sinkVec_shifterReg_27_0_valid | sinkVec_validSource_27_valid;
  assign sinkVec_sinkWire_26_ready = sinkVec_13_0_ready;
  assign sinkVec_sinkWire_27_ready = sinkVec_13_1_ready;
  reg          maskUnitFirst_13;
  wire         tryToRead_13 = sinkVec_13_0_valid | sinkVec_13_1_valid;
  wire         sinkWire_13_valid = maskUnitFirst_13 ? sinkVec_13_0_valid : sinkVec_13_1_valid;
  wire [4:0]   sinkWire_13_bits_vd = maskUnitFirst_13 ? sinkVec_13_0_bits_vd : sinkVec_13_1_bits_vd;
  wire [1:0]   sinkWire_13_bits_offset = maskUnitFirst_13 ? sinkVec_13_0_bits_offset : sinkVec_13_1_bits_offset;
  wire [3:0]   sinkWire_13_bits_mask = maskUnitFirst_13 ? sinkVec_13_0_bits_mask : sinkVec_13_1_bits_mask;
  wire [31:0]  sinkWire_13_bits_data = maskUnitFirst_13 ? sinkVec_13_0_bits_data : sinkVec_13_1_bits_data;
  wire         sinkWire_13_bits_last = maskUnitFirst_13 ? sinkVec_13_0_bits_last : sinkVec_13_1_bits_last;
  wire [2:0]   sinkWire_13_bits_instructionIndex = maskUnitFirst_13 ? sinkVec_13_0_bits_instructionIndex : sinkVec_13_1_bits_instructionIndex;
  wire         sinkWire_13_ready;
  assign sinkVec_13_1_ready = sinkWire_13_ready & ~maskUnitFirst_13;
  assign sinkVec_13_0_ready = sinkWire_13_ready & maskUnitFirst_13;
  reg          view__writeRelease_6_pipe_v;
  wire         view__writeRelease_6_pipe_out_valid = view__writeRelease_6_pipe_v;
  reg          pipe_v_18;
  wire         pipe_out_12_valid = pipe_v_18;
  wire         _probeWire_writeQueueEnqVec_6_valid_T = x22_6_0_ready & _maskUnit_exeResp_6_valid;
  reg          instructionFinishedPipe_pipe_v_6;
  wire         instructionFinishedPipe_pipe_out_6_valid = instructionFinishedPipe_pipe_v_6;
  reg  [7:0]   instructionFinishedPipe_pipe_b_6;
  wire [7:0]   instructionFinishedPipe_pipe_out_6_bits = instructionFinishedPipe_pipe_b_6;
  wire         instructionFinished_6_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_6_bits);
  assign vxsatReportVec_6 = _laneVec_6_vxsatReport[3:0];
  reg          pipe_v_19;
  reg  [31:0]  pipe_b_19;
  reg          pipe_pipe_v_6;
  wire         pipe_pipe_out_6_valid = pipe_pipe_v_6;
  reg  [31:0]  pipe_pipe_b_6;
  wire [31:0]  pipe_pipe_out_6_bits = pipe_pipe_b_6;
  reg          view__laneMaskSelect_6_pipe_v;
  reg  [5:0]   view__laneMaskSelect_6_pipe_b;
  reg          view__laneMaskSelect_6_pipe_pipe_v;
  wire         view__laneMaskSelect_6_pipe_pipe_out_valid = view__laneMaskSelect_6_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_6_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_6_pipe_pipe_out_bits = view__laneMaskSelect_6_pipe_pipe_b;
  reg          view__laneMaskSewSelect_6_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_6_pipe_b;
  reg          view__laneMaskSewSelect_6_pipe_pipe_v;
  wire         view__laneMaskSewSelect_6_pipe_pipe_out_valid = view__laneMaskSewSelect_6_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_6_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_6_pipe_pipe_out_bits = view__laneMaskSewSelect_6_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_6;
  wire         lsuLastPipe_pipe_out_6_valid = lsuLastPipe_pipe_v_6;
  reg  [7:0]   lsuLastPipe_pipe_b_6;
  wire [7:0]   lsuLastPipe_pipe_out_6_bits = lsuLastPipe_pipe_b_6;
  reg          maskLastPipe_pipe_v_6;
  wire         maskLastPipe_pipe_out_6_valid = maskLastPipe_pipe_v_6;
  reg  [7:0]   maskLastPipe_pipe_b_6;
  wire [7:0]   maskLastPipe_pipe_out_6_bits = maskLastPipe_pipe_b_6;
  wire [5:0]   writeCounter_6 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h18};
  reg          pipe_v_20;
  wire         pipe_out_13_valid = pipe_v_20;
  reg  [5:0]   pipe_b_20;
  wire [5:0]   pipe_out_13_bits = pipe_b_20;
  assign laneRequestSinkWire_7_ready = ~laneRequestSinkWire_7_bits_issueInst | _laneVec_7_laneRequest_ready;
  wire         sinkVec_tokenCheck_28;
  wire [4:0]   sinkVec_validSource_28_bits_vs = x13_7_0_bits_vs;
  wire [1:0]   sinkVec_validSource_28_bits_offset = x13_7_0_bits_offset;
  wire [2:0]   sinkVec_validSource_28_bits_instructionIndex = x13_7_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_29;
  wire [4:0]   sinkVec_validSource_29_bits_vs = x13_7_1_bits_vs;
  wire [1:0]   sinkVec_validSource_29_bits_offset = x13_7_1_bits_offset;
  wire [2:0]   sinkVec_validSource_29_bits_instructionIndex = x13_7_1_bits_instructionIndex;
  wire         sinkVec_14_0_ready;
  wire         sinkVec_queue_28_deq_ready = sinkVec_sinkWire_28_ready;
  wire         sinkVec_queue_28_deq_valid;
  wire [4:0]   sinkVec_queue_28_deq_bits_vs;
  wire         sinkVec_14_0_valid = sinkVec_sinkWire_28_valid;
  wire [1:0]   sinkVec_queue_28_deq_bits_readSource;
  wire [4:0]   sinkVec_14_0_bits_vs = sinkVec_sinkWire_28_bits_vs;
  wire [1:0]   sinkVec_queue_28_deq_bits_offset;
  wire [1:0]   sinkVec_14_0_bits_readSource = sinkVec_sinkWire_28_bits_readSource;
  wire [2:0]   sinkVec_queue_28_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_14_0_bits_offset = sinkVec_sinkWire_28_bits_offset;
  wire [2:0]   sinkVec_14_0_bits_instructionIndex = sinkVec_sinkWire_28_bits_instructionIndex;
  wire         sinkVec_validSink_28_valid;
  wire [4:0]   sinkVec_validSink_28_bits_vs;
  wire [1:0]   sinkVec_validSink_28_bits_readSource;
  wire [1:0]   sinkVec_validSink_28_bits_offset;
  wire [2:0]   sinkVec_validSink_28_bits_instructionIndex;
  assign sinkVec_sinkWire_28_valid = sinkVec_queue_28_deq_valid;
  assign sinkVec_sinkWire_28_bits_vs = sinkVec_queue_28_deq_bits_vs;
  assign sinkVec_sinkWire_28_bits_readSource = sinkVec_queue_28_deq_bits_readSource;
  assign sinkVec_sinkWire_28_bits_offset = sinkVec_queue_28_deq_bits_offset;
  assign sinkVec_sinkWire_28_bits_instructionIndex = sinkVec_queue_28_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_28_enq_bits_offset;
  wire [2:0]   sinkVec_queue_28_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_28 = {sinkVec_queue_28_enq_bits_offset, sinkVec_queue_28_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_28_enq_bits_vs;
  wire [1:0]   sinkVec_queue_28_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_28 = {sinkVec_queue_28_enq_bits_vs, sinkVec_queue_28_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_28 = {sinkVec_queue_dataIn_hi_28, sinkVec_queue_dataIn_lo_28};
  wire [2:0]   sinkVec_queue_dataOut_28_instructionIndex = _sinkVec_queue_fifo_28_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_28_offset = _sinkVec_queue_fifo_28_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_28_readSource = _sinkVec_queue_fifo_28_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_28_vs = _sinkVec_queue_fifo_28_data_out[11:7];
  wire         sinkVec_queue_28_enq_ready = ~_sinkVec_queue_fifo_28_full;
  wire         sinkVec_queue_28_enq_valid;
  assign sinkVec_queue_28_deq_valid = ~_sinkVec_queue_fifo_28_empty | sinkVec_queue_28_enq_valid;
  assign sinkVec_queue_28_deq_bits_vs = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_vs : sinkVec_queue_dataOut_28_vs;
  assign sinkVec_queue_28_deq_bits_readSource = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_readSource : sinkVec_queue_dataOut_28_readSource;
  assign sinkVec_queue_28_deq_bits_offset = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_offset : sinkVec_queue_dataOut_28_offset;
  assign sinkVec_queue_28_deq_bits_instructionIndex = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_instructionIndex : sinkVec_queue_dataOut_28_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_28;
  wire         sinkVec_releasePipe_pipe_out_28_valid = sinkVec_releasePipe_pipe_v_28;
  wire         x13_7_0_ready;
  wire         x13_7_0_valid;
  wire         sinkVec_validSource_28_valid = x13_7_0_ready & x13_7_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_28;
  wire [2:0]   sinkVec_tokenCheck_counterChange_28 = sinkVec_validSource_28_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_28 = ~(sinkVec_tokenCheck_counter_28[2]);
  assign x13_7_0_ready = sinkVec_tokenCheck_28;
  assign sinkVec_queue_28_enq_valid = sinkVec_validSink_28_valid;
  assign sinkVec_queue_28_enq_bits_vs = sinkVec_validSink_28_bits_vs;
  assign sinkVec_queue_28_enq_bits_readSource = sinkVec_validSink_28_bits_readSource;
  assign sinkVec_queue_28_enq_bits_offset = sinkVec_validSink_28_bits_offset;
  assign sinkVec_queue_28_enq_bits_instructionIndex = sinkVec_validSink_28_bits_instructionIndex;
  reg          sinkVec_shifterReg_28_0_valid;
  assign sinkVec_validSink_28_valid = sinkVec_shifterReg_28_0_valid;
  reg  [4:0]   sinkVec_shifterReg_28_0_bits_vs;
  assign sinkVec_validSink_28_bits_vs = sinkVec_shifterReg_28_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_28_0_bits_readSource;
  assign sinkVec_validSink_28_bits_readSource = sinkVec_shifterReg_28_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_28_0_bits_offset;
  assign sinkVec_validSink_28_bits_offset = sinkVec_shifterReg_28_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_28_0_bits_instructionIndex;
  assign sinkVec_validSink_28_bits_instructionIndex = sinkVec_shifterReg_28_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_28 = sinkVec_shifterReg_28_0_valid | sinkVec_validSource_28_valid;
  wire         sinkVec_14_1_ready;
  wire         sinkVec_queue_29_deq_ready = sinkVec_sinkWire_29_ready;
  wire         sinkVec_queue_29_deq_valid;
  wire [4:0]   sinkVec_queue_29_deq_bits_vs;
  wire         sinkVec_14_1_valid = sinkVec_sinkWire_29_valid;
  wire [1:0]   sinkVec_queue_29_deq_bits_readSource;
  wire [4:0]   sinkVec_14_1_bits_vs = sinkVec_sinkWire_29_bits_vs;
  wire [1:0]   sinkVec_queue_29_deq_bits_offset;
  wire [1:0]   sinkVec_14_1_bits_readSource = sinkVec_sinkWire_29_bits_readSource;
  wire [2:0]   sinkVec_queue_29_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_14_1_bits_offset = sinkVec_sinkWire_29_bits_offset;
  wire [2:0]   sinkVec_14_1_bits_instructionIndex = sinkVec_sinkWire_29_bits_instructionIndex;
  wire         sinkVec_validSink_29_valid;
  wire [4:0]   sinkVec_validSink_29_bits_vs;
  wire [1:0]   sinkVec_validSink_29_bits_readSource;
  wire [1:0]   sinkVec_validSink_29_bits_offset;
  wire [2:0]   sinkVec_validSink_29_bits_instructionIndex;
  assign sinkVec_sinkWire_29_valid = sinkVec_queue_29_deq_valid;
  assign sinkVec_sinkWire_29_bits_vs = sinkVec_queue_29_deq_bits_vs;
  assign sinkVec_sinkWire_29_bits_readSource = sinkVec_queue_29_deq_bits_readSource;
  assign sinkVec_sinkWire_29_bits_offset = sinkVec_queue_29_deq_bits_offset;
  assign sinkVec_sinkWire_29_bits_instructionIndex = sinkVec_queue_29_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_29_enq_bits_offset;
  wire [2:0]   sinkVec_queue_29_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_29 = {sinkVec_queue_29_enq_bits_offset, sinkVec_queue_29_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_29_enq_bits_vs;
  wire [1:0]   sinkVec_queue_29_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_29 = {sinkVec_queue_29_enq_bits_vs, sinkVec_queue_29_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_29 = {sinkVec_queue_dataIn_hi_29, sinkVec_queue_dataIn_lo_29};
  wire [2:0]   sinkVec_queue_dataOut_29_instructionIndex = _sinkVec_queue_fifo_29_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_29_offset = _sinkVec_queue_fifo_29_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_29_readSource = _sinkVec_queue_fifo_29_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_29_vs = _sinkVec_queue_fifo_29_data_out[11:7];
  wire         sinkVec_queue_29_enq_ready = ~_sinkVec_queue_fifo_29_full;
  wire         sinkVec_queue_29_enq_valid;
  assign sinkVec_queue_29_deq_valid = ~_sinkVec_queue_fifo_29_empty | sinkVec_queue_29_enq_valid;
  assign sinkVec_queue_29_deq_bits_vs = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_vs : sinkVec_queue_dataOut_29_vs;
  assign sinkVec_queue_29_deq_bits_readSource = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_readSource : sinkVec_queue_dataOut_29_readSource;
  assign sinkVec_queue_29_deq_bits_offset = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_offset : sinkVec_queue_dataOut_29_offset;
  assign sinkVec_queue_29_deq_bits_instructionIndex = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_instructionIndex : sinkVec_queue_dataOut_29_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_29;
  wire         sinkVec_releasePipe_pipe_out_29_valid = sinkVec_releasePipe_pipe_v_29;
  wire         x13_7_1_ready;
  wire         x13_7_1_valid;
  wire         sinkVec_validSource_29_valid = x13_7_1_ready & x13_7_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_29;
  wire [2:0]   sinkVec_tokenCheck_counterChange_29 = sinkVec_validSource_29_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_29 = ~(sinkVec_tokenCheck_counter_29[2]);
  assign x13_7_1_ready = sinkVec_tokenCheck_29;
  assign sinkVec_queue_29_enq_valid = sinkVec_validSink_29_valid;
  assign sinkVec_queue_29_enq_bits_vs = sinkVec_validSink_29_bits_vs;
  assign sinkVec_queue_29_enq_bits_readSource = sinkVec_validSink_29_bits_readSource;
  assign sinkVec_queue_29_enq_bits_offset = sinkVec_validSink_29_bits_offset;
  assign sinkVec_queue_29_enq_bits_instructionIndex = sinkVec_validSink_29_bits_instructionIndex;
  reg          sinkVec_shifterReg_29_0_valid;
  assign sinkVec_validSink_29_valid = sinkVec_shifterReg_29_0_valid;
  reg  [4:0]   sinkVec_shifterReg_29_0_bits_vs;
  assign sinkVec_validSink_29_bits_vs = sinkVec_shifterReg_29_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_29_0_bits_readSource;
  assign sinkVec_validSink_29_bits_readSource = sinkVec_shifterReg_29_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_29_0_bits_offset;
  assign sinkVec_validSink_29_bits_offset = sinkVec_shifterReg_29_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_29_0_bits_instructionIndex;
  assign sinkVec_validSink_29_bits_instructionIndex = sinkVec_shifterReg_29_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_29 = sinkVec_shifterReg_29_0_valid | sinkVec_validSource_29_valid;
  assign sinkVec_sinkWire_28_ready = sinkVec_14_0_ready;
  assign sinkVec_sinkWire_29_ready = sinkVec_14_1_ready;
  reg          maskUnitFirst_14;
  wire         tryToRead_14 = sinkVec_14_0_valid | sinkVec_14_1_valid;
  wire         sinkWire_14_valid = maskUnitFirst_14 ? sinkVec_14_0_valid : sinkVec_14_1_valid;
  wire [4:0]   sinkWire_14_bits_vs = maskUnitFirst_14 ? sinkVec_14_0_bits_vs : sinkVec_14_1_bits_vs;
  wire [1:0]   sinkWire_14_bits_readSource = maskUnitFirst_14 ? sinkVec_14_0_bits_readSource : sinkVec_14_1_bits_readSource;
  wire [1:0]   sinkWire_14_bits_offset = maskUnitFirst_14 ? sinkVec_14_0_bits_offset : sinkVec_14_1_bits_offset;
  wire [2:0]   sinkWire_14_bits_instructionIndex = maskUnitFirst_14 ? sinkVec_14_0_bits_instructionIndex : sinkVec_14_1_bits_instructionIndex;
  wire         sinkWire_14_ready;
  assign sinkVec_14_1_ready = sinkWire_14_ready & ~maskUnitFirst_14;
  assign sinkVec_14_0_ready = sinkWire_14_ready & maskUnitFirst_14;
  reg          accessDataValid_pipe_v_14;
  reg          accessDataValid_pipe_pipe_v_14;
  wire         accessDataValid_pipe_pipe_out_14_valid = accessDataValid_pipe_pipe_v_14;
  wire         accessDataSource_14_valid = accessDataValid_pipe_pipe_out_14_valid;
  reg          shifterReg_30_0_valid;
  reg  [31:0]  shifterReg_30_0_bits;
  wire         shifterValid_30 = shifterReg_30_0_valid | accessDataSource_14_valid;
  reg          accessDataValid_pipe_v_15;
  reg          accessDataValid_pipe_pipe_v_15;
  wire         accessDataValid_pipe_pipe_out_15_valid = accessDataValid_pipe_pipe_v_15;
  wire         accessDataSource_15_valid = accessDataValid_pipe_pipe_out_15_valid;
  reg          shifterReg_31_0_valid;
  reg  [31:0]  shifterReg_31_0_bits;
  wire         shifterValid_31 = shifterReg_31_0_valid | accessDataSource_15_valid;
  wire         sinkVec_tokenCheck_30;
  wire [4:0]   sinkVec_validSource_30_bits_vd = x22_7_0_bits_vd;
  wire [1:0]   sinkVec_validSource_30_bits_offset = x22_7_0_bits_offset;
  wire [3:0]   sinkVec_validSource_30_bits_mask = x22_7_0_bits_mask;
  wire [31:0]  sinkVec_validSource_30_bits_data = x22_7_0_bits_data;
  wire [2:0]   sinkVec_validSource_30_bits_instructionIndex = x22_7_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_31;
  wire [4:0]   sinkVec_validSource_31_bits_vd = x22_7_1_bits_vd;
  wire [1:0]   sinkVec_validSource_31_bits_offset = x22_7_1_bits_offset;
  wire [3:0]   sinkVec_validSource_31_bits_mask = x22_7_1_bits_mask;
  wire [31:0]  sinkVec_validSource_31_bits_data = x22_7_1_bits_data;
  wire         sinkVec_validSource_31_bits_last = x22_7_1_bits_last;
  wire [2:0]   sinkVec_validSource_31_bits_instructionIndex = x22_7_1_bits_instructionIndex;
  wire         sinkVec_15_0_ready;
  wire         sinkVec_queue_30_deq_ready = sinkVec_sinkWire_30_ready;
  wire         sinkVec_queue_30_deq_valid;
  wire [4:0]   sinkVec_queue_30_deq_bits_vd;
  wire         sinkVec_15_0_valid = sinkVec_sinkWire_30_valid;
  wire [1:0]   sinkVec_queue_30_deq_bits_offset;
  wire [4:0]   sinkVec_15_0_bits_vd = sinkVec_sinkWire_30_bits_vd;
  wire [3:0]   sinkVec_queue_30_deq_bits_mask;
  wire [1:0]   sinkVec_15_0_bits_offset = sinkVec_sinkWire_30_bits_offset;
  wire [31:0]  sinkVec_queue_30_deq_bits_data;
  wire [3:0]   sinkVec_15_0_bits_mask = sinkVec_sinkWire_30_bits_mask;
  wire         sinkVec_queue_30_deq_bits_last;
  wire [31:0]  sinkVec_15_0_bits_data = sinkVec_sinkWire_30_bits_data;
  wire [2:0]   sinkVec_queue_30_deq_bits_instructionIndex;
  wire         sinkVec_15_0_bits_last = sinkVec_sinkWire_30_bits_last;
  wire [2:0]   sinkVec_15_0_bits_instructionIndex = sinkVec_sinkWire_30_bits_instructionIndex;
  wire         sinkVec_validSink_30_valid;
  wire [4:0]   sinkVec_validSink_30_bits_vd;
  wire [1:0]   sinkVec_validSink_30_bits_offset;
  wire [3:0]   sinkVec_validSink_30_bits_mask;
  wire [31:0]  sinkVec_validSink_30_bits_data;
  wire [2:0]   sinkVec_validSink_30_bits_instructionIndex;
  assign sinkVec_sinkWire_30_valid = sinkVec_queue_30_deq_valid;
  assign sinkVec_sinkWire_30_bits_vd = sinkVec_queue_30_deq_bits_vd;
  assign sinkVec_sinkWire_30_bits_offset = sinkVec_queue_30_deq_bits_offset;
  assign sinkVec_sinkWire_30_bits_mask = sinkVec_queue_30_deq_bits_mask;
  assign sinkVec_sinkWire_30_bits_data = sinkVec_queue_30_deq_bits_data;
  assign sinkVec_sinkWire_30_bits_last = sinkVec_queue_30_deq_bits_last;
  assign sinkVec_sinkWire_30_bits_instructionIndex = sinkVec_queue_30_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_30_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_14 = {sinkVec_queue_30_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_30_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_30 = {sinkVec_queue_dataIn_lo_hi_14, sinkVec_queue_30_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_30_enq_bits_vd;
  wire [1:0]   sinkVec_queue_30_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_14 = {sinkVec_queue_30_enq_bits_vd, sinkVec_queue_30_enq_bits_offset};
  wire [3:0]   sinkVec_queue_30_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_30 = {sinkVec_queue_dataIn_hi_hi_14, sinkVec_queue_30_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_30 = {sinkVec_queue_dataIn_hi_30, sinkVec_queue_dataIn_lo_30};
  wire [2:0]   sinkVec_queue_dataOut_30_instructionIndex = _sinkVec_queue_fifo_30_data_out[2:0];
  wire         sinkVec_queue_dataOut_30_last = _sinkVec_queue_fifo_30_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_30_data = _sinkVec_queue_fifo_30_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_30_mask = _sinkVec_queue_fifo_30_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_30_offset = _sinkVec_queue_fifo_30_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_30_vd = _sinkVec_queue_fifo_30_data_out[46:42];
  wire         sinkVec_queue_30_enq_ready = ~_sinkVec_queue_fifo_30_full;
  wire         sinkVec_queue_30_enq_valid;
  assign sinkVec_queue_30_deq_valid = ~_sinkVec_queue_fifo_30_empty | sinkVec_queue_30_enq_valid;
  assign sinkVec_queue_30_deq_bits_vd = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_vd : sinkVec_queue_dataOut_30_vd;
  assign sinkVec_queue_30_deq_bits_offset = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_offset : sinkVec_queue_dataOut_30_offset;
  assign sinkVec_queue_30_deq_bits_mask = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_mask : sinkVec_queue_dataOut_30_mask;
  assign sinkVec_queue_30_deq_bits_data = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_data : sinkVec_queue_dataOut_30_data;
  assign sinkVec_queue_30_deq_bits_last = ~_sinkVec_queue_fifo_30_empty & sinkVec_queue_dataOut_30_last;
  assign sinkVec_queue_30_deq_bits_instructionIndex = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_instructionIndex : sinkVec_queue_dataOut_30_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_30;
  wire         sinkVec_releasePipe_pipe_out_30_valid = sinkVec_releasePipe_pipe_v_30;
  wire         x22_7_0_ready;
  wire         x22_7_0_valid;
  wire         sinkVec_validSource_30_valid = x22_7_0_ready & x22_7_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_30;
  wire [2:0]   sinkVec_tokenCheck_counterChange_30 = sinkVec_validSource_30_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_30 = ~(sinkVec_tokenCheck_counter_30[2]);
  assign x22_7_0_ready = sinkVec_tokenCheck_30;
  assign sinkVec_queue_30_enq_valid = sinkVec_validSink_30_valid;
  assign sinkVec_queue_30_enq_bits_vd = sinkVec_validSink_30_bits_vd;
  assign sinkVec_queue_30_enq_bits_offset = sinkVec_validSink_30_bits_offset;
  assign sinkVec_queue_30_enq_bits_mask = sinkVec_validSink_30_bits_mask;
  assign sinkVec_queue_30_enq_bits_data = sinkVec_validSink_30_bits_data;
  assign sinkVec_queue_30_enq_bits_instructionIndex = sinkVec_validSink_30_bits_instructionIndex;
  reg          sinkVec_shifterReg_30_0_valid;
  assign sinkVec_validSink_30_valid = sinkVec_shifterReg_30_0_valid;
  reg  [4:0]   sinkVec_shifterReg_30_0_bits_vd;
  assign sinkVec_validSink_30_bits_vd = sinkVec_shifterReg_30_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_30_0_bits_offset;
  assign sinkVec_validSink_30_bits_offset = sinkVec_shifterReg_30_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_30_0_bits_mask;
  assign sinkVec_validSink_30_bits_mask = sinkVec_shifterReg_30_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_30_0_bits_data;
  assign sinkVec_validSink_30_bits_data = sinkVec_shifterReg_30_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_30_0_bits_instructionIndex;
  assign sinkVec_validSink_30_bits_instructionIndex = sinkVec_shifterReg_30_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_30 = sinkVec_shifterReg_30_0_valid | sinkVec_validSource_30_valid;
  wire         sinkVec_15_1_ready;
  wire         sinkVec_queue_31_deq_ready = sinkVec_sinkWire_31_ready;
  wire         sinkVec_queue_31_deq_valid;
  wire [4:0]   sinkVec_queue_31_deq_bits_vd;
  wire         sinkVec_15_1_valid = sinkVec_sinkWire_31_valid;
  wire [1:0]   sinkVec_queue_31_deq_bits_offset;
  wire [4:0]   sinkVec_15_1_bits_vd = sinkVec_sinkWire_31_bits_vd;
  wire [3:0]   sinkVec_queue_31_deq_bits_mask;
  wire [1:0]   sinkVec_15_1_bits_offset = sinkVec_sinkWire_31_bits_offset;
  wire [31:0]  sinkVec_queue_31_deq_bits_data;
  wire [3:0]   sinkVec_15_1_bits_mask = sinkVec_sinkWire_31_bits_mask;
  wire         sinkVec_queue_31_deq_bits_last;
  wire [31:0]  sinkVec_15_1_bits_data = sinkVec_sinkWire_31_bits_data;
  wire [2:0]   sinkVec_queue_31_deq_bits_instructionIndex;
  wire         sinkVec_15_1_bits_last = sinkVec_sinkWire_31_bits_last;
  wire [2:0]   sinkVec_15_1_bits_instructionIndex = sinkVec_sinkWire_31_bits_instructionIndex;
  wire         sinkVec_validSink_31_valid;
  wire [4:0]   sinkVec_validSink_31_bits_vd;
  wire [1:0]   sinkVec_validSink_31_bits_offset;
  wire [3:0]   sinkVec_validSink_31_bits_mask;
  wire [31:0]  sinkVec_validSink_31_bits_data;
  wire         sinkVec_validSink_31_bits_last;
  wire [2:0]   sinkVec_validSink_31_bits_instructionIndex;
  assign sinkVec_sinkWire_31_valid = sinkVec_queue_31_deq_valid;
  assign sinkVec_sinkWire_31_bits_vd = sinkVec_queue_31_deq_bits_vd;
  assign sinkVec_sinkWire_31_bits_offset = sinkVec_queue_31_deq_bits_offset;
  assign sinkVec_sinkWire_31_bits_mask = sinkVec_queue_31_deq_bits_mask;
  assign sinkVec_sinkWire_31_bits_data = sinkVec_queue_31_deq_bits_data;
  assign sinkVec_sinkWire_31_bits_last = sinkVec_queue_31_deq_bits_last;
  assign sinkVec_sinkWire_31_bits_instructionIndex = sinkVec_queue_31_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_31_enq_bits_data;
  wire         sinkVec_queue_31_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_15 = {sinkVec_queue_31_enq_bits_data, sinkVec_queue_31_enq_bits_last};
  wire [2:0]   sinkVec_queue_31_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_31 = {sinkVec_queue_dataIn_lo_hi_15, sinkVec_queue_31_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_31_enq_bits_vd;
  wire [1:0]   sinkVec_queue_31_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_15 = {sinkVec_queue_31_enq_bits_vd, sinkVec_queue_31_enq_bits_offset};
  wire [3:0]   sinkVec_queue_31_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_31 = {sinkVec_queue_dataIn_hi_hi_15, sinkVec_queue_31_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_31 = {sinkVec_queue_dataIn_hi_31, sinkVec_queue_dataIn_lo_31};
  wire [2:0]   sinkVec_queue_dataOut_31_instructionIndex = _sinkVec_queue_fifo_31_data_out[2:0];
  wire         sinkVec_queue_dataOut_31_last = _sinkVec_queue_fifo_31_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_31_data = _sinkVec_queue_fifo_31_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_31_mask = _sinkVec_queue_fifo_31_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_31_offset = _sinkVec_queue_fifo_31_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_31_vd = _sinkVec_queue_fifo_31_data_out[46:42];
  wire         sinkVec_queue_31_enq_ready = ~_sinkVec_queue_fifo_31_full;
  wire         sinkVec_queue_31_enq_valid;
  assign sinkVec_queue_31_deq_valid = ~_sinkVec_queue_fifo_31_empty | sinkVec_queue_31_enq_valid;
  assign sinkVec_queue_31_deq_bits_vd = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_vd : sinkVec_queue_dataOut_31_vd;
  assign sinkVec_queue_31_deq_bits_offset = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_offset : sinkVec_queue_dataOut_31_offset;
  assign sinkVec_queue_31_deq_bits_mask = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_mask : sinkVec_queue_dataOut_31_mask;
  assign sinkVec_queue_31_deq_bits_data = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_data : sinkVec_queue_dataOut_31_data;
  assign sinkVec_queue_31_deq_bits_last = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_last : sinkVec_queue_dataOut_31_last;
  assign sinkVec_queue_31_deq_bits_instructionIndex = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_instructionIndex : sinkVec_queue_dataOut_31_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_31;
  wire         sinkVec_releasePipe_pipe_out_31_valid = sinkVec_releasePipe_pipe_v_31;
  wire         x22_7_1_ready;
  wire         x22_7_1_valid;
  wire         sinkVec_validSource_31_valid = x22_7_1_ready & x22_7_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_31;
  wire [2:0]   sinkVec_tokenCheck_counterChange_31 = sinkVec_validSource_31_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_31 = ~(sinkVec_tokenCheck_counter_31[2]);
  assign x22_7_1_ready = sinkVec_tokenCheck_31;
  assign sinkVec_queue_31_enq_valid = sinkVec_validSink_31_valid;
  assign sinkVec_queue_31_enq_bits_vd = sinkVec_validSink_31_bits_vd;
  assign sinkVec_queue_31_enq_bits_offset = sinkVec_validSink_31_bits_offset;
  assign sinkVec_queue_31_enq_bits_mask = sinkVec_validSink_31_bits_mask;
  assign sinkVec_queue_31_enq_bits_data = sinkVec_validSink_31_bits_data;
  assign sinkVec_queue_31_enq_bits_last = sinkVec_validSink_31_bits_last;
  assign sinkVec_queue_31_enq_bits_instructionIndex = sinkVec_validSink_31_bits_instructionIndex;
  reg          sinkVec_shifterReg_31_0_valid;
  assign sinkVec_validSink_31_valid = sinkVec_shifterReg_31_0_valid;
  reg  [4:0]   sinkVec_shifterReg_31_0_bits_vd;
  assign sinkVec_validSink_31_bits_vd = sinkVec_shifterReg_31_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_31_0_bits_offset;
  assign sinkVec_validSink_31_bits_offset = sinkVec_shifterReg_31_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_31_0_bits_mask;
  assign sinkVec_validSink_31_bits_mask = sinkVec_shifterReg_31_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_31_0_bits_data;
  assign sinkVec_validSink_31_bits_data = sinkVec_shifterReg_31_0_bits_data;
  reg          sinkVec_shifterReg_31_0_bits_last;
  assign sinkVec_validSink_31_bits_last = sinkVec_shifterReg_31_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_31_0_bits_instructionIndex;
  assign sinkVec_validSink_31_bits_instructionIndex = sinkVec_shifterReg_31_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_31 = sinkVec_shifterReg_31_0_valid | sinkVec_validSource_31_valid;
  assign sinkVec_sinkWire_30_ready = sinkVec_15_0_ready;
  assign sinkVec_sinkWire_31_ready = sinkVec_15_1_ready;
  reg          maskUnitFirst_15;
  wire         tryToRead_15 = sinkVec_15_0_valid | sinkVec_15_1_valid;
  wire         sinkWire_15_valid = maskUnitFirst_15 ? sinkVec_15_0_valid : sinkVec_15_1_valid;
  wire [4:0]   sinkWire_15_bits_vd = maskUnitFirst_15 ? sinkVec_15_0_bits_vd : sinkVec_15_1_bits_vd;
  wire [1:0]   sinkWire_15_bits_offset = maskUnitFirst_15 ? sinkVec_15_0_bits_offset : sinkVec_15_1_bits_offset;
  wire [3:0]   sinkWire_15_bits_mask = maskUnitFirst_15 ? sinkVec_15_0_bits_mask : sinkVec_15_1_bits_mask;
  wire [31:0]  sinkWire_15_bits_data = maskUnitFirst_15 ? sinkVec_15_0_bits_data : sinkVec_15_1_bits_data;
  wire         sinkWire_15_bits_last = maskUnitFirst_15 ? sinkVec_15_0_bits_last : sinkVec_15_1_bits_last;
  wire [2:0]   sinkWire_15_bits_instructionIndex = maskUnitFirst_15 ? sinkVec_15_0_bits_instructionIndex : sinkVec_15_1_bits_instructionIndex;
  wire         sinkWire_15_ready;
  assign sinkVec_15_1_ready = sinkWire_15_ready & ~maskUnitFirst_15;
  assign sinkVec_15_0_ready = sinkWire_15_ready & maskUnitFirst_15;
  reg          view__writeRelease_7_pipe_v;
  wire         view__writeRelease_7_pipe_out_valid = view__writeRelease_7_pipe_v;
  reg          pipe_v_21;
  wire         pipe_out_14_valid = pipe_v_21;
  wire         _probeWire_writeQueueEnqVec_7_valid_T = x22_7_0_ready & _maskUnit_exeResp_7_valid;
  reg          instructionFinishedPipe_pipe_v_7;
  wire         instructionFinishedPipe_pipe_out_7_valid = instructionFinishedPipe_pipe_v_7;
  reg  [7:0]   instructionFinishedPipe_pipe_b_7;
  wire [7:0]   instructionFinishedPipe_pipe_out_7_bits = instructionFinishedPipe_pipe_b_7;
  wire         instructionFinished_7_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_7_bits);
  assign vxsatReportVec_7 = _laneVec_7_vxsatReport[3:0];
  reg          pipe_v_22;
  reg  [31:0]  pipe_b_22;
  reg          pipe_pipe_v_7;
  wire         pipe_pipe_out_7_valid = pipe_pipe_v_7;
  reg  [31:0]  pipe_pipe_b_7;
  wire [31:0]  pipe_pipe_out_7_bits = pipe_pipe_b_7;
  reg          view__laneMaskSelect_7_pipe_v;
  reg  [5:0]   view__laneMaskSelect_7_pipe_b;
  reg          view__laneMaskSelect_7_pipe_pipe_v;
  wire         view__laneMaskSelect_7_pipe_pipe_out_valid = view__laneMaskSelect_7_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_7_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_7_pipe_pipe_out_bits = view__laneMaskSelect_7_pipe_pipe_b;
  reg          view__laneMaskSewSelect_7_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_7_pipe_b;
  reg          view__laneMaskSewSelect_7_pipe_pipe_v;
  wire         view__laneMaskSewSelect_7_pipe_pipe_out_valid = view__laneMaskSewSelect_7_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_7_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_7_pipe_pipe_out_bits = view__laneMaskSewSelect_7_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_7;
  wire         lsuLastPipe_pipe_out_7_valid = lsuLastPipe_pipe_v_7;
  reg  [7:0]   lsuLastPipe_pipe_b_7;
  wire [7:0]   lsuLastPipe_pipe_out_7_bits = lsuLastPipe_pipe_b_7;
  reg          maskLastPipe_pipe_v_7;
  wire         maskLastPipe_pipe_out_7_valid = maskLastPipe_pipe_v_7;
  reg  [7:0]   maskLastPipe_pipe_b_7;
  wire [7:0]   maskLastPipe_pipe_out_7_bits = maskLastPipe_pipe_b_7;
  wire [5:0]   writeCounter_7 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h1C};
  reg          pipe_v_23;
  wire         pipe_out_15_valid = pipe_v_23;
  reg  [5:0]   pipe_b_23;
  wire [5:0]   pipe_out_15_bits = pipe_b_23;
  assign laneRequestSinkWire_8_ready = ~laneRequestSinkWire_8_bits_issueInst | _laneVec_8_laneRequest_ready;
  wire         sinkVec_tokenCheck_32;
  wire [4:0]   sinkVec_validSource_32_bits_vs = x13_8_0_bits_vs;
  wire [1:0]   sinkVec_validSource_32_bits_offset = x13_8_0_bits_offset;
  wire [2:0]   sinkVec_validSource_32_bits_instructionIndex = x13_8_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_33;
  wire [4:0]   sinkVec_validSource_33_bits_vs = x13_8_1_bits_vs;
  wire [1:0]   sinkVec_validSource_33_bits_offset = x13_8_1_bits_offset;
  wire [2:0]   sinkVec_validSource_33_bits_instructionIndex = x13_8_1_bits_instructionIndex;
  wire         sinkVec_16_0_ready;
  wire         sinkVec_queue_32_deq_ready = sinkVec_sinkWire_32_ready;
  wire         sinkVec_queue_32_deq_valid;
  wire [4:0]   sinkVec_queue_32_deq_bits_vs;
  wire         sinkVec_16_0_valid = sinkVec_sinkWire_32_valid;
  wire [1:0]   sinkVec_queue_32_deq_bits_readSource;
  wire [4:0]   sinkVec_16_0_bits_vs = sinkVec_sinkWire_32_bits_vs;
  wire [1:0]   sinkVec_queue_32_deq_bits_offset;
  wire [1:0]   sinkVec_16_0_bits_readSource = sinkVec_sinkWire_32_bits_readSource;
  wire [2:0]   sinkVec_queue_32_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_16_0_bits_offset = sinkVec_sinkWire_32_bits_offset;
  wire [2:0]   sinkVec_16_0_bits_instructionIndex = sinkVec_sinkWire_32_bits_instructionIndex;
  wire         sinkVec_validSink_32_valid;
  wire [4:0]   sinkVec_validSink_32_bits_vs;
  wire [1:0]   sinkVec_validSink_32_bits_readSource;
  wire [1:0]   sinkVec_validSink_32_bits_offset;
  wire [2:0]   sinkVec_validSink_32_bits_instructionIndex;
  assign sinkVec_sinkWire_32_valid = sinkVec_queue_32_deq_valid;
  assign sinkVec_sinkWire_32_bits_vs = sinkVec_queue_32_deq_bits_vs;
  assign sinkVec_sinkWire_32_bits_readSource = sinkVec_queue_32_deq_bits_readSource;
  assign sinkVec_sinkWire_32_bits_offset = sinkVec_queue_32_deq_bits_offset;
  assign sinkVec_sinkWire_32_bits_instructionIndex = sinkVec_queue_32_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_32_enq_bits_offset;
  wire [2:0]   sinkVec_queue_32_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_32 = {sinkVec_queue_32_enq_bits_offset, sinkVec_queue_32_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_32_enq_bits_vs;
  wire [1:0]   sinkVec_queue_32_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_32 = {sinkVec_queue_32_enq_bits_vs, sinkVec_queue_32_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_32 = {sinkVec_queue_dataIn_hi_32, sinkVec_queue_dataIn_lo_32};
  wire [2:0]   sinkVec_queue_dataOut_32_instructionIndex = _sinkVec_queue_fifo_32_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_32_offset = _sinkVec_queue_fifo_32_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_32_readSource = _sinkVec_queue_fifo_32_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_32_vs = _sinkVec_queue_fifo_32_data_out[11:7];
  wire         sinkVec_queue_32_enq_ready = ~_sinkVec_queue_fifo_32_full;
  wire         sinkVec_queue_32_enq_valid;
  assign sinkVec_queue_32_deq_valid = ~_sinkVec_queue_fifo_32_empty | sinkVec_queue_32_enq_valid;
  assign sinkVec_queue_32_deq_bits_vs = _sinkVec_queue_fifo_32_empty ? sinkVec_queue_32_enq_bits_vs : sinkVec_queue_dataOut_32_vs;
  assign sinkVec_queue_32_deq_bits_readSource = _sinkVec_queue_fifo_32_empty ? sinkVec_queue_32_enq_bits_readSource : sinkVec_queue_dataOut_32_readSource;
  assign sinkVec_queue_32_deq_bits_offset = _sinkVec_queue_fifo_32_empty ? sinkVec_queue_32_enq_bits_offset : sinkVec_queue_dataOut_32_offset;
  assign sinkVec_queue_32_deq_bits_instructionIndex = _sinkVec_queue_fifo_32_empty ? sinkVec_queue_32_enq_bits_instructionIndex : sinkVec_queue_dataOut_32_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_32;
  wire         sinkVec_releasePipe_pipe_out_32_valid = sinkVec_releasePipe_pipe_v_32;
  wire         x13_8_0_ready;
  wire         x13_8_0_valid;
  wire         sinkVec_validSource_32_valid = x13_8_0_ready & x13_8_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_32;
  wire [2:0]   sinkVec_tokenCheck_counterChange_32 = sinkVec_validSource_32_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_32 = ~(sinkVec_tokenCheck_counter_32[2]);
  assign x13_8_0_ready = sinkVec_tokenCheck_32;
  assign sinkVec_queue_32_enq_valid = sinkVec_validSink_32_valid;
  assign sinkVec_queue_32_enq_bits_vs = sinkVec_validSink_32_bits_vs;
  assign sinkVec_queue_32_enq_bits_readSource = sinkVec_validSink_32_bits_readSource;
  assign sinkVec_queue_32_enq_bits_offset = sinkVec_validSink_32_bits_offset;
  assign sinkVec_queue_32_enq_bits_instructionIndex = sinkVec_validSink_32_bits_instructionIndex;
  reg          sinkVec_shifterReg_32_0_valid;
  assign sinkVec_validSink_32_valid = sinkVec_shifterReg_32_0_valid;
  reg  [4:0]   sinkVec_shifterReg_32_0_bits_vs;
  assign sinkVec_validSink_32_bits_vs = sinkVec_shifterReg_32_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_32_0_bits_readSource;
  assign sinkVec_validSink_32_bits_readSource = sinkVec_shifterReg_32_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_32_0_bits_offset;
  assign sinkVec_validSink_32_bits_offset = sinkVec_shifterReg_32_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_32_0_bits_instructionIndex;
  assign sinkVec_validSink_32_bits_instructionIndex = sinkVec_shifterReg_32_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_32 = sinkVec_shifterReg_32_0_valid | sinkVec_validSource_32_valid;
  wire         sinkVec_16_1_ready;
  wire         sinkVec_queue_33_deq_ready = sinkVec_sinkWire_33_ready;
  wire         sinkVec_queue_33_deq_valid;
  wire [4:0]   sinkVec_queue_33_deq_bits_vs;
  wire         sinkVec_16_1_valid = sinkVec_sinkWire_33_valid;
  wire [1:0]   sinkVec_queue_33_deq_bits_readSource;
  wire [4:0]   sinkVec_16_1_bits_vs = sinkVec_sinkWire_33_bits_vs;
  wire [1:0]   sinkVec_queue_33_deq_bits_offset;
  wire [1:0]   sinkVec_16_1_bits_readSource = sinkVec_sinkWire_33_bits_readSource;
  wire [2:0]   sinkVec_queue_33_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_16_1_bits_offset = sinkVec_sinkWire_33_bits_offset;
  wire [2:0]   sinkVec_16_1_bits_instructionIndex = sinkVec_sinkWire_33_bits_instructionIndex;
  wire         sinkVec_validSink_33_valid;
  wire [4:0]   sinkVec_validSink_33_bits_vs;
  wire [1:0]   sinkVec_validSink_33_bits_readSource;
  wire [1:0]   sinkVec_validSink_33_bits_offset;
  wire [2:0]   sinkVec_validSink_33_bits_instructionIndex;
  assign sinkVec_sinkWire_33_valid = sinkVec_queue_33_deq_valid;
  assign sinkVec_sinkWire_33_bits_vs = sinkVec_queue_33_deq_bits_vs;
  assign sinkVec_sinkWire_33_bits_readSource = sinkVec_queue_33_deq_bits_readSource;
  assign sinkVec_sinkWire_33_bits_offset = sinkVec_queue_33_deq_bits_offset;
  assign sinkVec_sinkWire_33_bits_instructionIndex = sinkVec_queue_33_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_33_enq_bits_offset;
  wire [2:0]   sinkVec_queue_33_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_33 = {sinkVec_queue_33_enq_bits_offset, sinkVec_queue_33_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_33_enq_bits_vs;
  wire [1:0]   sinkVec_queue_33_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_33 = {sinkVec_queue_33_enq_bits_vs, sinkVec_queue_33_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_33 = {sinkVec_queue_dataIn_hi_33, sinkVec_queue_dataIn_lo_33};
  wire [2:0]   sinkVec_queue_dataOut_33_instructionIndex = _sinkVec_queue_fifo_33_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_33_offset = _sinkVec_queue_fifo_33_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_33_readSource = _sinkVec_queue_fifo_33_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_33_vs = _sinkVec_queue_fifo_33_data_out[11:7];
  wire         sinkVec_queue_33_enq_ready = ~_sinkVec_queue_fifo_33_full;
  wire         sinkVec_queue_33_enq_valid;
  assign sinkVec_queue_33_deq_valid = ~_sinkVec_queue_fifo_33_empty | sinkVec_queue_33_enq_valid;
  assign sinkVec_queue_33_deq_bits_vs = _sinkVec_queue_fifo_33_empty ? sinkVec_queue_33_enq_bits_vs : sinkVec_queue_dataOut_33_vs;
  assign sinkVec_queue_33_deq_bits_readSource = _sinkVec_queue_fifo_33_empty ? sinkVec_queue_33_enq_bits_readSource : sinkVec_queue_dataOut_33_readSource;
  assign sinkVec_queue_33_deq_bits_offset = _sinkVec_queue_fifo_33_empty ? sinkVec_queue_33_enq_bits_offset : sinkVec_queue_dataOut_33_offset;
  assign sinkVec_queue_33_deq_bits_instructionIndex = _sinkVec_queue_fifo_33_empty ? sinkVec_queue_33_enq_bits_instructionIndex : sinkVec_queue_dataOut_33_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_33;
  wire         sinkVec_releasePipe_pipe_out_33_valid = sinkVec_releasePipe_pipe_v_33;
  wire         x13_8_1_ready;
  wire         x13_8_1_valid;
  wire         sinkVec_validSource_33_valid = x13_8_1_ready & x13_8_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_33;
  wire [2:0]   sinkVec_tokenCheck_counterChange_33 = sinkVec_validSource_33_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_33 = ~(sinkVec_tokenCheck_counter_33[2]);
  assign x13_8_1_ready = sinkVec_tokenCheck_33;
  assign sinkVec_queue_33_enq_valid = sinkVec_validSink_33_valid;
  assign sinkVec_queue_33_enq_bits_vs = sinkVec_validSink_33_bits_vs;
  assign sinkVec_queue_33_enq_bits_readSource = sinkVec_validSink_33_bits_readSource;
  assign sinkVec_queue_33_enq_bits_offset = sinkVec_validSink_33_bits_offset;
  assign sinkVec_queue_33_enq_bits_instructionIndex = sinkVec_validSink_33_bits_instructionIndex;
  reg          sinkVec_shifterReg_33_0_valid;
  assign sinkVec_validSink_33_valid = sinkVec_shifterReg_33_0_valid;
  reg  [4:0]   sinkVec_shifterReg_33_0_bits_vs;
  assign sinkVec_validSink_33_bits_vs = sinkVec_shifterReg_33_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_33_0_bits_readSource;
  assign sinkVec_validSink_33_bits_readSource = sinkVec_shifterReg_33_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_33_0_bits_offset;
  assign sinkVec_validSink_33_bits_offset = sinkVec_shifterReg_33_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_33_0_bits_instructionIndex;
  assign sinkVec_validSink_33_bits_instructionIndex = sinkVec_shifterReg_33_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_33 = sinkVec_shifterReg_33_0_valid | sinkVec_validSource_33_valid;
  assign sinkVec_sinkWire_32_ready = sinkVec_16_0_ready;
  assign sinkVec_sinkWire_33_ready = sinkVec_16_1_ready;
  reg          maskUnitFirst_16;
  wire         tryToRead_16 = sinkVec_16_0_valid | sinkVec_16_1_valid;
  wire         sinkWire_16_valid = maskUnitFirst_16 ? sinkVec_16_0_valid : sinkVec_16_1_valid;
  wire [4:0]   sinkWire_16_bits_vs = maskUnitFirst_16 ? sinkVec_16_0_bits_vs : sinkVec_16_1_bits_vs;
  wire [1:0]   sinkWire_16_bits_readSource = maskUnitFirst_16 ? sinkVec_16_0_bits_readSource : sinkVec_16_1_bits_readSource;
  wire [1:0]   sinkWire_16_bits_offset = maskUnitFirst_16 ? sinkVec_16_0_bits_offset : sinkVec_16_1_bits_offset;
  wire [2:0]   sinkWire_16_bits_instructionIndex = maskUnitFirst_16 ? sinkVec_16_0_bits_instructionIndex : sinkVec_16_1_bits_instructionIndex;
  wire         sinkWire_16_ready;
  assign sinkVec_16_1_ready = sinkWire_16_ready & ~maskUnitFirst_16;
  assign sinkVec_16_0_ready = sinkWire_16_ready & maskUnitFirst_16;
  reg          accessDataValid_pipe_v_16;
  reg          accessDataValid_pipe_pipe_v_16;
  wire         accessDataValid_pipe_pipe_out_16_valid = accessDataValid_pipe_pipe_v_16;
  wire         accessDataSource_16_valid = accessDataValid_pipe_pipe_out_16_valid;
  reg          shifterReg_32_0_valid;
  reg  [31:0]  shifterReg_32_0_bits;
  wire         shifterValid_32 = shifterReg_32_0_valid | accessDataSource_16_valid;
  reg          accessDataValid_pipe_v_17;
  reg          accessDataValid_pipe_pipe_v_17;
  wire         accessDataValid_pipe_pipe_out_17_valid = accessDataValid_pipe_pipe_v_17;
  wire         accessDataSource_17_valid = accessDataValid_pipe_pipe_out_17_valid;
  reg          shifterReg_33_0_valid;
  reg  [31:0]  shifterReg_33_0_bits;
  wire         shifterValid_33 = shifterReg_33_0_valid | accessDataSource_17_valid;
  wire         sinkVec_tokenCheck_34;
  wire [4:0]   sinkVec_validSource_34_bits_vd = x22_8_0_bits_vd;
  wire [1:0]   sinkVec_validSource_34_bits_offset = x22_8_0_bits_offset;
  wire [3:0]   sinkVec_validSource_34_bits_mask = x22_8_0_bits_mask;
  wire [31:0]  sinkVec_validSource_34_bits_data = x22_8_0_bits_data;
  wire [2:0]   sinkVec_validSource_34_bits_instructionIndex = x22_8_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_35;
  wire [4:0]   sinkVec_validSource_35_bits_vd = x22_8_1_bits_vd;
  wire [1:0]   sinkVec_validSource_35_bits_offset = x22_8_1_bits_offset;
  wire [3:0]   sinkVec_validSource_35_bits_mask = x22_8_1_bits_mask;
  wire [31:0]  sinkVec_validSource_35_bits_data = x22_8_1_bits_data;
  wire         sinkVec_validSource_35_bits_last = x22_8_1_bits_last;
  wire [2:0]   sinkVec_validSource_35_bits_instructionIndex = x22_8_1_bits_instructionIndex;
  wire         sinkVec_17_0_ready;
  wire         sinkVec_queue_34_deq_ready = sinkVec_sinkWire_34_ready;
  wire         sinkVec_queue_34_deq_valid;
  wire [4:0]   sinkVec_queue_34_deq_bits_vd;
  wire         sinkVec_17_0_valid = sinkVec_sinkWire_34_valid;
  wire [1:0]   sinkVec_queue_34_deq_bits_offset;
  wire [4:0]   sinkVec_17_0_bits_vd = sinkVec_sinkWire_34_bits_vd;
  wire [3:0]   sinkVec_queue_34_deq_bits_mask;
  wire [1:0]   sinkVec_17_0_bits_offset = sinkVec_sinkWire_34_bits_offset;
  wire [31:0]  sinkVec_queue_34_deq_bits_data;
  wire [3:0]   sinkVec_17_0_bits_mask = sinkVec_sinkWire_34_bits_mask;
  wire         sinkVec_queue_34_deq_bits_last;
  wire [31:0]  sinkVec_17_0_bits_data = sinkVec_sinkWire_34_bits_data;
  wire [2:0]   sinkVec_queue_34_deq_bits_instructionIndex;
  wire         sinkVec_17_0_bits_last = sinkVec_sinkWire_34_bits_last;
  wire [2:0]   sinkVec_17_0_bits_instructionIndex = sinkVec_sinkWire_34_bits_instructionIndex;
  wire         sinkVec_validSink_34_valid;
  wire [4:0]   sinkVec_validSink_34_bits_vd;
  wire [1:0]   sinkVec_validSink_34_bits_offset;
  wire [3:0]   sinkVec_validSink_34_bits_mask;
  wire [31:0]  sinkVec_validSink_34_bits_data;
  wire [2:0]   sinkVec_validSink_34_bits_instructionIndex;
  assign sinkVec_sinkWire_34_valid = sinkVec_queue_34_deq_valid;
  assign sinkVec_sinkWire_34_bits_vd = sinkVec_queue_34_deq_bits_vd;
  assign sinkVec_sinkWire_34_bits_offset = sinkVec_queue_34_deq_bits_offset;
  assign sinkVec_sinkWire_34_bits_mask = sinkVec_queue_34_deq_bits_mask;
  assign sinkVec_sinkWire_34_bits_data = sinkVec_queue_34_deq_bits_data;
  assign sinkVec_sinkWire_34_bits_last = sinkVec_queue_34_deq_bits_last;
  assign sinkVec_sinkWire_34_bits_instructionIndex = sinkVec_queue_34_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_34_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_16 = {sinkVec_queue_34_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_34_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_34 = {sinkVec_queue_dataIn_lo_hi_16, sinkVec_queue_34_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_34_enq_bits_vd;
  wire [1:0]   sinkVec_queue_34_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_16 = {sinkVec_queue_34_enq_bits_vd, sinkVec_queue_34_enq_bits_offset};
  wire [3:0]   sinkVec_queue_34_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_34 = {sinkVec_queue_dataIn_hi_hi_16, sinkVec_queue_34_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_34 = {sinkVec_queue_dataIn_hi_34, sinkVec_queue_dataIn_lo_34};
  wire [2:0]   sinkVec_queue_dataOut_34_instructionIndex = _sinkVec_queue_fifo_34_data_out[2:0];
  wire         sinkVec_queue_dataOut_34_last = _sinkVec_queue_fifo_34_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_34_data = _sinkVec_queue_fifo_34_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_34_mask = _sinkVec_queue_fifo_34_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_34_offset = _sinkVec_queue_fifo_34_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_34_vd = _sinkVec_queue_fifo_34_data_out[46:42];
  wire         sinkVec_queue_34_enq_ready = ~_sinkVec_queue_fifo_34_full;
  wire         sinkVec_queue_34_enq_valid;
  assign sinkVec_queue_34_deq_valid = ~_sinkVec_queue_fifo_34_empty | sinkVec_queue_34_enq_valid;
  assign sinkVec_queue_34_deq_bits_vd = _sinkVec_queue_fifo_34_empty ? sinkVec_queue_34_enq_bits_vd : sinkVec_queue_dataOut_34_vd;
  assign sinkVec_queue_34_deq_bits_offset = _sinkVec_queue_fifo_34_empty ? sinkVec_queue_34_enq_bits_offset : sinkVec_queue_dataOut_34_offset;
  assign sinkVec_queue_34_deq_bits_mask = _sinkVec_queue_fifo_34_empty ? sinkVec_queue_34_enq_bits_mask : sinkVec_queue_dataOut_34_mask;
  assign sinkVec_queue_34_deq_bits_data = _sinkVec_queue_fifo_34_empty ? sinkVec_queue_34_enq_bits_data : sinkVec_queue_dataOut_34_data;
  assign sinkVec_queue_34_deq_bits_last = ~_sinkVec_queue_fifo_34_empty & sinkVec_queue_dataOut_34_last;
  assign sinkVec_queue_34_deq_bits_instructionIndex = _sinkVec_queue_fifo_34_empty ? sinkVec_queue_34_enq_bits_instructionIndex : sinkVec_queue_dataOut_34_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_34;
  wire         sinkVec_releasePipe_pipe_out_34_valid = sinkVec_releasePipe_pipe_v_34;
  wire         x22_8_0_ready;
  wire         x22_8_0_valid;
  wire         sinkVec_validSource_34_valid = x22_8_0_ready & x22_8_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_34;
  wire [2:0]   sinkVec_tokenCheck_counterChange_34 = sinkVec_validSource_34_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_34 = ~(sinkVec_tokenCheck_counter_34[2]);
  assign x22_8_0_ready = sinkVec_tokenCheck_34;
  assign sinkVec_queue_34_enq_valid = sinkVec_validSink_34_valid;
  assign sinkVec_queue_34_enq_bits_vd = sinkVec_validSink_34_bits_vd;
  assign sinkVec_queue_34_enq_bits_offset = sinkVec_validSink_34_bits_offset;
  assign sinkVec_queue_34_enq_bits_mask = sinkVec_validSink_34_bits_mask;
  assign sinkVec_queue_34_enq_bits_data = sinkVec_validSink_34_bits_data;
  assign sinkVec_queue_34_enq_bits_instructionIndex = sinkVec_validSink_34_bits_instructionIndex;
  reg          sinkVec_shifterReg_34_0_valid;
  assign sinkVec_validSink_34_valid = sinkVec_shifterReg_34_0_valid;
  reg  [4:0]   sinkVec_shifterReg_34_0_bits_vd;
  assign sinkVec_validSink_34_bits_vd = sinkVec_shifterReg_34_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_34_0_bits_offset;
  assign sinkVec_validSink_34_bits_offset = sinkVec_shifterReg_34_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_34_0_bits_mask;
  assign sinkVec_validSink_34_bits_mask = sinkVec_shifterReg_34_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_34_0_bits_data;
  assign sinkVec_validSink_34_bits_data = sinkVec_shifterReg_34_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_34_0_bits_instructionIndex;
  assign sinkVec_validSink_34_bits_instructionIndex = sinkVec_shifterReg_34_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_34 = sinkVec_shifterReg_34_0_valid | sinkVec_validSource_34_valid;
  wire         sinkVec_17_1_ready;
  wire         sinkVec_queue_35_deq_ready = sinkVec_sinkWire_35_ready;
  wire         sinkVec_queue_35_deq_valid;
  wire [4:0]   sinkVec_queue_35_deq_bits_vd;
  wire         sinkVec_17_1_valid = sinkVec_sinkWire_35_valid;
  wire [1:0]   sinkVec_queue_35_deq_bits_offset;
  wire [4:0]   sinkVec_17_1_bits_vd = sinkVec_sinkWire_35_bits_vd;
  wire [3:0]   sinkVec_queue_35_deq_bits_mask;
  wire [1:0]   sinkVec_17_1_bits_offset = sinkVec_sinkWire_35_bits_offset;
  wire [31:0]  sinkVec_queue_35_deq_bits_data;
  wire [3:0]   sinkVec_17_1_bits_mask = sinkVec_sinkWire_35_bits_mask;
  wire         sinkVec_queue_35_deq_bits_last;
  wire [31:0]  sinkVec_17_1_bits_data = sinkVec_sinkWire_35_bits_data;
  wire [2:0]   sinkVec_queue_35_deq_bits_instructionIndex;
  wire         sinkVec_17_1_bits_last = sinkVec_sinkWire_35_bits_last;
  wire [2:0]   sinkVec_17_1_bits_instructionIndex = sinkVec_sinkWire_35_bits_instructionIndex;
  wire         sinkVec_validSink_35_valid;
  wire [4:0]   sinkVec_validSink_35_bits_vd;
  wire [1:0]   sinkVec_validSink_35_bits_offset;
  wire [3:0]   sinkVec_validSink_35_bits_mask;
  wire [31:0]  sinkVec_validSink_35_bits_data;
  wire         sinkVec_validSink_35_bits_last;
  wire [2:0]   sinkVec_validSink_35_bits_instructionIndex;
  assign sinkVec_sinkWire_35_valid = sinkVec_queue_35_deq_valid;
  assign sinkVec_sinkWire_35_bits_vd = sinkVec_queue_35_deq_bits_vd;
  assign sinkVec_sinkWire_35_bits_offset = sinkVec_queue_35_deq_bits_offset;
  assign sinkVec_sinkWire_35_bits_mask = sinkVec_queue_35_deq_bits_mask;
  assign sinkVec_sinkWire_35_bits_data = sinkVec_queue_35_deq_bits_data;
  assign sinkVec_sinkWire_35_bits_last = sinkVec_queue_35_deq_bits_last;
  assign sinkVec_sinkWire_35_bits_instructionIndex = sinkVec_queue_35_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_35_enq_bits_data;
  wire         sinkVec_queue_35_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_17 = {sinkVec_queue_35_enq_bits_data, sinkVec_queue_35_enq_bits_last};
  wire [2:0]   sinkVec_queue_35_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_35 = {sinkVec_queue_dataIn_lo_hi_17, sinkVec_queue_35_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_35_enq_bits_vd;
  wire [1:0]   sinkVec_queue_35_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_17 = {sinkVec_queue_35_enq_bits_vd, sinkVec_queue_35_enq_bits_offset};
  wire [3:0]   sinkVec_queue_35_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_35 = {sinkVec_queue_dataIn_hi_hi_17, sinkVec_queue_35_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_35 = {sinkVec_queue_dataIn_hi_35, sinkVec_queue_dataIn_lo_35};
  wire [2:0]   sinkVec_queue_dataOut_35_instructionIndex = _sinkVec_queue_fifo_35_data_out[2:0];
  wire         sinkVec_queue_dataOut_35_last = _sinkVec_queue_fifo_35_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_35_data = _sinkVec_queue_fifo_35_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_35_mask = _sinkVec_queue_fifo_35_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_35_offset = _sinkVec_queue_fifo_35_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_35_vd = _sinkVec_queue_fifo_35_data_out[46:42];
  wire         sinkVec_queue_35_enq_ready = ~_sinkVec_queue_fifo_35_full;
  wire         sinkVec_queue_35_enq_valid;
  assign sinkVec_queue_35_deq_valid = ~_sinkVec_queue_fifo_35_empty | sinkVec_queue_35_enq_valid;
  assign sinkVec_queue_35_deq_bits_vd = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_vd : sinkVec_queue_dataOut_35_vd;
  assign sinkVec_queue_35_deq_bits_offset = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_offset : sinkVec_queue_dataOut_35_offset;
  assign sinkVec_queue_35_deq_bits_mask = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_mask : sinkVec_queue_dataOut_35_mask;
  assign sinkVec_queue_35_deq_bits_data = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_data : sinkVec_queue_dataOut_35_data;
  assign sinkVec_queue_35_deq_bits_last = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_last : sinkVec_queue_dataOut_35_last;
  assign sinkVec_queue_35_deq_bits_instructionIndex = _sinkVec_queue_fifo_35_empty ? sinkVec_queue_35_enq_bits_instructionIndex : sinkVec_queue_dataOut_35_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_35;
  wire         sinkVec_releasePipe_pipe_out_35_valid = sinkVec_releasePipe_pipe_v_35;
  wire         x22_8_1_ready;
  wire         x22_8_1_valid;
  wire         sinkVec_validSource_35_valid = x22_8_1_ready & x22_8_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_35;
  wire [2:0]   sinkVec_tokenCheck_counterChange_35 = sinkVec_validSource_35_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_35 = ~(sinkVec_tokenCheck_counter_35[2]);
  assign x22_8_1_ready = sinkVec_tokenCheck_35;
  assign sinkVec_queue_35_enq_valid = sinkVec_validSink_35_valid;
  assign sinkVec_queue_35_enq_bits_vd = sinkVec_validSink_35_bits_vd;
  assign sinkVec_queue_35_enq_bits_offset = sinkVec_validSink_35_bits_offset;
  assign sinkVec_queue_35_enq_bits_mask = sinkVec_validSink_35_bits_mask;
  assign sinkVec_queue_35_enq_bits_data = sinkVec_validSink_35_bits_data;
  assign sinkVec_queue_35_enq_bits_last = sinkVec_validSink_35_bits_last;
  assign sinkVec_queue_35_enq_bits_instructionIndex = sinkVec_validSink_35_bits_instructionIndex;
  reg          sinkVec_shifterReg_35_0_valid;
  assign sinkVec_validSink_35_valid = sinkVec_shifterReg_35_0_valid;
  reg  [4:0]   sinkVec_shifterReg_35_0_bits_vd;
  assign sinkVec_validSink_35_bits_vd = sinkVec_shifterReg_35_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_35_0_bits_offset;
  assign sinkVec_validSink_35_bits_offset = sinkVec_shifterReg_35_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_35_0_bits_mask;
  assign sinkVec_validSink_35_bits_mask = sinkVec_shifterReg_35_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_35_0_bits_data;
  assign sinkVec_validSink_35_bits_data = sinkVec_shifterReg_35_0_bits_data;
  reg          sinkVec_shifterReg_35_0_bits_last;
  assign sinkVec_validSink_35_bits_last = sinkVec_shifterReg_35_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_35_0_bits_instructionIndex;
  assign sinkVec_validSink_35_bits_instructionIndex = sinkVec_shifterReg_35_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_35 = sinkVec_shifterReg_35_0_valid | sinkVec_validSource_35_valid;
  assign sinkVec_sinkWire_34_ready = sinkVec_17_0_ready;
  assign sinkVec_sinkWire_35_ready = sinkVec_17_1_ready;
  reg          maskUnitFirst_17;
  wire         tryToRead_17 = sinkVec_17_0_valid | sinkVec_17_1_valid;
  wire         sinkWire_17_valid = maskUnitFirst_17 ? sinkVec_17_0_valid : sinkVec_17_1_valid;
  wire [4:0]   sinkWire_17_bits_vd = maskUnitFirst_17 ? sinkVec_17_0_bits_vd : sinkVec_17_1_bits_vd;
  wire [1:0]   sinkWire_17_bits_offset = maskUnitFirst_17 ? sinkVec_17_0_bits_offset : sinkVec_17_1_bits_offset;
  wire [3:0]   sinkWire_17_bits_mask = maskUnitFirst_17 ? sinkVec_17_0_bits_mask : sinkVec_17_1_bits_mask;
  wire [31:0]  sinkWire_17_bits_data = maskUnitFirst_17 ? sinkVec_17_0_bits_data : sinkVec_17_1_bits_data;
  wire         sinkWire_17_bits_last = maskUnitFirst_17 ? sinkVec_17_0_bits_last : sinkVec_17_1_bits_last;
  wire [2:0]   sinkWire_17_bits_instructionIndex = maskUnitFirst_17 ? sinkVec_17_0_bits_instructionIndex : sinkVec_17_1_bits_instructionIndex;
  wire         sinkWire_17_ready;
  assign sinkVec_17_1_ready = sinkWire_17_ready & ~maskUnitFirst_17;
  assign sinkVec_17_0_ready = sinkWire_17_ready & maskUnitFirst_17;
  reg          view__writeRelease_8_pipe_v;
  wire         view__writeRelease_8_pipe_out_valid = view__writeRelease_8_pipe_v;
  reg          pipe_v_24;
  wire         pipe_out_16_valid = pipe_v_24;
  wire         _probeWire_writeQueueEnqVec_8_valid_T = x22_8_0_ready & _maskUnit_exeResp_8_valid;
  reg          instructionFinishedPipe_pipe_v_8;
  wire         instructionFinishedPipe_pipe_out_8_valid = instructionFinishedPipe_pipe_v_8;
  reg  [7:0]   instructionFinishedPipe_pipe_b_8;
  wire [7:0]   instructionFinishedPipe_pipe_out_8_bits = instructionFinishedPipe_pipe_b_8;
  wire         instructionFinished_8_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_8_bits);
  wire         instructionFinished_8_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_8_bits);
  wire         instructionFinished_8_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_8_bits);
  wire         instructionFinished_8_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_8_bits);
  assign vxsatReportVec_8 = _laneVec_8_vxsatReport[3:0];
  reg          pipe_v_25;
  reg  [31:0]  pipe_b_25;
  reg          pipe_pipe_v_8;
  wire         pipe_pipe_out_8_valid = pipe_pipe_v_8;
  reg  [31:0]  pipe_pipe_b_8;
  wire [31:0]  pipe_pipe_out_8_bits = pipe_pipe_b_8;
  reg          view__laneMaskSelect_8_pipe_v;
  reg  [5:0]   view__laneMaskSelect_8_pipe_b;
  reg          view__laneMaskSelect_8_pipe_pipe_v;
  wire         view__laneMaskSelect_8_pipe_pipe_out_valid = view__laneMaskSelect_8_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_8_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_8_pipe_pipe_out_bits = view__laneMaskSelect_8_pipe_pipe_b;
  reg          view__laneMaskSewSelect_8_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_8_pipe_b;
  reg          view__laneMaskSewSelect_8_pipe_pipe_v;
  wire         view__laneMaskSewSelect_8_pipe_pipe_out_valid = view__laneMaskSewSelect_8_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_8_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_8_pipe_pipe_out_bits = view__laneMaskSewSelect_8_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_8;
  wire         lsuLastPipe_pipe_out_8_valid = lsuLastPipe_pipe_v_8;
  reg  [7:0]   lsuLastPipe_pipe_b_8;
  wire [7:0]   lsuLastPipe_pipe_out_8_bits = lsuLastPipe_pipe_b_8;
  reg          maskLastPipe_pipe_v_8;
  wire         maskLastPipe_pipe_out_8_valid = maskLastPipe_pipe_v_8;
  reg  [7:0]   maskLastPipe_pipe_b_8;
  wire [7:0]   maskLastPipe_pipe_out_8_bits = maskLastPipe_pipe_b_8;
  wire [5:0]   writeCounter_8 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h20};
  reg          pipe_v_26;
  wire         pipe_out_17_valid = pipe_v_26;
  reg  [5:0]   pipe_b_26;
  wire [5:0]   pipe_out_17_bits = pipe_b_26;
  assign laneRequestSinkWire_9_ready = ~laneRequestSinkWire_9_bits_issueInst | _laneVec_9_laneRequest_ready;
  wire         sinkVec_tokenCheck_36;
  wire [4:0]   sinkVec_validSource_36_bits_vs = x13_9_0_bits_vs;
  wire [1:0]   sinkVec_validSource_36_bits_offset = x13_9_0_bits_offset;
  wire [2:0]   sinkVec_validSource_36_bits_instructionIndex = x13_9_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_37;
  wire [4:0]   sinkVec_validSource_37_bits_vs = x13_9_1_bits_vs;
  wire [1:0]   sinkVec_validSource_37_bits_offset = x13_9_1_bits_offset;
  wire [2:0]   sinkVec_validSource_37_bits_instructionIndex = x13_9_1_bits_instructionIndex;
  wire         sinkVec_18_0_ready;
  wire         sinkVec_queue_36_deq_ready = sinkVec_sinkWire_36_ready;
  wire         sinkVec_queue_36_deq_valid;
  wire [4:0]   sinkVec_queue_36_deq_bits_vs;
  wire         sinkVec_18_0_valid = sinkVec_sinkWire_36_valid;
  wire [1:0]   sinkVec_queue_36_deq_bits_readSource;
  wire [4:0]   sinkVec_18_0_bits_vs = sinkVec_sinkWire_36_bits_vs;
  wire [1:0]   sinkVec_queue_36_deq_bits_offset;
  wire [1:0]   sinkVec_18_0_bits_readSource = sinkVec_sinkWire_36_bits_readSource;
  wire [2:0]   sinkVec_queue_36_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_18_0_bits_offset = sinkVec_sinkWire_36_bits_offset;
  wire [2:0]   sinkVec_18_0_bits_instructionIndex = sinkVec_sinkWire_36_bits_instructionIndex;
  wire         sinkVec_validSink_36_valid;
  wire [4:0]   sinkVec_validSink_36_bits_vs;
  wire [1:0]   sinkVec_validSink_36_bits_readSource;
  wire [1:0]   sinkVec_validSink_36_bits_offset;
  wire [2:0]   sinkVec_validSink_36_bits_instructionIndex;
  assign sinkVec_sinkWire_36_valid = sinkVec_queue_36_deq_valid;
  assign sinkVec_sinkWire_36_bits_vs = sinkVec_queue_36_deq_bits_vs;
  assign sinkVec_sinkWire_36_bits_readSource = sinkVec_queue_36_deq_bits_readSource;
  assign sinkVec_sinkWire_36_bits_offset = sinkVec_queue_36_deq_bits_offset;
  assign sinkVec_sinkWire_36_bits_instructionIndex = sinkVec_queue_36_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_36_enq_bits_offset;
  wire [2:0]   sinkVec_queue_36_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_36 = {sinkVec_queue_36_enq_bits_offset, sinkVec_queue_36_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_36_enq_bits_vs;
  wire [1:0]   sinkVec_queue_36_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_36 = {sinkVec_queue_36_enq_bits_vs, sinkVec_queue_36_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_36 = {sinkVec_queue_dataIn_hi_36, sinkVec_queue_dataIn_lo_36};
  wire [2:0]   sinkVec_queue_dataOut_36_instructionIndex = _sinkVec_queue_fifo_36_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_36_offset = _sinkVec_queue_fifo_36_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_36_readSource = _sinkVec_queue_fifo_36_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_36_vs = _sinkVec_queue_fifo_36_data_out[11:7];
  wire         sinkVec_queue_36_enq_ready = ~_sinkVec_queue_fifo_36_full;
  wire         sinkVec_queue_36_enq_valid;
  assign sinkVec_queue_36_deq_valid = ~_sinkVec_queue_fifo_36_empty | sinkVec_queue_36_enq_valid;
  assign sinkVec_queue_36_deq_bits_vs = _sinkVec_queue_fifo_36_empty ? sinkVec_queue_36_enq_bits_vs : sinkVec_queue_dataOut_36_vs;
  assign sinkVec_queue_36_deq_bits_readSource = _sinkVec_queue_fifo_36_empty ? sinkVec_queue_36_enq_bits_readSource : sinkVec_queue_dataOut_36_readSource;
  assign sinkVec_queue_36_deq_bits_offset = _sinkVec_queue_fifo_36_empty ? sinkVec_queue_36_enq_bits_offset : sinkVec_queue_dataOut_36_offset;
  assign sinkVec_queue_36_deq_bits_instructionIndex = _sinkVec_queue_fifo_36_empty ? sinkVec_queue_36_enq_bits_instructionIndex : sinkVec_queue_dataOut_36_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_36;
  wire         sinkVec_releasePipe_pipe_out_36_valid = sinkVec_releasePipe_pipe_v_36;
  wire         x13_9_0_ready;
  wire         x13_9_0_valid;
  wire         sinkVec_validSource_36_valid = x13_9_0_ready & x13_9_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_36;
  wire [2:0]   sinkVec_tokenCheck_counterChange_36 = sinkVec_validSource_36_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_36 = ~(sinkVec_tokenCheck_counter_36[2]);
  assign x13_9_0_ready = sinkVec_tokenCheck_36;
  assign sinkVec_queue_36_enq_valid = sinkVec_validSink_36_valid;
  assign sinkVec_queue_36_enq_bits_vs = sinkVec_validSink_36_bits_vs;
  assign sinkVec_queue_36_enq_bits_readSource = sinkVec_validSink_36_bits_readSource;
  assign sinkVec_queue_36_enq_bits_offset = sinkVec_validSink_36_bits_offset;
  assign sinkVec_queue_36_enq_bits_instructionIndex = sinkVec_validSink_36_bits_instructionIndex;
  reg          sinkVec_shifterReg_36_0_valid;
  assign sinkVec_validSink_36_valid = sinkVec_shifterReg_36_0_valid;
  reg  [4:0]   sinkVec_shifterReg_36_0_bits_vs;
  assign sinkVec_validSink_36_bits_vs = sinkVec_shifterReg_36_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_36_0_bits_readSource;
  assign sinkVec_validSink_36_bits_readSource = sinkVec_shifterReg_36_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_36_0_bits_offset;
  assign sinkVec_validSink_36_bits_offset = sinkVec_shifterReg_36_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_36_0_bits_instructionIndex;
  assign sinkVec_validSink_36_bits_instructionIndex = sinkVec_shifterReg_36_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_36 = sinkVec_shifterReg_36_0_valid | sinkVec_validSource_36_valid;
  wire         sinkVec_18_1_ready;
  wire         sinkVec_queue_37_deq_ready = sinkVec_sinkWire_37_ready;
  wire         sinkVec_queue_37_deq_valid;
  wire [4:0]   sinkVec_queue_37_deq_bits_vs;
  wire         sinkVec_18_1_valid = sinkVec_sinkWire_37_valid;
  wire [1:0]   sinkVec_queue_37_deq_bits_readSource;
  wire [4:0]   sinkVec_18_1_bits_vs = sinkVec_sinkWire_37_bits_vs;
  wire [1:0]   sinkVec_queue_37_deq_bits_offset;
  wire [1:0]   sinkVec_18_1_bits_readSource = sinkVec_sinkWire_37_bits_readSource;
  wire [2:0]   sinkVec_queue_37_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_18_1_bits_offset = sinkVec_sinkWire_37_bits_offset;
  wire [2:0]   sinkVec_18_1_bits_instructionIndex = sinkVec_sinkWire_37_bits_instructionIndex;
  wire         sinkVec_validSink_37_valid;
  wire [4:0]   sinkVec_validSink_37_bits_vs;
  wire [1:0]   sinkVec_validSink_37_bits_readSource;
  wire [1:0]   sinkVec_validSink_37_bits_offset;
  wire [2:0]   sinkVec_validSink_37_bits_instructionIndex;
  assign sinkVec_sinkWire_37_valid = sinkVec_queue_37_deq_valid;
  assign sinkVec_sinkWire_37_bits_vs = sinkVec_queue_37_deq_bits_vs;
  assign sinkVec_sinkWire_37_bits_readSource = sinkVec_queue_37_deq_bits_readSource;
  assign sinkVec_sinkWire_37_bits_offset = sinkVec_queue_37_deq_bits_offset;
  assign sinkVec_sinkWire_37_bits_instructionIndex = sinkVec_queue_37_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_37_enq_bits_offset;
  wire [2:0]   sinkVec_queue_37_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_37 = {sinkVec_queue_37_enq_bits_offset, sinkVec_queue_37_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_37_enq_bits_vs;
  wire [1:0]   sinkVec_queue_37_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_37 = {sinkVec_queue_37_enq_bits_vs, sinkVec_queue_37_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_37 = {sinkVec_queue_dataIn_hi_37, sinkVec_queue_dataIn_lo_37};
  wire [2:0]   sinkVec_queue_dataOut_37_instructionIndex = _sinkVec_queue_fifo_37_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_37_offset = _sinkVec_queue_fifo_37_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_37_readSource = _sinkVec_queue_fifo_37_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_37_vs = _sinkVec_queue_fifo_37_data_out[11:7];
  wire         sinkVec_queue_37_enq_ready = ~_sinkVec_queue_fifo_37_full;
  wire         sinkVec_queue_37_enq_valid;
  assign sinkVec_queue_37_deq_valid = ~_sinkVec_queue_fifo_37_empty | sinkVec_queue_37_enq_valid;
  assign sinkVec_queue_37_deq_bits_vs = _sinkVec_queue_fifo_37_empty ? sinkVec_queue_37_enq_bits_vs : sinkVec_queue_dataOut_37_vs;
  assign sinkVec_queue_37_deq_bits_readSource = _sinkVec_queue_fifo_37_empty ? sinkVec_queue_37_enq_bits_readSource : sinkVec_queue_dataOut_37_readSource;
  assign sinkVec_queue_37_deq_bits_offset = _sinkVec_queue_fifo_37_empty ? sinkVec_queue_37_enq_bits_offset : sinkVec_queue_dataOut_37_offset;
  assign sinkVec_queue_37_deq_bits_instructionIndex = _sinkVec_queue_fifo_37_empty ? sinkVec_queue_37_enq_bits_instructionIndex : sinkVec_queue_dataOut_37_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_37;
  wire         sinkVec_releasePipe_pipe_out_37_valid = sinkVec_releasePipe_pipe_v_37;
  wire         x13_9_1_ready;
  wire         x13_9_1_valid;
  wire         sinkVec_validSource_37_valid = x13_9_1_ready & x13_9_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_37;
  wire [2:0]   sinkVec_tokenCheck_counterChange_37 = sinkVec_validSource_37_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_37 = ~(sinkVec_tokenCheck_counter_37[2]);
  assign x13_9_1_ready = sinkVec_tokenCheck_37;
  assign sinkVec_queue_37_enq_valid = sinkVec_validSink_37_valid;
  assign sinkVec_queue_37_enq_bits_vs = sinkVec_validSink_37_bits_vs;
  assign sinkVec_queue_37_enq_bits_readSource = sinkVec_validSink_37_bits_readSource;
  assign sinkVec_queue_37_enq_bits_offset = sinkVec_validSink_37_bits_offset;
  assign sinkVec_queue_37_enq_bits_instructionIndex = sinkVec_validSink_37_bits_instructionIndex;
  reg          sinkVec_shifterReg_37_0_valid;
  assign sinkVec_validSink_37_valid = sinkVec_shifterReg_37_0_valid;
  reg  [4:0]   sinkVec_shifterReg_37_0_bits_vs;
  assign sinkVec_validSink_37_bits_vs = sinkVec_shifterReg_37_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_37_0_bits_readSource;
  assign sinkVec_validSink_37_bits_readSource = sinkVec_shifterReg_37_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_37_0_bits_offset;
  assign sinkVec_validSink_37_bits_offset = sinkVec_shifterReg_37_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_37_0_bits_instructionIndex;
  assign sinkVec_validSink_37_bits_instructionIndex = sinkVec_shifterReg_37_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_37 = sinkVec_shifterReg_37_0_valid | sinkVec_validSource_37_valid;
  assign sinkVec_sinkWire_36_ready = sinkVec_18_0_ready;
  assign sinkVec_sinkWire_37_ready = sinkVec_18_1_ready;
  reg          maskUnitFirst_18;
  wire         tryToRead_18 = sinkVec_18_0_valid | sinkVec_18_1_valid;
  wire         sinkWire_18_valid = maskUnitFirst_18 ? sinkVec_18_0_valid : sinkVec_18_1_valid;
  wire [4:0]   sinkWire_18_bits_vs = maskUnitFirst_18 ? sinkVec_18_0_bits_vs : sinkVec_18_1_bits_vs;
  wire [1:0]   sinkWire_18_bits_readSource = maskUnitFirst_18 ? sinkVec_18_0_bits_readSource : sinkVec_18_1_bits_readSource;
  wire [1:0]   sinkWire_18_bits_offset = maskUnitFirst_18 ? sinkVec_18_0_bits_offset : sinkVec_18_1_bits_offset;
  wire [2:0]   sinkWire_18_bits_instructionIndex = maskUnitFirst_18 ? sinkVec_18_0_bits_instructionIndex : sinkVec_18_1_bits_instructionIndex;
  wire         sinkWire_18_ready;
  assign sinkVec_18_1_ready = sinkWire_18_ready & ~maskUnitFirst_18;
  assign sinkVec_18_0_ready = sinkWire_18_ready & maskUnitFirst_18;
  reg          accessDataValid_pipe_v_18;
  reg          accessDataValid_pipe_pipe_v_18;
  wire         accessDataValid_pipe_pipe_out_18_valid = accessDataValid_pipe_pipe_v_18;
  wire         accessDataSource_18_valid = accessDataValid_pipe_pipe_out_18_valid;
  reg          shifterReg_34_0_valid;
  reg  [31:0]  shifterReg_34_0_bits;
  wire         shifterValid_34 = shifterReg_34_0_valid | accessDataSource_18_valid;
  reg          accessDataValid_pipe_v_19;
  reg          accessDataValid_pipe_pipe_v_19;
  wire         accessDataValid_pipe_pipe_out_19_valid = accessDataValid_pipe_pipe_v_19;
  wire         accessDataSource_19_valid = accessDataValid_pipe_pipe_out_19_valid;
  reg          shifterReg_35_0_valid;
  reg  [31:0]  shifterReg_35_0_bits;
  wire         shifterValid_35 = shifterReg_35_0_valid | accessDataSource_19_valid;
  wire         sinkVec_tokenCheck_38;
  wire [4:0]   sinkVec_validSource_38_bits_vd = x22_9_0_bits_vd;
  wire [1:0]   sinkVec_validSource_38_bits_offset = x22_9_0_bits_offset;
  wire [3:0]   sinkVec_validSource_38_bits_mask = x22_9_0_bits_mask;
  wire [31:0]  sinkVec_validSource_38_bits_data = x22_9_0_bits_data;
  wire [2:0]   sinkVec_validSource_38_bits_instructionIndex = x22_9_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_39;
  wire [4:0]   sinkVec_validSource_39_bits_vd = x22_9_1_bits_vd;
  wire [1:0]   sinkVec_validSource_39_bits_offset = x22_9_1_bits_offset;
  wire [3:0]   sinkVec_validSource_39_bits_mask = x22_9_1_bits_mask;
  wire [31:0]  sinkVec_validSource_39_bits_data = x22_9_1_bits_data;
  wire         sinkVec_validSource_39_bits_last = x22_9_1_bits_last;
  wire [2:0]   sinkVec_validSource_39_bits_instructionIndex = x22_9_1_bits_instructionIndex;
  wire         sinkVec_19_0_ready;
  wire         sinkVec_queue_38_deq_ready = sinkVec_sinkWire_38_ready;
  wire         sinkVec_queue_38_deq_valid;
  wire [4:0]   sinkVec_queue_38_deq_bits_vd;
  wire         sinkVec_19_0_valid = sinkVec_sinkWire_38_valid;
  wire [1:0]   sinkVec_queue_38_deq_bits_offset;
  wire [4:0]   sinkVec_19_0_bits_vd = sinkVec_sinkWire_38_bits_vd;
  wire [3:0]   sinkVec_queue_38_deq_bits_mask;
  wire [1:0]   sinkVec_19_0_bits_offset = sinkVec_sinkWire_38_bits_offset;
  wire [31:0]  sinkVec_queue_38_deq_bits_data;
  wire [3:0]   sinkVec_19_0_bits_mask = sinkVec_sinkWire_38_bits_mask;
  wire         sinkVec_queue_38_deq_bits_last;
  wire [31:0]  sinkVec_19_0_bits_data = sinkVec_sinkWire_38_bits_data;
  wire [2:0]   sinkVec_queue_38_deq_bits_instructionIndex;
  wire         sinkVec_19_0_bits_last = sinkVec_sinkWire_38_bits_last;
  wire [2:0]   sinkVec_19_0_bits_instructionIndex = sinkVec_sinkWire_38_bits_instructionIndex;
  wire         sinkVec_validSink_38_valid;
  wire [4:0]   sinkVec_validSink_38_bits_vd;
  wire [1:0]   sinkVec_validSink_38_bits_offset;
  wire [3:0]   sinkVec_validSink_38_bits_mask;
  wire [31:0]  sinkVec_validSink_38_bits_data;
  wire [2:0]   sinkVec_validSink_38_bits_instructionIndex;
  assign sinkVec_sinkWire_38_valid = sinkVec_queue_38_deq_valid;
  assign sinkVec_sinkWire_38_bits_vd = sinkVec_queue_38_deq_bits_vd;
  assign sinkVec_sinkWire_38_bits_offset = sinkVec_queue_38_deq_bits_offset;
  assign sinkVec_sinkWire_38_bits_mask = sinkVec_queue_38_deq_bits_mask;
  assign sinkVec_sinkWire_38_bits_data = sinkVec_queue_38_deq_bits_data;
  assign sinkVec_sinkWire_38_bits_last = sinkVec_queue_38_deq_bits_last;
  assign sinkVec_sinkWire_38_bits_instructionIndex = sinkVec_queue_38_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_38_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_18 = {sinkVec_queue_38_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_38_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_38 = {sinkVec_queue_dataIn_lo_hi_18, sinkVec_queue_38_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_38_enq_bits_vd;
  wire [1:0]   sinkVec_queue_38_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_18 = {sinkVec_queue_38_enq_bits_vd, sinkVec_queue_38_enq_bits_offset};
  wire [3:0]   sinkVec_queue_38_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_38 = {sinkVec_queue_dataIn_hi_hi_18, sinkVec_queue_38_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_38 = {sinkVec_queue_dataIn_hi_38, sinkVec_queue_dataIn_lo_38};
  wire [2:0]   sinkVec_queue_dataOut_38_instructionIndex = _sinkVec_queue_fifo_38_data_out[2:0];
  wire         sinkVec_queue_dataOut_38_last = _sinkVec_queue_fifo_38_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_38_data = _sinkVec_queue_fifo_38_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_38_mask = _sinkVec_queue_fifo_38_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_38_offset = _sinkVec_queue_fifo_38_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_38_vd = _sinkVec_queue_fifo_38_data_out[46:42];
  wire         sinkVec_queue_38_enq_ready = ~_sinkVec_queue_fifo_38_full;
  wire         sinkVec_queue_38_enq_valid;
  assign sinkVec_queue_38_deq_valid = ~_sinkVec_queue_fifo_38_empty | sinkVec_queue_38_enq_valid;
  assign sinkVec_queue_38_deq_bits_vd = _sinkVec_queue_fifo_38_empty ? sinkVec_queue_38_enq_bits_vd : sinkVec_queue_dataOut_38_vd;
  assign sinkVec_queue_38_deq_bits_offset = _sinkVec_queue_fifo_38_empty ? sinkVec_queue_38_enq_bits_offset : sinkVec_queue_dataOut_38_offset;
  assign sinkVec_queue_38_deq_bits_mask = _sinkVec_queue_fifo_38_empty ? sinkVec_queue_38_enq_bits_mask : sinkVec_queue_dataOut_38_mask;
  assign sinkVec_queue_38_deq_bits_data = _sinkVec_queue_fifo_38_empty ? sinkVec_queue_38_enq_bits_data : sinkVec_queue_dataOut_38_data;
  assign sinkVec_queue_38_deq_bits_last = ~_sinkVec_queue_fifo_38_empty & sinkVec_queue_dataOut_38_last;
  assign sinkVec_queue_38_deq_bits_instructionIndex = _sinkVec_queue_fifo_38_empty ? sinkVec_queue_38_enq_bits_instructionIndex : sinkVec_queue_dataOut_38_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_38;
  wire         sinkVec_releasePipe_pipe_out_38_valid = sinkVec_releasePipe_pipe_v_38;
  wire         x22_9_0_ready;
  wire         x22_9_0_valid;
  wire         sinkVec_validSource_38_valid = x22_9_0_ready & x22_9_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_38;
  wire [2:0]   sinkVec_tokenCheck_counterChange_38 = sinkVec_validSource_38_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_38 = ~(sinkVec_tokenCheck_counter_38[2]);
  assign x22_9_0_ready = sinkVec_tokenCheck_38;
  assign sinkVec_queue_38_enq_valid = sinkVec_validSink_38_valid;
  assign sinkVec_queue_38_enq_bits_vd = sinkVec_validSink_38_bits_vd;
  assign sinkVec_queue_38_enq_bits_offset = sinkVec_validSink_38_bits_offset;
  assign sinkVec_queue_38_enq_bits_mask = sinkVec_validSink_38_bits_mask;
  assign sinkVec_queue_38_enq_bits_data = sinkVec_validSink_38_bits_data;
  assign sinkVec_queue_38_enq_bits_instructionIndex = sinkVec_validSink_38_bits_instructionIndex;
  reg          sinkVec_shifterReg_38_0_valid;
  assign sinkVec_validSink_38_valid = sinkVec_shifterReg_38_0_valid;
  reg  [4:0]   sinkVec_shifterReg_38_0_bits_vd;
  assign sinkVec_validSink_38_bits_vd = sinkVec_shifterReg_38_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_38_0_bits_offset;
  assign sinkVec_validSink_38_bits_offset = sinkVec_shifterReg_38_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_38_0_bits_mask;
  assign sinkVec_validSink_38_bits_mask = sinkVec_shifterReg_38_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_38_0_bits_data;
  assign sinkVec_validSink_38_bits_data = sinkVec_shifterReg_38_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_38_0_bits_instructionIndex;
  assign sinkVec_validSink_38_bits_instructionIndex = sinkVec_shifterReg_38_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_38 = sinkVec_shifterReg_38_0_valid | sinkVec_validSource_38_valid;
  wire         sinkVec_19_1_ready;
  wire         sinkVec_queue_39_deq_ready = sinkVec_sinkWire_39_ready;
  wire         sinkVec_queue_39_deq_valid;
  wire [4:0]   sinkVec_queue_39_deq_bits_vd;
  wire         sinkVec_19_1_valid = sinkVec_sinkWire_39_valid;
  wire [1:0]   sinkVec_queue_39_deq_bits_offset;
  wire [4:0]   sinkVec_19_1_bits_vd = sinkVec_sinkWire_39_bits_vd;
  wire [3:0]   sinkVec_queue_39_deq_bits_mask;
  wire [1:0]   sinkVec_19_1_bits_offset = sinkVec_sinkWire_39_bits_offset;
  wire [31:0]  sinkVec_queue_39_deq_bits_data;
  wire [3:0]   sinkVec_19_1_bits_mask = sinkVec_sinkWire_39_bits_mask;
  wire         sinkVec_queue_39_deq_bits_last;
  wire [31:0]  sinkVec_19_1_bits_data = sinkVec_sinkWire_39_bits_data;
  wire [2:0]   sinkVec_queue_39_deq_bits_instructionIndex;
  wire         sinkVec_19_1_bits_last = sinkVec_sinkWire_39_bits_last;
  wire [2:0]   sinkVec_19_1_bits_instructionIndex = sinkVec_sinkWire_39_bits_instructionIndex;
  wire         sinkVec_validSink_39_valid;
  wire [4:0]   sinkVec_validSink_39_bits_vd;
  wire [1:0]   sinkVec_validSink_39_bits_offset;
  wire [3:0]   sinkVec_validSink_39_bits_mask;
  wire [31:0]  sinkVec_validSink_39_bits_data;
  wire         sinkVec_validSink_39_bits_last;
  wire [2:0]   sinkVec_validSink_39_bits_instructionIndex;
  assign sinkVec_sinkWire_39_valid = sinkVec_queue_39_deq_valid;
  assign sinkVec_sinkWire_39_bits_vd = sinkVec_queue_39_deq_bits_vd;
  assign sinkVec_sinkWire_39_bits_offset = sinkVec_queue_39_deq_bits_offset;
  assign sinkVec_sinkWire_39_bits_mask = sinkVec_queue_39_deq_bits_mask;
  assign sinkVec_sinkWire_39_bits_data = sinkVec_queue_39_deq_bits_data;
  assign sinkVec_sinkWire_39_bits_last = sinkVec_queue_39_deq_bits_last;
  assign sinkVec_sinkWire_39_bits_instructionIndex = sinkVec_queue_39_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_39_enq_bits_data;
  wire         sinkVec_queue_39_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_19 = {sinkVec_queue_39_enq_bits_data, sinkVec_queue_39_enq_bits_last};
  wire [2:0]   sinkVec_queue_39_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_39 = {sinkVec_queue_dataIn_lo_hi_19, sinkVec_queue_39_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_39_enq_bits_vd;
  wire [1:0]   sinkVec_queue_39_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_19 = {sinkVec_queue_39_enq_bits_vd, sinkVec_queue_39_enq_bits_offset};
  wire [3:0]   sinkVec_queue_39_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_39 = {sinkVec_queue_dataIn_hi_hi_19, sinkVec_queue_39_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_39 = {sinkVec_queue_dataIn_hi_39, sinkVec_queue_dataIn_lo_39};
  wire [2:0]   sinkVec_queue_dataOut_39_instructionIndex = _sinkVec_queue_fifo_39_data_out[2:0];
  wire         sinkVec_queue_dataOut_39_last = _sinkVec_queue_fifo_39_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_39_data = _sinkVec_queue_fifo_39_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_39_mask = _sinkVec_queue_fifo_39_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_39_offset = _sinkVec_queue_fifo_39_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_39_vd = _sinkVec_queue_fifo_39_data_out[46:42];
  wire         sinkVec_queue_39_enq_ready = ~_sinkVec_queue_fifo_39_full;
  wire         sinkVec_queue_39_enq_valid;
  assign sinkVec_queue_39_deq_valid = ~_sinkVec_queue_fifo_39_empty | sinkVec_queue_39_enq_valid;
  assign sinkVec_queue_39_deq_bits_vd = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_vd : sinkVec_queue_dataOut_39_vd;
  assign sinkVec_queue_39_deq_bits_offset = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_offset : sinkVec_queue_dataOut_39_offset;
  assign sinkVec_queue_39_deq_bits_mask = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_mask : sinkVec_queue_dataOut_39_mask;
  assign sinkVec_queue_39_deq_bits_data = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_data : sinkVec_queue_dataOut_39_data;
  assign sinkVec_queue_39_deq_bits_last = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_last : sinkVec_queue_dataOut_39_last;
  assign sinkVec_queue_39_deq_bits_instructionIndex = _sinkVec_queue_fifo_39_empty ? sinkVec_queue_39_enq_bits_instructionIndex : sinkVec_queue_dataOut_39_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_39;
  wire         sinkVec_releasePipe_pipe_out_39_valid = sinkVec_releasePipe_pipe_v_39;
  wire         x22_9_1_ready;
  wire         x22_9_1_valid;
  wire         sinkVec_validSource_39_valid = x22_9_1_ready & x22_9_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_39;
  wire [2:0]   sinkVec_tokenCheck_counterChange_39 = sinkVec_validSource_39_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_39 = ~(sinkVec_tokenCheck_counter_39[2]);
  assign x22_9_1_ready = sinkVec_tokenCheck_39;
  assign sinkVec_queue_39_enq_valid = sinkVec_validSink_39_valid;
  assign sinkVec_queue_39_enq_bits_vd = sinkVec_validSink_39_bits_vd;
  assign sinkVec_queue_39_enq_bits_offset = sinkVec_validSink_39_bits_offset;
  assign sinkVec_queue_39_enq_bits_mask = sinkVec_validSink_39_bits_mask;
  assign sinkVec_queue_39_enq_bits_data = sinkVec_validSink_39_bits_data;
  assign sinkVec_queue_39_enq_bits_last = sinkVec_validSink_39_bits_last;
  assign sinkVec_queue_39_enq_bits_instructionIndex = sinkVec_validSink_39_bits_instructionIndex;
  reg          sinkVec_shifterReg_39_0_valid;
  assign sinkVec_validSink_39_valid = sinkVec_shifterReg_39_0_valid;
  reg  [4:0]   sinkVec_shifterReg_39_0_bits_vd;
  assign sinkVec_validSink_39_bits_vd = sinkVec_shifterReg_39_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_39_0_bits_offset;
  assign sinkVec_validSink_39_bits_offset = sinkVec_shifterReg_39_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_39_0_bits_mask;
  assign sinkVec_validSink_39_bits_mask = sinkVec_shifterReg_39_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_39_0_bits_data;
  assign sinkVec_validSink_39_bits_data = sinkVec_shifterReg_39_0_bits_data;
  reg          sinkVec_shifterReg_39_0_bits_last;
  assign sinkVec_validSink_39_bits_last = sinkVec_shifterReg_39_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_39_0_bits_instructionIndex;
  assign sinkVec_validSink_39_bits_instructionIndex = sinkVec_shifterReg_39_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_39 = sinkVec_shifterReg_39_0_valid | sinkVec_validSource_39_valid;
  assign sinkVec_sinkWire_38_ready = sinkVec_19_0_ready;
  assign sinkVec_sinkWire_39_ready = sinkVec_19_1_ready;
  reg          maskUnitFirst_19;
  wire         tryToRead_19 = sinkVec_19_0_valid | sinkVec_19_1_valid;
  wire         sinkWire_19_valid = maskUnitFirst_19 ? sinkVec_19_0_valid : sinkVec_19_1_valid;
  wire [4:0]   sinkWire_19_bits_vd = maskUnitFirst_19 ? sinkVec_19_0_bits_vd : sinkVec_19_1_bits_vd;
  wire [1:0]   sinkWire_19_bits_offset = maskUnitFirst_19 ? sinkVec_19_0_bits_offset : sinkVec_19_1_bits_offset;
  wire [3:0]   sinkWire_19_bits_mask = maskUnitFirst_19 ? sinkVec_19_0_bits_mask : sinkVec_19_1_bits_mask;
  wire [31:0]  sinkWire_19_bits_data = maskUnitFirst_19 ? sinkVec_19_0_bits_data : sinkVec_19_1_bits_data;
  wire         sinkWire_19_bits_last = maskUnitFirst_19 ? sinkVec_19_0_bits_last : sinkVec_19_1_bits_last;
  wire [2:0]   sinkWire_19_bits_instructionIndex = maskUnitFirst_19 ? sinkVec_19_0_bits_instructionIndex : sinkVec_19_1_bits_instructionIndex;
  wire         sinkWire_19_ready;
  assign sinkVec_19_1_ready = sinkWire_19_ready & ~maskUnitFirst_19;
  assign sinkVec_19_0_ready = sinkWire_19_ready & maskUnitFirst_19;
  reg          view__writeRelease_9_pipe_v;
  wire         view__writeRelease_9_pipe_out_valid = view__writeRelease_9_pipe_v;
  reg          pipe_v_27;
  wire         pipe_out_18_valid = pipe_v_27;
  wire         _probeWire_writeQueueEnqVec_9_valid_T = x22_9_0_ready & _maskUnit_exeResp_9_valid;
  reg          instructionFinishedPipe_pipe_v_9;
  wire         instructionFinishedPipe_pipe_out_9_valid = instructionFinishedPipe_pipe_v_9;
  reg  [7:0]   instructionFinishedPipe_pipe_b_9;
  wire [7:0]   instructionFinishedPipe_pipe_out_9_bits = instructionFinishedPipe_pipe_b_9;
  wire         instructionFinished_9_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_9_bits);
  wire         instructionFinished_9_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_9_bits);
  wire         instructionFinished_9_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_9_bits);
  wire         instructionFinished_9_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_9_bits);
  assign vxsatReportVec_9 = _laneVec_9_vxsatReport[3:0];
  reg          pipe_v_28;
  reg  [31:0]  pipe_b_28;
  reg          pipe_pipe_v_9;
  wire         pipe_pipe_out_9_valid = pipe_pipe_v_9;
  reg  [31:0]  pipe_pipe_b_9;
  wire [31:0]  pipe_pipe_out_9_bits = pipe_pipe_b_9;
  reg          view__laneMaskSelect_9_pipe_v;
  reg  [5:0]   view__laneMaskSelect_9_pipe_b;
  reg          view__laneMaskSelect_9_pipe_pipe_v;
  wire         view__laneMaskSelect_9_pipe_pipe_out_valid = view__laneMaskSelect_9_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_9_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_9_pipe_pipe_out_bits = view__laneMaskSelect_9_pipe_pipe_b;
  reg          view__laneMaskSewSelect_9_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_9_pipe_b;
  reg          view__laneMaskSewSelect_9_pipe_pipe_v;
  wire         view__laneMaskSewSelect_9_pipe_pipe_out_valid = view__laneMaskSewSelect_9_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_9_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_9_pipe_pipe_out_bits = view__laneMaskSewSelect_9_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_9;
  wire         lsuLastPipe_pipe_out_9_valid = lsuLastPipe_pipe_v_9;
  reg  [7:0]   lsuLastPipe_pipe_b_9;
  wire [7:0]   lsuLastPipe_pipe_out_9_bits = lsuLastPipe_pipe_b_9;
  reg          maskLastPipe_pipe_v_9;
  wire         maskLastPipe_pipe_out_9_valid = maskLastPipe_pipe_v_9;
  reg  [7:0]   maskLastPipe_pipe_b_9;
  wire [7:0]   maskLastPipe_pipe_out_9_bits = maskLastPipe_pipe_b_9;
  wire [5:0]   writeCounter_9 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h24};
  reg          pipe_v_29;
  wire         pipe_out_19_valid = pipe_v_29;
  reg  [5:0]   pipe_b_29;
  wire [5:0]   pipe_out_19_bits = pipe_b_29;
  assign laneRequestSinkWire_10_ready = ~laneRequestSinkWire_10_bits_issueInst | _laneVec_10_laneRequest_ready;
  wire         sinkVec_tokenCheck_40;
  wire [4:0]   sinkVec_validSource_40_bits_vs = x13_10_0_bits_vs;
  wire [1:0]   sinkVec_validSource_40_bits_offset = x13_10_0_bits_offset;
  wire [2:0]   sinkVec_validSource_40_bits_instructionIndex = x13_10_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_41;
  wire [4:0]   sinkVec_validSource_41_bits_vs = x13_10_1_bits_vs;
  wire [1:0]   sinkVec_validSource_41_bits_offset = x13_10_1_bits_offset;
  wire [2:0]   sinkVec_validSource_41_bits_instructionIndex = x13_10_1_bits_instructionIndex;
  wire         sinkVec_20_0_ready;
  wire         sinkVec_queue_40_deq_ready = sinkVec_sinkWire_40_ready;
  wire         sinkVec_queue_40_deq_valid;
  wire [4:0]   sinkVec_queue_40_deq_bits_vs;
  wire         sinkVec_20_0_valid = sinkVec_sinkWire_40_valid;
  wire [1:0]   sinkVec_queue_40_deq_bits_readSource;
  wire [4:0]   sinkVec_20_0_bits_vs = sinkVec_sinkWire_40_bits_vs;
  wire [1:0]   sinkVec_queue_40_deq_bits_offset;
  wire [1:0]   sinkVec_20_0_bits_readSource = sinkVec_sinkWire_40_bits_readSource;
  wire [2:0]   sinkVec_queue_40_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_20_0_bits_offset = sinkVec_sinkWire_40_bits_offset;
  wire [2:0]   sinkVec_20_0_bits_instructionIndex = sinkVec_sinkWire_40_bits_instructionIndex;
  wire         sinkVec_validSink_40_valid;
  wire [4:0]   sinkVec_validSink_40_bits_vs;
  wire [1:0]   sinkVec_validSink_40_bits_readSource;
  wire [1:0]   sinkVec_validSink_40_bits_offset;
  wire [2:0]   sinkVec_validSink_40_bits_instructionIndex;
  assign sinkVec_sinkWire_40_valid = sinkVec_queue_40_deq_valid;
  assign sinkVec_sinkWire_40_bits_vs = sinkVec_queue_40_deq_bits_vs;
  assign sinkVec_sinkWire_40_bits_readSource = sinkVec_queue_40_deq_bits_readSource;
  assign sinkVec_sinkWire_40_bits_offset = sinkVec_queue_40_deq_bits_offset;
  assign sinkVec_sinkWire_40_bits_instructionIndex = sinkVec_queue_40_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_40_enq_bits_offset;
  wire [2:0]   sinkVec_queue_40_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_40 = {sinkVec_queue_40_enq_bits_offset, sinkVec_queue_40_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_40_enq_bits_vs;
  wire [1:0]   sinkVec_queue_40_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_40 = {sinkVec_queue_40_enq_bits_vs, sinkVec_queue_40_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_40 = {sinkVec_queue_dataIn_hi_40, sinkVec_queue_dataIn_lo_40};
  wire [2:0]   sinkVec_queue_dataOut_40_instructionIndex = _sinkVec_queue_fifo_40_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_40_offset = _sinkVec_queue_fifo_40_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_40_readSource = _sinkVec_queue_fifo_40_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_40_vs = _sinkVec_queue_fifo_40_data_out[11:7];
  wire         sinkVec_queue_40_enq_ready = ~_sinkVec_queue_fifo_40_full;
  wire         sinkVec_queue_40_enq_valid;
  assign sinkVec_queue_40_deq_valid = ~_sinkVec_queue_fifo_40_empty | sinkVec_queue_40_enq_valid;
  assign sinkVec_queue_40_deq_bits_vs = _sinkVec_queue_fifo_40_empty ? sinkVec_queue_40_enq_bits_vs : sinkVec_queue_dataOut_40_vs;
  assign sinkVec_queue_40_deq_bits_readSource = _sinkVec_queue_fifo_40_empty ? sinkVec_queue_40_enq_bits_readSource : sinkVec_queue_dataOut_40_readSource;
  assign sinkVec_queue_40_deq_bits_offset = _sinkVec_queue_fifo_40_empty ? sinkVec_queue_40_enq_bits_offset : sinkVec_queue_dataOut_40_offset;
  assign sinkVec_queue_40_deq_bits_instructionIndex = _sinkVec_queue_fifo_40_empty ? sinkVec_queue_40_enq_bits_instructionIndex : sinkVec_queue_dataOut_40_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_40;
  wire         sinkVec_releasePipe_pipe_out_40_valid = sinkVec_releasePipe_pipe_v_40;
  wire         x13_10_0_ready;
  wire         x13_10_0_valid;
  wire         sinkVec_validSource_40_valid = x13_10_0_ready & x13_10_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_40;
  wire [2:0]   sinkVec_tokenCheck_counterChange_40 = sinkVec_validSource_40_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_40 = ~(sinkVec_tokenCheck_counter_40[2]);
  assign x13_10_0_ready = sinkVec_tokenCheck_40;
  assign sinkVec_queue_40_enq_valid = sinkVec_validSink_40_valid;
  assign sinkVec_queue_40_enq_bits_vs = sinkVec_validSink_40_bits_vs;
  assign sinkVec_queue_40_enq_bits_readSource = sinkVec_validSink_40_bits_readSource;
  assign sinkVec_queue_40_enq_bits_offset = sinkVec_validSink_40_bits_offset;
  assign sinkVec_queue_40_enq_bits_instructionIndex = sinkVec_validSink_40_bits_instructionIndex;
  reg          sinkVec_shifterReg_40_0_valid;
  assign sinkVec_validSink_40_valid = sinkVec_shifterReg_40_0_valid;
  reg  [4:0]   sinkVec_shifterReg_40_0_bits_vs;
  assign sinkVec_validSink_40_bits_vs = sinkVec_shifterReg_40_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_40_0_bits_readSource;
  assign sinkVec_validSink_40_bits_readSource = sinkVec_shifterReg_40_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_40_0_bits_offset;
  assign sinkVec_validSink_40_bits_offset = sinkVec_shifterReg_40_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_40_0_bits_instructionIndex;
  assign sinkVec_validSink_40_bits_instructionIndex = sinkVec_shifterReg_40_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_40 = sinkVec_shifterReg_40_0_valid | sinkVec_validSource_40_valid;
  wire         sinkVec_20_1_ready;
  wire         sinkVec_queue_41_deq_ready = sinkVec_sinkWire_41_ready;
  wire         sinkVec_queue_41_deq_valid;
  wire [4:0]   sinkVec_queue_41_deq_bits_vs;
  wire         sinkVec_20_1_valid = sinkVec_sinkWire_41_valid;
  wire [1:0]   sinkVec_queue_41_deq_bits_readSource;
  wire [4:0]   sinkVec_20_1_bits_vs = sinkVec_sinkWire_41_bits_vs;
  wire [1:0]   sinkVec_queue_41_deq_bits_offset;
  wire [1:0]   sinkVec_20_1_bits_readSource = sinkVec_sinkWire_41_bits_readSource;
  wire [2:0]   sinkVec_queue_41_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_20_1_bits_offset = sinkVec_sinkWire_41_bits_offset;
  wire [2:0]   sinkVec_20_1_bits_instructionIndex = sinkVec_sinkWire_41_bits_instructionIndex;
  wire         sinkVec_validSink_41_valid;
  wire [4:0]   sinkVec_validSink_41_bits_vs;
  wire [1:0]   sinkVec_validSink_41_bits_readSource;
  wire [1:0]   sinkVec_validSink_41_bits_offset;
  wire [2:0]   sinkVec_validSink_41_bits_instructionIndex;
  assign sinkVec_sinkWire_41_valid = sinkVec_queue_41_deq_valid;
  assign sinkVec_sinkWire_41_bits_vs = sinkVec_queue_41_deq_bits_vs;
  assign sinkVec_sinkWire_41_bits_readSource = sinkVec_queue_41_deq_bits_readSource;
  assign sinkVec_sinkWire_41_bits_offset = sinkVec_queue_41_deq_bits_offset;
  assign sinkVec_sinkWire_41_bits_instructionIndex = sinkVec_queue_41_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_41_enq_bits_offset;
  wire [2:0]   sinkVec_queue_41_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_41 = {sinkVec_queue_41_enq_bits_offset, sinkVec_queue_41_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_41_enq_bits_vs;
  wire [1:0]   sinkVec_queue_41_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_41 = {sinkVec_queue_41_enq_bits_vs, sinkVec_queue_41_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_41 = {sinkVec_queue_dataIn_hi_41, sinkVec_queue_dataIn_lo_41};
  wire [2:0]   sinkVec_queue_dataOut_41_instructionIndex = _sinkVec_queue_fifo_41_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_41_offset = _sinkVec_queue_fifo_41_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_41_readSource = _sinkVec_queue_fifo_41_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_41_vs = _sinkVec_queue_fifo_41_data_out[11:7];
  wire         sinkVec_queue_41_enq_ready = ~_sinkVec_queue_fifo_41_full;
  wire         sinkVec_queue_41_enq_valid;
  assign sinkVec_queue_41_deq_valid = ~_sinkVec_queue_fifo_41_empty | sinkVec_queue_41_enq_valid;
  assign sinkVec_queue_41_deq_bits_vs = _sinkVec_queue_fifo_41_empty ? sinkVec_queue_41_enq_bits_vs : sinkVec_queue_dataOut_41_vs;
  assign sinkVec_queue_41_deq_bits_readSource = _sinkVec_queue_fifo_41_empty ? sinkVec_queue_41_enq_bits_readSource : sinkVec_queue_dataOut_41_readSource;
  assign sinkVec_queue_41_deq_bits_offset = _sinkVec_queue_fifo_41_empty ? sinkVec_queue_41_enq_bits_offset : sinkVec_queue_dataOut_41_offset;
  assign sinkVec_queue_41_deq_bits_instructionIndex = _sinkVec_queue_fifo_41_empty ? sinkVec_queue_41_enq_bits_instructionIndex : sinkVec_queue_dataOut_41_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_41;
  wire         sinkVec_releasePipe_pipe_out_41_valid = sinkVec_releasePipe_pipe_v_41;
  wire         x13_10_1_ready;
  wire         x13_10_1_valid;
  wire         sinkVec_validSource_41_valid = x13_10_1_ready & x13_10_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_41;
  wire [2:0]   sinkVec_tokenCheck_counterChange_41 = sinkVec_validSource_41_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_41 = ~(sinkVec_tokenCheck_counter_41[2]);
  assign x13_10_1_ready = sinkVec_tokenCheck_41;
  assign sinkVec_queue_41_enq_valid = sinkVec_validSink_41_valid;
  assign sinkVec_queue_41_enq_bits_vs = sinkVec_validSink_41_bits_vs;
  assign sinkVec_queue_41_enq_bits_readSource = sinkVec_validSink_41_bits_readSource;
  assign sinkVec_queue_41_enq_bits_offset = sinkVec_validSink_41_bits_offset;
  assign sinkVec_queue_41_enq_bits_instructionIndex = sinkVec_validSink_41_bits_instructionIndex;
  reg          sinkVec_shifterReg_41_0_valid;
  assign sinkVec_validSink_41_valid = sinkVec_shifterReg_41_0_valid;
  reg  [4:0]   sinkVec_shifterReg_41_0_bits_vs;
  assign sinkVec_validSink_41_bits_vs = sinkVec_shifterReg_41_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_41_0_bits_readSource;
  assign sinkVec_validSink_41_bits_readSource = sinkVec_shifterReg_41_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_41_0_bits_offset;
  assign sinkVec_validSink_41_bits_offset = sinkVec_shifterReg_41_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_41_0_bits_instructionIndex;
  assign sinkVec_validSink_41_bits_instructionIndex = sinkVec_shifterReg_41_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_41 = sinkVec_shifterReg_41_0_valid | sinkVec_validSource_41_valid;
  assign sinkVec_sinkWire_40_ready = sinkVec_20_0_ready;
  assign sinkVec_sinkWire_41_ready = sinkVec_20_1_ready;
  reg          maskUnitFirst_20;
  wire         tryToRead_20 = sinkVec_20_0_valid | sinkVec_20_1_valid;
  wire         sinkWire_20_valid = maskUnitFirst_20 ? sinkVec_20_0_valid : sinkVec_20_1_valid;
  wire [4:0]   sinkWire_20_bits_vs = maskUnitFirst_20 ? sinkVec_20_0_bits_vs : sinkVec_20_1_bits_vs;
  wire [1:0]   sinkWire_20_bits_readSource = maskUnitFirst_20 ? sinkVec_20_0_bits_readSource : sinkVec_20_1_bits_readSource;
  wire [1:0]   sinkWire_20_bits_offset = maskUnitFirst_20 ? sinkVec_20_0_bits_offset : sinkVec_20_1_bits_offset;
  wire [2:0]   sinkWire_20_bits_instructionIndex = maskUnitFirst_20 ? sinkVec_20_0_bits_instructionIndex : sinkVec_20_1_bits_instructionIndex;
  wire         sinkWire_20_ready;
  assign sinkVec_20_1_ready = sinkWire_20_ready & ~maskUnitFirst_20;
  assign sinkVec_20_0_ready = sinkWire_20_ready & maskUnitFirst_20;
  reg          accessDataValid_pipe_v_20;
  reg          accessDataValid_pipe_pipe_v_20;
  wire         accessDataValid_pipe_pipe_out_20_valid = accessDataValid_pipe_pipe_v_20;
  wire         accessDataSource_20_valid = accessDataValid_pipe_pipe_out_20_valid;
  reg          shifterReg_36_0_valid;
  reg  [31:0]  shifterReg_36_0_bits;
  wire         shifterValid_36 = shifterReg_36_0_valid | accessDataSource_20_valid;
  reg          accessDataValid_pipe_v_21;
  reg          accessDataValid_pipe_pipe_v_21;
  wire         accessDataValid_pipe_pipe_out_21_valid = accessDataValid_pipe_pipe_v_21;
  wire         accessDataSource_21_valid = accessDataValid_pipe_pipe_out_21_valid;
  reg          shifterReg_37_0_valid;
  reg  [31:0]  shifterReg_37_0_bits;
  wire         shifterValid_37 = shifterReg_37_0_valid | accessDataSource_21_valid;
  wire         sinkVec_tokenCheck_42;
  wire [4:0]   sinkVec_validSource_42_bits_vd = x22_10_0_bits_vd;
  wire [1:0]   sinkVec_validSource_42_bits_offset = x22_10_0_bits_offset;
  wire [3:0]   sinkVec_validSource_42_bits_mask = x22_10_0_bits_mask;
  wire [31:0]  sinkVec_validSource_42_bits_data = x22_10_0_bits_data;
  wire [2:0]   sinkVec_validSource_42_bits_instructionIndex = x22_10_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_43;
  wire [4:0]   sinkVec_validSource_43_bits_vd = x22_10_1_bits_vd;
  wire [1:0]   sinkVec_validSource_43_bits_offset = x22_10_1_bits_offset;
  wire [3:0]   sinkVec_validSource_43_bits_mask = x22_10_1_bits_mask;
  wire [31:0]  sinkVec_validSource_43_bits_data = x22_10_1_bits_data;
  wire         sinkVec_validSource_43_bits_last = x22_10_1_bits_last;
  wire [2:0]   sinkVec_validSource_43_bits_instructionIndex = x22_10_1_bits_instructionIndex;
  wire         sinkVec_21_0_ready;
  wire         sinkVec_queue_42_deq_ready = sinkVec_sinkWire_42_ready;
  wire         sinkVec_queue_42_deq_valid;
  wire [4:0]   sinkVec_queue_42_deq_bits_vd;
  wire         sinkVec_21_0_valid = sinkVec_sinkWire_42_valid;
  wire [1:0]   sinkVec_queue_42_deq_bits_offset;
  wire [4:0]   sinkVec_21_0_bits_vd = sinkVec_sinkWire_42_bits_vd;
  wire [3:0]   sinkVec_queue_42_deq_bits_mask;
  wire [1:0]   sinkVec_21_0_bits_offset = sinkVec_sinkWire_42_bits_offset;
  wire [31:0]  sinkVec_queue_42_deq_bits_data;
  wire [3:0]   sinkVec_21_0_bits_mask = sinkVec_sinkWire_42_bits_mask;
  wire         sinkVec_queue_42_deq_bits_last;
  wire [31:0]  sinkVec_21_0_bits_data = sinkVec_sinkWire_42_bits_data;
  wire [2:0]   sinkVec_queue_42_deq_bits_instructionIndex;
  wire         sinkVec_21_0_bits_last = sinkVec_sinkWire_42_bits_last;
  wire [2:0]   sinkVec_21_0_bits_instructionIndex = sinkVec_sinkWire_42_bits_instructionIndex;
  wire         sinkVec_validSink_42_valid;
  wire [4:0]   sinkVec_validSink_42_bits_vd;
  wire [1:0]   sinkVec_validSink_42_bits_offset;
  wire [3:0]   sinkVec_validSink_42_bits_mask;
  wire [31:0]  sinkVec_validSink_42_bits_data;
  wire [2:0]   sinkVec_validSink_42_bits_instructionIndex;
  assign sinkVec_sinkWire_42_valid = sinkVec_queue_42_deq_valid;
  assign sinkVec_sinkWire_42_bits_vd = sinkVec_queue_42_deq_bits_vd;
  assign sinkVec_sinkWire_42_bits_offset = sinkVec_queue_42_deq_bits_offset;
  assign sinkVec_sinkWire_42_bits_mask = sinkVec_queue_42_deq_bits_mask;
  assign sinkVec_sinkWire_42_bits_data = sinkVec_queue_42_deq_bits_data;
  assign sinkVec_sinkWire_42_bits_last = sinkVec_queue_42_deq_bits_last;
  assign sinkVec_sinkWire_42_bits_instructionIndex = sinkVec_queue_42_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_42_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_20 = {sinkVec_queue_42_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_42_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_42 = {sinkVec_queue_dataIn_lo_hi_20, sinkVec_queue_42_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_42_enq_bits_vd;
  wire [1:0]   sinkVec_queue_42_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_20 = {sinkVec_queue_42_enq_bits_vd, sinkVec_queue_42_enq_bits_offset};
  wire [3:0]   sinkVec_queue_42_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_42 = {sinkVec_queue_dataIn_hi_hi_20, sinkVec_queue_42_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_42 = {sinkVec_queue_dataIn_hi_42, sinkVec_queue_dataIn_lo_42};
  wire [2:0]   sinkVec_queue_dataOut_42_instructionIndex = _sinkVec_queue_fifo_42_data_out[2:0];
  wire         sinkVec_queue_dataOut_42_last = _sinkVec_queue_fifo_42_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_42_data = _sinkVec_queue_fifo_42_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_42_mask = _sinkVec_queue_fifo_42_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_42_offset = _sinkVec_queue_fifo_42_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_42_vd = _sinkVec_queue_fifo_42_data_out[46:42];
  wire         sinkVec_queue_42_enq_ready = ~_sinkVec_queue_fifo_42_full;
  wire         sinkVec_queue_42_enq_valid;
  assign sinkVec_queue_42_deq_valid = ~_sinkVec_queue_fifo_42_empty | sinkVec_queue_42_enq_valid;
  assign sinkVec_queue_42_deq_bits_vd = _sinkVec_queue_fifo_42_empty ? sinkVec_queue_42_enq_bits_vd : sinkVec_queue_dataOut_42_vd;
  assign sinkVec_queue_42_deq_bits_offset = _sinkVec_queue_fifo_42_empty ? sinkVec_queue_42_enq_bits_offset : sinkVec_queue_dataOut_42_offset;
  assign sinkVec_queue_42_deq_bits_mask = _sinkVec_queue_fifo_42_empty ? sinkVec_queue_42_enq_bits_mask : sinkVec_queue_dataOut_42_mask;
  assign sinkVec_queue_42_deq_bits_data = _sinkVec_queue_fifo_42_empty ? sinkVec_queue_42_enq_bits_data : sinkVec_queue_dataOut_42_data;
  assign sinkVec_queue_42_deq_bits_last = ~_sinkVec_queue_fifo_42_empty & sinkVec_queue_dataOut_42_last;
  assign sinkVec_queue_42_deq_bits_instructionIndex = _sinkVec_queue_fifo_42_empty ? sinkVec_queue_42_enq_bits_instructionIndex : sinkVec_queue_dataOut_42_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_42;
  wire         sinkVec_releasePipe_pipe_out_42_valid = sinkVec_releasePipe_pipe_v_42;
  wire         x22_10_0_ready;
  wire         x22_10_0_valid;
  wire         sinkVec_validSource_42_valid = x22_10_0_ready & x22_10_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_42;
  wire [2:0]   sinkVec_tokenCheck_counterChange_42 = sinkVec_validSource_42_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_42 = ~(sinkVec_tokenCheck_counter_42[2]);
  assign x22_10_0_ready = sinkVec_tokenCheck_42;
  assign sinkVec_queue_42_enq_valid = sinkVec_validSink_42_valid;
  assign sinkVec_queue_42_enq_bits_vd = sinkVec_validSink_42_bits_vd;
  assign sinkVec_queue_42_enq_bits_offset = sinkVec_validSink_42_bits_offset;
  assign sinkVec_queue_42_enq_bits_mask = sinkVec_validSink_42_bits_mask;
  assign sinkVec_queue_42_enq_bits_data = sinkVec_validSink_42_bits_data;
  assign sinkVec_queue_42_enq_bits_instructionIndex = sinkVec_validSink_42_bits_instructionIndex;
  reg          sinkVec_shifterReg_42_0_valid;
  assign sinkVec_validSink_42_valid = sinkVec_shifterReg_42_0_valid;
  reg  [4:0]   sinkVec_shifterReg_42_0_bits_vd;
  assign sinkVec_validSink_42_bits_vd = sinkVec_shifterReg_42_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_42_0_bits_offset;
  assign sinkVec_validSink_42_bits_offset = sinkVec_shifterReg_42_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_42_0_bits_mask;
  assign sinkVec_validSink_42_bits_mask = sinkVec_shifterReg_42_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_42_0_bits_data;
  assign sinkVec_validSink_42_bits_data = sinkVec_shifterReg_42_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_42_0_bits_instructionIndex;
  assign sinkVec_validSink_42_bits_instructionIndex = sinkVec_shifterReg_42_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_42 = sinkVec_shifterReg_42_0_valid | sinkVec_validSource_42_valid;
  wire         sinkVec_21_1_ready;
  wire         sinkVec_queue_43_deq_ready = sinkVec_sinkWire_43_ready;
  wire         sinkVec_queue_43_deq_valid;
  wire [4:0]   sinkVec_queue_43_deq_bits_vd;
  wire         sinkVec_21_1_valid = sinkVec_sinkWire_43_valid;
  wire [1:0]   sinkVec_queue_43_deq_bits_offset;
  wire [4:0]   sinkVec_21_1_bits_vd = sinkVec_sinkWire_43_bits_vd;
  wire [3:0]   sinkVec_queue_43_deq_bits_mask;
  wire [1:0]   sinkVec_21_1_bits_offset = sinkVec_sinkWire_43_bits_offset;
  wire [31:0]  sinkVec_queue_43_deq_bits_data;
  wire [3:0]   sinkVec_21_1_bits_mask = sinkVec_sinkWire_43_bits_mask;
  wire         sinkVec_queue_43_deq_bits_last;
  wire [31:0]  sinkVec_21_1_bits_data = sinkVec_sinkWire_43_bits_data;
  wire [2:0]   sinkVec_queue_43_deq_bits_instructionIndex;
  wire         sinkVec_21_1_bits_last = sinkVec_sinkWire_43_bits_last;
  wire [2:0]   sinkVec_21_1_bits_instructionIndex = sinkVec_sinkWire_43_bits_instructionIndex;
  wire         sinkVec_validSink_43_valid;
  wire [4:0]   sinkVec_validSink_43_bits_vd;
  wire [1:0]   sinkVec_validSink_43_bits_offset;
  wire [3:0]   sinkVec_validSink_43_bits_mask;
  wire [31:0]  sinkVec_validSink_43_bits_data;
  wire         sinkVec_validSink_43_bits_last;
  wire [2:0]   sinkVec_validSink_43_bits_instructionIndex;
  assign sinkVec_sinkWire_43_valid = sinkVec_queue_43_deq_valid;
  assign sinkVec_sinkWire_43_bits_vd = sinkVec_queue_43_deq_bits_vd;
  assign sinkVec_sinkWire_43_bits_offset = sinkVec_queue_43_deq_bits_offset;
  assign sinkVec_sinkWire_43_bits_mask = sinkVec_queue_43_deq_bits_mask;
  assign sinkVec_sinkWire_43_bits_data = sinkVec_queue_43_deq_bits_data;
  assign sinkVec_sinkWire_43_bits_last = sinkVec_queue_43_deq_bits_last;
  assign sinkVec_sinkWire_43_bits_instructionIndex = sinkVec_queue_43_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_43_enq_bits_data;
  wire         sinkVec_queue_43_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_21 = {sinkVec_queue_43_enq_bits_data, sinkVec_queue_43_enq_bits_last};
  wire [2:0]   sinkVec_queue_43_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_43 = {sinkVec_queue_dataIn_lo_hi_21, sinkVec_queue_43_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_43_enq_bits_vd;
  wire [1:0]   sinkVec_queue_43_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_21 = {sinkVec_queue_43_enq_bits_vd, sinkVec_queue_43_enq_bits_offset};
  wire [3:0]   sinkVec_queue_43_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_43 = {sinkVec_queue_dataIn_hi_hi_21, sinkVec_queue_43_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_43 = {sinkVec_queue_dataIn_hi_43, sinkVec_queue_dataIn_lo_43};
  wire [2:0]   sinkVec_queue_dataOut_43_instructionIndex = _sinkVec_queue_fifo_43_data_out[2:0];
  wire         sinkVec_queue_dataOut_43_last = _sinkVec_queue_fifo_43_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_43_data = _sinkVec_queue_fifo_43_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_43_mask = _sinkVec_queue_fifo_43_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_43_offset = _sinkVec_queue_fifo_43_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_43_vd = _sinkVec_queue_fifo_43_data_out[46:42];
  wire         sinkVec_queue_43_enq_ready = ~_sinkVec_queue_fifo_43_full;
  wire         sinkVec_queue_43_enq_valid;
  assign sinkVec_queue_43_deq_valid = ~_sinkVec_queue_fifo_43_empty | sinkVec_queue_43_enq_valid;
  assign sinkVec_queue_43_deq_bits_vd = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_vd : sinkVec_queue_dataOut_43_vd;
  assign sinkVec_queue_43_deq_bits_offset = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_offset : sinkVec_queue_dataOut_43_offset;
  assign sinkVec_queue_43_deq_bits_mask = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_mask : sinkVec_queue_dataOut_43_mask;
  assign sinkVec_queue_43_deq_bits_data = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_data : sinkVec_queue_dataOut_43_data;
  assign sinkVec_queue_43_deq_bits_last = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_last : sinkVec_queue_dataOut_43_last;
  assign sinkVec_queue_43_deq_bits_instructionIndex = _sinkVec_queue_fifo_43_empty ? sinkVec_queue_43_enq_bits_instructionIndex : sinkVec_queue_dataOut_43_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_43;
  wire         sinkVec_releasePipe_pipe_out_43_valid = sinkVec_releasePipe_pipe_v_43;
  wire         x22_10_1_ready;
  wire         x22_10_1_valid;
  wire         sinkVec_validSource_43_valid = x22_10_1_ready & x22_10_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_43;
  wire [2:0]   sinkVec_tokenCheck_counterChange_43 = sinkVec_validSource_43_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_43 = ~(sinkVec_tokenCheck_counter_43[2]);
  assign x22_10_1_ready = sinkVec_tokenCheck_43;
  assign sinkVec_queue_43_enq_valid = sinkVec_validSink_43_valid;
  assign sinkVec_queue_43_enq_bits_vd = sinkVec_validSink_43_bits_vd;
  assign sinkVec_queue_43_enq_bits_offset = sinkVec_validSink_43_bits_offset;
  assign sinkVec_queue_43_enq_bits_mask = sinkVec_validSink_43_bits_mask;
  assign sinkVec_queue_43_enq_bits_data = sinkVec_validSink_43_bits_data;
  assign sinkVec_queue_43_enq_bits_last = sinkVec_validSink_43_bits_last;
  assign sinkVec_queue_43_enq_bits_instructionIndex = sinkVec_validSink_43_bits_instructionIndex;
  reg          sinkVec_shifterReg_43_0_valid;
  assign sinkVec_validSink_43_valid = sinkVec_shifterReg_43_0_valid;
  reg  [4:0]   sinkVec_shifterReg_43_0_bits_vd;
  assign sinkVec_validSink_43_bits_vd = sinkVec_shifterReg_43_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_43_0_bits_offset;
  assign sinkVec_validSink_43_bits_offset = sinkVec_shifterReg_43_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_43_0_bits_mask;
  assign sinkVec_validSink_43_bits_mask = sinkVec_shifterReg_43_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_43_0_bits_data;
  assign sinkVec_validSink_43_bits_data = sinkVec_shifterReg_43_0_bits_data;
  reg          sinkVec_shifterReg_43_0_bits_last;
  assign sinkVec_validSink_43_bits_last = sinkVec_shifterReg_43_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_43_0_bits_instructionIndex;
  assign sinkVec_validSink_43_bits_instructionIndex = sinkVec_shifterReg_43_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_43 = sinkVec_shifterReg_43_0_valid | sinkVec_validSource_43_valid;
  assign sinkVec_sinkWire_42_ready = sinkVec_21_0_ready;
  assign sinkVec_sinkWire_43_ready = sinkVec_21_1_ready;
  reg          maskUnitFirst_21;
  wire         tryToRead_21 = sinkVec_21_0_valid | sinkVec_21_1_valid;
  wire         sinkWire_21_valid = maskUnitFirst_21 ? sinkVec_21_0_valid : sinkVec_21_1_valid;
  wire [4:0]   sinkWire_21_bits_vd = maskUnitFirst_21 ? sinkVec_21_0_bits_vd : sinkVec_21_1_bits_vd;
  wire [1:0]   sinkWire_21_bits_offset = maskUnitFirst_21 ? sinkVec_21_0_bits_offset : sinkVec_21_1_bits_offset;
  wire [3:0]   sinkWire_21_bits_mask = maskUnitFirst_21 ? sinkVec_21_0_bits_mask : sinkVec_21_1_bits_mask;
  wire [31:0]  sinkWire_21_bits_data = maskUnitFirst_21 ? sinkVec_21_0_bits_data : sinkVec_21_1_bits_data;
  wire         sinkWire_21_bits_last = maskUnitFirst_21 ? sinkVec_21_0_bits_last : sinkVec_21_1_bits_last;
  wire [2:0]   sinkWire_21_bits_instructionIndex = maskUnitFirst_21 ? sinkVec_21_0_bits_instructionIndex : sinkVec_21_1_bits_instructionIndex;
  wire         sinkWire_21_ready;
  assign sinkVec_21_1_ready = sinkWire_21_ready & ~maskUnitFirst_21;
  assign sinkVec_21_0_ready = sinkWire_21_ready & maskUnitFirst_21;
  reg          view__writeRelease_10_pipe_v;
  wire         view__writeRelease_10_pipe_out_valid = view__writeRelease_10_pipe_v;
  reg          pipe_v_30;
  wire         pipe_out_20_valid = pipe_v_30;
  wire         _probeWire_writeQueueEnqVec_10_valid_T = x22_10_0_ready & _maskUnit_exeResp_10_valid;
  reg          instructionFinishedPipe_pipe_v_10;
  wire         instructionFinishedPipe_pipe_out_10_valid = instructionFinishedPipe_pipe_v_10;
  reg  [7:0]   instructionFinishedPipe_pipe_b_10;
  wire [7:0]   instructionFinishedPipe_pipe_out_10_bits = instructionFinishedPipe_pipe_b_10;
  wire         instructionFinished_10_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_10_bits);
  wire         instructionFinished_10_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_10_bits);
  wire         instructionFinished_10_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_10_bits);
  wire         instructionFinished_10_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_10_bits);
  assign vxsatReportVec_10 = _laneVec_10_vxsatReport[3:0];
  reg          pipe_v_31;
  reg  [31:0]  pipe_b_31;
  reg          pipe_pipe_v_10;
  wire         pipe_pipe_out_10_valid = pipe_pipe_v_10;
  reg  [31:0]  pipe_pipe_b_10;
  wire [31:0]  pipe_pipe_out_10_bits = pipe_pipe_b_10;
  reg          view__laneMaskSelect_10_pipe_v;
  reg  [5:0]   view__laneMaskSelect_10_pipe_b;
  reg          view__laneMaskSelect_10_pipe_pipe_v;
  wire         view__laneMaskSelect_10_pipe_pipe_out_valid = view__laneMaskSelect_10_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_10_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_10_pipe_pipe_out_bits = view__laneMaskSelect_10_pipe_pipe_b;
  reg          view__laneMaskSewSelect_10_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_10_pipe_b;
  reg          view__laneMaskSewSelect_10_pipe_pipe_v;
  wire         view__laneMaskSewSelect_10_pipe_pipe_out_valid = view__laneMaskSewSelect_10_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_10_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_10_pipe_pipe_out_bits = view__laneMaskSewSelect_10_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_10;
  wire         lsuLastPipe_pipe_out_10_valid = lsuLastPipe_pipe_v_10;
  reg  [7:0]   lsuLastPipe_pipe_b_10;
  wire [7:0]   lsuLastPipe_pipe_out_10_bits = lsuLastPipe_pipe_b_10;
  reg          maskLastPipe_pipe_v_10;
  wire         maskLastPipe_pipe_out_10_valid = maskLastPipe_pipe_v_10;
  reg  [7:0]   maskLastPipe_pipe_b_10;
  wire [7:0]   maskLastPipe_pipe_out_10_bits = maskLastPipe_pipe_b_10;
  wire [5:0]   writeCounter_10 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h28};
  reg          pipe_v_32;
  wire         pipe_out_21_valid = pipe_v_32;
  reg  [5:0]   pipe_b_32;
  wire [5:0]   pipe_out_21_bits = pipe_b_32;
  assign laneRequestSinkWire_11_ready = ~laneRequestSinkWire_11_bits_issueInst | _laneVec_11_laneRequest_ready;
  wire         sinkVec_tokenCheck_44;
  wire [4:0]   sinkVec_validSource_44_bits_vs = x13_11_0_bits_vs;
  wire [1:0]   sinkVec_validSource_44_bits_offset = x13_11_0_bits_offset;
  wire [2:0]   sinkVec_validSource_44_bits_instructionIndex = x13_11_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_45;
  wire [4:0]   sinkVec_validSource_45_bits_vs = x13_11_1_bits_vs;
  wire [1:0]   sinkVec_validSource_45_bits_offset = x13_11_1_bits_offset;
  wire [2:0]   sinkVec_validSource_45_bits_instructionIndex = x13_11_1_bits_instructionIndex;
  wire         sinkVec_22_0_ready;
  wire         sinkVec_queue_44_deq_ready = sinkVec_sinkWire_44_ready;
  wire         sinkVec_queue_44_deq_valid;
  wire [4:0]   sinkVec_queue_44_deq_bits_vs;
  wire         sinkVec_22_0_valid = sinkVec_sinkWire_44_valid;
  wire [1:0]   sinkVec_queue_44_deq_bits_readSource;
  wire [4:0]   sinkVec_22_0_bits_vs = sinkVec_sinkWire_44_bits_vs;
  wire [1:0]   sinkVec_queue_44_deq_bits_offset;
  wire [1:0]   sinkVec_22_0_bits_readSource = sinkVec_sinkWire_44_bits_readSource;
  wire [2:0]   sinkVec_queue_44_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_22_0_bits_offset = sinkVec_sinkWire_44_bits_offset;
  wire [2:0]   sinkVec_22_0_bits_instructionIndex = sinkVec_sinkWire_44_bits_instructionIndex;
  wire         sinkVec_validSink_44_valid;
  wire [4:0]   sinkVec_validSink_44_bits_vs;
  wire [1:0]   sinkVec_validSink_44_bits_readSource;
  wire [1:0]   sinkVec_validSink_44_bits_offset;
  wire [2:0]   sinkVec_validSink_44_bits_instructionIndex;
  assign sinkVec_sinkWire_44_valid = sinkVec_queue_44_deq_valid;
  assign sinkVec_sinkWire_44_bits_vs = sinkVec_queue_44_deq_bits_vs;
  assign sinkVec_sinkWire_44_bits_readSource = sinkVec_queue_44_deq_bits_readSource;
  assign sinkVec_sinkWire_44_bits_offset = sinkVec_queue_44_deq_bits_offset;
  assign sinkVec_sinkWire_44_bits_instructionIndex = sinkVec_queue_44_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_44_enq_bits_offset;
  wire [2:0]   sinkVec_queue_44_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_44 = {sinkVec_queue_44_enq_bits_offset, sinkVec_queue_44_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_44_enq_bits_vs;
  wire [1:0]   sinkVec_queue_44_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_44 = {sinkVec_queue_44_enq_bits_vs, sinkVec_queue_44_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_44 = {sinkVec_queue_dataIn_hi_44, sinkVec_queue_dataIn_lo_44};
  wire [2:0]   sinkVec_queue_dataOut_44_instructionIndex = _sinkVec_queue_fifo_44_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_44_offset = _sinkVec_queue_fifo_44_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_44_readSource = _sinkVec_queue_fifo_44_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_44_vs = _sinkVec_queue_fifo_44_data_out[11:7];
  wire         sinkVec_queue_44_enq_ready = ~_sinkVec_queue_fifo_44_full;
  wire         sinkVec_queue_44_enq_valid;
  assign sinkVec_queue_44_deq_valid = ~_sinkVec_queue_fifo_44_empty | sinkVec_queue_44_enq_valid;
  assign sinkVec_queue_44_deq_bits_vs = _sinkVec_queue_fifo_44_empty ? sinkVec_queue_44_enq_bits_vs : sinkVec_queue_dataOut_44_vs;
  assign sinkVec_queue_44_deq_bits_readSource = _sinkVec_queue_fifo_44_empty ? sinkVec_queue_44_enq_bits_readSource : sinkVec_queue_dataOut_44_readSource;
  assign sinkVec_queue_44_deq_bits_offset = _sinkVec_queue_fifo_44_empty ? sinkVec_queue_44_enq_bits_offset : sinkVec_queue_dataOut_44_offset;
  assign sinkVec_queue_44_deq_bits_instructionIndex = _sinkVec_queue_fifo_44_empty ? sinkVec_queue_44_enq_bits_instructionIndex : sinkVec_queue_dataOut_44_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_44;
  wire         sinkVec_releasePipe_pipe_out_44_valid = sinkVec_releasePipe_pipe_v_44;
  wire         x13_11_0_ready;
  wire         x13_11_0_valid;
  wire         sinkVec_validSource_44_valid = x13_11_0_ready & x13_11_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_44;
  wire [2:0]   sinkVec_tokenCheck_counterChange_44 = sinkVec_validSource_44_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_44 = ~(sinkVec_tokenCheck_counter_44[2]);
  assign x13_11_0_ready = sinkVec_tokenCheck_44;
  assign sinkVec_queue_44_enq_valid = sinkVec_validSink_44_valid;
  assign sinkVec_queue_44_enq_bits_vs = sinkVec_validSink_44_bits_vs;
  assign sinkVec_queue_44_enq_bits_readSource = sinkVec_validSink_44_bits_readSource;
  assign sinkVec_queue_44_enq_bits_offset = sinkVec_validSink_44_bits_offset;
  assign sinkVec_queue_44_enq_bits_instructionIndex = sinkVec_validSink_44_bits_instructionIndex;
  reg          sinkVec_shifterReg_44_0_valid;
  assign sinkVec_validSink_44_valid = sinkVec_shifterReg_44_0_valid;
  reg  [4:0]   sinkVec_shifterReg_44_0_bits_vs;
  assign sinkVec_validSink_44_bits_vs = sinkVec_shifterReg_44_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_44_0_bits_readSource;
  assign sinkVec_validSink_44_bits_readSource = sinkVec_shifterReg_44_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_44_0_bits_offset;
  assign sinkVec_validSink_44_bits_offset = sinkVec_shifterReg_44_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_44_0_bits_instructionIndex;
  assign sinkVec_validSink_44_bits_instructionIndex = sinkVec_shifterReg_44_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_44 = sinkVec_shifterReg_44_0_valid | sinkVec_validSource_44_valid;
  wire         sinkVec_22_1_ready;
  wire         sinkVec_queue_45_deq_ready = sinkVec_sinkWire_45_ready;
  wire         sinkVec_queue_45_deq_valid;
  wire [4:0]   sinkVec_queue_45_deq_bits_vs;
  wire         sinkVec_22_1_valid = sinkVec_sinkWire_45_valid;
  wire [1:0]   sinkVec_queue_45_deq_bits_readSource;
  wire [4:0]   sinkVec_22_1_bits_vs = sinkVec_sinkWire_45_bits_vs;
  wire [1:0]   sinkVec_queue_45_deq_bits_offset;
  wire [1:0]   sinkVec_22_1_bits_readSource = sinkVec_sinkWire_45_bits_readSource;
  wire [2:0]   sinkVec_queue_45_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_22_1_bits_offset = sinkVec_sinkWire_45_bits_offset;
  wire [2:0]   sinkVec_22_1_bits_instructionIndex = sinkVec_sinkWire_45_bits_instructionIndex;
  wire         sinkVec_validSink_45_valid;
  wire [4:0]   sinkVec_validSink_45_bits_vs;
  wire [1:0]   sinkVec_validSink_45_bits_readSource;
  wire [1:0]   sinkVec_validSink_45_bits_offset;
  wire [2:0]   sinkVec_validSink_45_bits_instructionIndex;
  assign sinkVec_sinkWire_45_valid = sinkVec_queue_45_deq_valid;
  assign sinkVec_sinkWire_45_bits_vs = sinkVec_queue_45_deq_bits_vs;
  assign sinkVec_sinkWire_45_bits_readSource = sinkVec_queue_45_deq_bits_readSource;
  assign sinkVec_sinkWire_45_bits_offset = sinkVec_queue_45_deq_bits_offset;
  assign sinkVec_sinkWire_45_bits_instructionIndex = sinkVec_queue_45_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_45_enq_bits_offset;
  wire [2:0]   sinkVec_queue_45_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_45 = {sinkVec_queue_45_enq_bits_offset, sinkVec_queue_45_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_45_enq_bits_vs;
  wire [1:0]   sinkVec_queue_45_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_45 = {sinkVec_queue_45_enq_bits_vs, sinkVec_queue_45_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_45 = {sinkVec_queue_dataIn_hi_45, sinkVec_queue_dataIn_lo_45};
  wire [2:0]   sinkVec_queue_dataOut_45_instructionIndex = _sinkVec_queue_fifo_45_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_45_offset = _sinkVec_queue_fifo_45_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_45_readSource = _sinkVec_queue_fifo_45_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_45_vs = _sinkVec_queue_fifo_45_data_out[11:7];
  wire         sinkVec_queue_45_enq_ready = ~_sinkVec_queue_fifo_45_full;
  wire         sinkVec_queue_45_enq_valid;
  assign sinkVec_queue_45_deq_valid = ~_sinkVec_queue_fifo_45_empty | sinkVec_queue_45_enq_valid;
  assign sinkVec_queue_45_deq_bits_vs = _sinkVec_queue_fifo_45_empty ? sinkVec_queue_45_enq_bits_vs : sinkVec_queue_dataOut_45_vs;
  assign sinkVec_queue_45_deq_bits_readSource = _sinkVec_queue_fifo_45_empty ? sinkVec_queue_45_enq_bits_readSource : sinkVec_queue_dataOut_45_readSource;
  assign sinkVec_queue_45_deq_bits_offset = _sinkVec_queue_fifo_45_empty ? sinkVec_queue_45_enq_bits_offset : sinkVec_queue_dataOut_45_offset;
  assign sinkVec_queue_45_deq_bits_instructionIndex = _sinkVec_queue_fifo_45_empty ? sinkVec_queue_45_enq_bits_instructionIndex : sinkVec_queue_dataOut_45_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_45;
  wire         sinkVec_releasePipe_pipe_out_45_valid = sinkVec_releasePipe_pipe_v_45;
  wire         x13_11_1_ready;
  wire         x13_11_1_valid;
  wire         sinkVec_validSource_45_valid = x13_11_1_ready & x13_11_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_45;
  wire [2:0]   sinkVec_tokenCheck_counterChange_45 = sinkVec_validSource_45_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_45 = ~(sinkVec_tokenCheck_counter_45[2]);
  assign x13_11_1_ready = sinkVec_tokenCheck_45;
  assign sinkVec_queue_45_enq_valid = sinkVec_validSink_45_valid;
  assign sinkVec_queue_45_enq_bits_vs = sinkVec_validSink_45_bits_vs;
  assign sinkVec_queue_45_enq_bits_readSource = sinkVec_validSink_45_bits_readSource;
  assign sinkVec_queue_45_enq_bits_offset = sinkVec_validSink_45_bits_offset;
  assign sinkVec_queue_45_enq_bits_instructionIndex = sinkVec_validSink_45_bits_instructionIndex;
  reg          sinkVec_shifterReg_45_0_valid;
  assign sinkVec_validSink_45_valid = sinkVec_shifterReg_45_0_valid;
  reg  [4:0]   sinkVec_shifterReg_45_0_bits_vs;
  assign sinkVec_validSink_45_bits_vs = sinkVec_shifterReg_45_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_45_0_bits_readSource;
  assign sinkVec_validSink_45_bits_readSource = sinkVec_shifterReg_45_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_45_0_bits_offset;
  assign sinkVec_validSink_45_bits_offset = sinkVec_shifterReg_45_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_45_0_bits_instructionIndex;
  assign sinkVec_validSink_45_bits_instructionIndex = sinkVec_shifterReg_45_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_45 = sinkVec_shifterReg_45_0_valid | sinkVec_validSource_45_valid;
  assign sinkVec_sinkWire_44_ready = sinkVec_22_0_ready;
  assign sinkVec_sinkWire_45_ready = sinkVec_22_1_ready;
  reg          maskUnitFirst_22;
  wire         tryToRead_22 = sinkVec_22_0_valid | sinkVec_22_1_valid;
  wire         sinkWire_22_valid = maskUnitFirst_22 ? sinkVec_22_0_valid : sinkVec_22_1_valid;
  wire [4:0]   sinkWire_22_bits_vs = maskUnitFirst_22 ? sinkVec_22_0_bits_vs : sinkVec_22_1_bits_vs;
  wire [1:0]   sinkWire_22_bits_readSource = maskUnitFirst_22 ? sinkVec_22_0_bits_readSource : sinkVec_22_1_bits_readSource;
  wire [1:0]   sinkWire_22_bits_offset = maskUnitFirst_22 ? sinkVec_22_0_bits_offset : sinkVec_22_1_bits_offset;
  wire [2:0]   sinkWire_22_bits_instructionIndex = maskUnitFirst_22 ? sinkVec_22_0_bits_instructionIndex : sinkVec_22_1_bits_instructionIndex;
  wire         sinkWire_22_ready;
  assign sinkVec_22_1_ready = sinkWire_22_ready & ~maskUnitFirst_22;
  assign sinkVec_22_0_ready = sinkWire_22_ready & maskUnitFirst_22;
  reg          accessDataValid_pipe_v_22;
  reg          accessDataValid_pipe_pipe_v_22;
  wire         accessDataValid_pipe_pipe_out_22_valid = accessDataValid_pipe_pipe_v_22;
  wire         accessDataSource_22_valid = accessDataValid_pipe_pipe_out_22_valid;
  reg          shifterReg_38_0_valid;
  reg  [31:0]  shifterReg_38_0_bits;
  wire         shifterValid_38 = shifterReg_38_0_valid | accessDataSource_22_valid;
  reg          accessDataValid_pipe_v_23;
  reg          accessDataValid_pipe_pipe_v_23;
  wire         accessDataValid_pipe_pipe_out_23_valid = accessDataValid_pipe_pipe_v_23;
  wire         accessDataSource_23_valid = accessDataValid_pipe_pipe_out_23_valid;
  reg          shifterReg_39_0_valid;
  reg  [31:0]  shifterReg_39_0_bits;
  wire         shifterValid_39 = shifterReg_39_0_valid | accessDataSource_23_valid;
  wire         sinkVec_tokenCheck_46;
  wire [4:0]   sinkVec_validSource_46_bits_vd = x22_11_0_bits_vd;
  wire [1:0]   sinkVec_validSource_46_bits_offset = x22_11_0_bits_offset;
  wire [3:0]   sinkVec_validSource_46_bits_mask = x22_11_0_bits_mask;
  wire [31:0]  sinkVec_validSource_46_bits_data = x22_11_0_bits_data;
  wire [2:0]   sinkVec_validSource_46_bits_instructionIndex = x22_11_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_47;
  wire [4:0]   sinkVec_validSource_47_bits_vd = x22_11_1_bits_vd;
  wire [1:0]   sinkVec_validSource_47_bits_offset = x22_11_1_bits_offset;
  wire [3:0]   sinkVec_validSource_47_bits_mask = x22_11_1_bits_mask;
  wire [31:0]  sinkVec_validSource_47_bits_data = x22_11_1_bits_data;
  wire         sinkVec_validSource_47_bits_last = x22_11_1_bits_last;
  wire [2:0]   sinkVec_validSource_47_bits_instructionIndex = x22_11_1_bits_instructionIndex;
  wire         sinkVec_23_0_ready;
  wire         sinkVec_queue_46_deq_ready = sinkVec_sinkWire_46_ready;
  wire         sinkVec_queue_46_deq_valid;
  wire [4:0]   sinkVec_queue_46_deq_bits_vd;
  wire         sinkVec_23_0_valid = sinkVec_sinkWire_46_valid;
  wire [1:0]   sinkVec_queue_46_deq_bits_offset;
  wire [4:0]   sinkVec_23_0_bits_vd = sinkVec_sinkWire_46_bits_vd;
  wire [3:0]   sinkVec_queue_46_deq_bits_mask;
  wire [1:0]   sinkVec_23_0_bits_offset = sinkVec_sinkWire_46_bits_offset;
  wire [31:0]  sinkVec_queue_46_deq_bits_data;
  wire [3:0]   sinkVec_23_0_bits_mask = sinkVec_sinkWire_46_bits_mask;
  wire         sinkVec_queue_46_deq_bits_last;
  wire [31:0]  sinkVec_23_0_bits_data = sinkVec_sinkWire_46_bits_data;
  wire [2:0]   sinkVec_queue_46_deq_bits_instructionIndex;
  wire         sinkVec_23_0_bits_last = sinkVec_sinkWire_46_bits_last;
  wire [2:0]   sinkVec_23_0_bits_instructionIndex = sinkVec_sinkWire_46_bits_instructionIndex;
  wire         sinkVec_validSink_46_valid;
  wire [4:0]   sinkVec_validSink_46_bits_vd;
  wire [1:0]   sinkVec_validSink_46_bits_offset;
  wire [3:0]   sinkVec_validSink_46_bits_mask;
  wire [31:0]  sinkVec_validSink_46_bits_data;
  wire [2:0]   sinkVec_validSink_46_bits_instructionIndex;
  assign sinkVec_sinkWire_46_valid = sinkVec_queue_46_deq_valid;
  assign sinkVec_sinkWire_46_bits_vd = sinkVec_queue_46_deq_bits_vd;
  assign sinkVec_sinkWire_46_bits_offset = sinkVec_queue_46_deq_bits_offset;
  assign sinkVec_sinkWire_46_bits_mask = sinkVec_queue_46_deq_bits_mask;
  assign sinkVec_sinkWire_46_bits_data = sinkVec_queue_46_deq_bits_data;
  assign sinkVec_sinkWire_46_bits_last = sinkVec_queue_46_deq_bits_last;
  assign sinkVec_sinkWire_46_bits_instructionIndex = sinkVec_queue_46_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_46_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_22 = {sinkVec_queue_46_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_46_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_46 = {sinkVec_queue_dataIn_lo_hi_22, sinkVec_queue_46_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_46_enq_bits_vd;
  wire [1:0]   sinkVec_queue_46_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_22 = {sinkVec_queue_46_enq_bits_vd, sinkVec_queue_46_enq_bits_offset};
  wire [3:0]   sinkVec_queue_46_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_46 = {sinkVec_queue_dataIn_hi_hi_22, sinkVec_queue_46_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_46 = {sinkVec_queue_dataIn_hi_46, sinkVec_queue_dataIn_lo_46};
  wire [2:0]   sinkVec_queue_dataOut_46_instructionIndex = _sinkVec_queue_fifo_46_data_out[2:0];
  wire         sinkVec_queue_dataOut_46_last = _sinkVec_queue_fifo_46_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_46_data = _sinkVec_queue_fifo_46_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_46_mask = _sinkVec_queue_fifo_46_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_46_offset = _sinkVec_queue_fifo_46_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_46_vd = _sinkVec_queue_fifo_46_data_out[46:42];
  wire         sinkVec_queue_46_enq_ready = ~_sinkVec_queue_fifo_46_full;
  wire         sinkVec_queue_46_enq_valid;
  assign sinkVec_queue_46_deq_valid = ~_sinkVec_queue_fifo_46_empty | sinkVec_queue_46_enq_valid;
  assign sinkVec_queue_46_deq_bits_vd = _sinkVec_queue_fifo_46_empty ? sinkVec_queue_46_enq_bits_vd : sinkVec_queue_dataOut_46_vd;
  assign sinkVec_queue_46_deq_bits_offset = _sinkVec_queue_fifo_46_empty ? sinkVec_queue_46_enq_bits_offset : sinkVec_queue_dataOut_46_offset;
  assign sinkVec_queue_46_deq_bits_mask = _sinkVec_queue_fifo_46_empty ? sinkVec_queue_46_enq_bits_mask : sinkVec_queue_dataOut_46_mask;
  assign sinkVec_queue_46_deq_bits_data = _sinkVec_queue_fifo_46_empty ? sinkVec_queue_46_enq_bits_data : sinkVec_queue_dataOut_46_data;
  assign sinkVec_queue_46_deq_bits_last = ~_sinkVec_queue_fifo_46_empty & sinkVec_queue_dataOut_46_last;
  assign sinkVec_queue_46_deq_bits_instructionIndex = _sinkVec_queue_fifo_46_empty ? sinkVec_queue_46_enq_bits_instructionIndex : sinkVec_queue_dataOut_46_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_46;
  wire         sinkVec_releasePipe_pipe_out_46_valid = sinkVec_releasePipe_pipe_v_46;
  wire         x22_11_0_ready;
  wire         x22_11_0_valid;
  wire         sinkVec_validSource_46_valid = x22_11_0_ready & x22_11_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_46;
  wire [2:0]   sinkVec_tokenCheck_counterChange_46 = sinkVec_validSource_46_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_46 = ~(sinkVec_tokenCheck_counter_46[2]);
  assign x22_11_0_ready = sinkVec_tokenCheck_46;
  assign sinkVec_queue_46_enq_valid = sinkVec_validSink_46_valid;
  assign sinkVec_queue_46_enq_bits_vd = sinkVec_validSink_46_bits_vd;
  assign sinkVec_queue_46_enq_bits_offset = sinkVec_validSink_46_bits_offset;
  assign sinkVec_queue_46_enq_bits_mask = sinkVec_validSink_46_bits_mask;
  assign sinkVec_queue_46_enq_bits_data = sinkVec_validSink_46_bits_data;
  assign sinkVec_queue_46_enq_bits_instructionIndex = sinkVec_validSink_46_bits_instructionIndex;
  reg          sinkVec_shifterReg_46_0_valid;
  assign sinkVec_validSink_46_valid = sinkVec_shifterReg_46_0_valid;
  reg  [4:0]   sinkVec_shifterReg_46_0_bits_vd;
  assign sinkVec_validSink_46_bits_vd = sinkVec_shifterReg_46_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_46_0_bits_offset;
  assign sinkVec_validSink_46_bits_offset = sinkVec_shifterReg_46_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_46_0_bits_mask;
  assign sinkVec_validSink_46_bits_mask = sinkVec_shifterReg_46_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_46_0_bits_data;
  assign sinkVec_validSink_46_bits_data = sinkVec_shifterReg_46_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_46_0_bits_instructionIndex;
  assign sinkVec_validSink_46_bits_instructionIndex = sinkVec_shifterReg_46_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_46 = sinkVec_shifterReg_46_0_valid | sinkVec_validSource_46_valid;
  wire         sinkVec_23_1_ready;
  wire         sinkVec_queue_47_deq_ready = sinkVec_sinkWire_47_ready;
  wire         sinkVec_queue_47_deq_valid;
  wire [4:0]   sinkVec_queue_47_deq_bits_vd;
  wire         sinkVec_23_1_valid = sinkVec_sinkWire_47_valid;
  wire [1:0]   sinkVec_queue_47_deq_bits_offset;
  wire [4:0]   sinkVec_23_1_bits_vd = sinkVec_sinkWire_47_bits_vd;
  wire [3:0]   sinkVec_queue_47_deq_bits_mask;
  wire [1:0]   sinkVec_23_1_bits_offset = sinkVec_sinkWire_47_bits_offset;
  wire [31:0]  sinkVec_queue_47_deq_bits_data;
  wire [3:0]   sinkVec_23_1_bits_mask = sinkVec_sinkWire_47_bits_mask;
  wire         sinkVec_queue_47_deq_bits_last;
  wire [31:0]  sinkVec_23_1_bits_data = sinkVec_sinkWire_47_bits_data;
  wire [2:0]   sinkVec_queue_47_deq_bits_instructionIndex;
  wire         sinkVec_23_1_bits_last = sinkVec_sinkWire_47_bits_last;
  wire [2:0]   sinkVec_23_1_bits_instructionIndex = sinkVec_sinkWire_47_bits_instructionIndex;
  wire         sinkVec_validSink_47_valid;
  wire [4:0]   sinkVec_validSink_47_bits_vd;
  wire [1:0]   sinkVec_validSink_47_bits_offset;
  wire [3:0]   sinkVec_validSink_47_bits_mask;
  wire [31:0]  sinkVec_validSink_47_bits_data;
  wire         sinkVec_validSink_47_bits_last;
  wire [2:0]   sinkVec_validSink_47_bits_instructionIndex;
  assign sinkVec_sinkWire_47_valid = sinkVec_queue_47_deq_valid;
  assign sinkVec_sinkWire_47_bits_vd = sinkVec_queue_47_deq_bits_vd;
  assign sinkVec_sinkWire_47_bits_offset = sinkVec_queue_47_deq_bits_offset;
  assign sinkVec_sinkWire_47_bits_mask = sinkVec_queue_47_deq_bits_mask;
  assign sinkVec_sinkWire_47_bits_data = sinkVec_queue_47_deq_bits_data;
  assign sinkVec_sinkWire_47_bits_last = sinkVec_queue_47_deq_bits_last;
  assign sinkVec_sinkWire_47_bits_instructionIndex = sinkVec_queue_47_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_47_enq_bits_data;
  wire         sinkVec_queue_47_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_23 = {sinkVec_queue_47_enq_bits_data, sinkVec_queue_47_enq_bits_last};
  wire [2:0]   sinkVec_queue_47_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_47 = {sinkVec_queue_dataIn_lo_hi_23, sinkVec_queue_47_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_47_enq_bits_vd;
  wire [1:0]   sinkVec_queue_47_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_23 = {sinkVec_queue_47_enq_bits_vd, sinkVec_queue_47_enq_bits_offset};
  wire [3:0]   sinkVec_queue_47_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_47 = {sinkVec_queue_dataIn_hi_hi_23, sinkVec_queue_47_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_47 = {sinkVec_queue_dataIn_hi_47, sinkVec_queue_dataIn_lo_47};
  wire [2:0]   sinkVec_queue_dataOut_47_instructionIndex = _sinkVec_queue_fifo_47_data_out[2:0];
  wire         sinkVec_queue_dataOut_47_last = _sinkVec_queue_fifo_47_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_47_data = _sinkVec_queue_fifo_47_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_47_mask = _sinkVec_queue_fifo_47_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_47_offset = _sinkVec_queue_fifo_47_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_47_vd = _sinkVec_queue_fifo_47_data_out[46:42];
  wire         sinkVec_queue_47_enq_ready = ~_sinkVec_queue_fifo_47_full;
  wire         sinkVec_queue_47_enq_valid;
  assign sinkVec_queue_47_deq_valid = ~_sinkVec_queue_fifo_47_empty | sinkVec_queue_47_enq_valid;
  assign sinkVec_queue_47_deq_bits_vd = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_vd : sinkVec_queue_dataOut_47_vd;
  assign sinkVec_queue_47_deq_bits_offset = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_offset : sinkVec_queue_dataOut_47_offset;
  assign sinkVec_queue_47_deq_bits_mask = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_mask : sinkVec_queue_dataOut_47_mask;
  assign sinkVec_queue_47_deq_bits_data = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_data : sinkVec_queue_dataOut_47_data;
  assign sinkVec_queue_47_deq_bits_last = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_last : sinkVec_queue_dataOut_47_last;
  assign sinkVec_queue_47_deq_bits_instructionIndex = _sinkVec_queue_fifo_47_empty ? sinkVec_queue_47_enq_bits_instructionIndex : sinkVec_queue_dataOut_47_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_47;
  wire         sinkVec_releasePipe_pipe_out_47_valid = sinkVec_releasePipe_pipe_v_47;
  wire         x22_11_1_ready;
  wire         x22_11_1_valid;
  wire         sinkVec_validSource_47_valid = x22_11_1_ready & x22_11_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_47;
  wire [2:0]   sinkVec_tokenCheck_counterChange_47 = sinkVec_validSource_47_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_47 = ~(sinkVec_tokenCheck_counter_47[2]);
  assign x22_11_1_ready = sinkVec_tokenCheck_47;
  assign sinkVec_queue_47_enq_valid = sinkVec_validSink_47_valid;
  assign sinkVec_queue_47_enq_bits_vd = sinkVec_validSink_47_bits_vd;
  assign sinkVec_queue_47_enq_bits_offset = sinkVec_validSink_47_bits_offset;
  assign sinkVec_queue_47_enq_bits_mask = sinkVec_validSink_47_bits_mask;
  assign sinkVec_queue_47_enq_bits_data = sinkVec_validSink_47_bits_data;
  assign sinkVec_queue_47_enq_bits_last = sinkVec_validSink_47_bits_last;
  assign sinkVec_queue_47_enq_bits_instructionIndex = sinkVec_validSink_47_bits_instructionIndex;
  reg          sinkVec_shifterReg_47_0_valid;
  assign sinkVec_validSink_47_valid = sinkVec_shifterReg_47_0_valid;
  reg  [4:0]   sinkVec_shifterReg_47_0_bits_vd;
  assign sinkVec_validSink_47_bits_vd = sinkVec_shifterReg_47_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_47_0_bits_offset;
  assign sinkVec_validSink_47_bits_offset = sinkVec_shifterReg_47_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_47_0_bits_mask;
  assign sinkVec_validSink_47_bits_mask = sinkVec_shifterReg_47_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_47_0_bits_data;
  assign sinkVec_validSink_47_bits_data = sinkVec_shifterReg_47_0_bits_data;
  reg          sinkVec_shifterReg_47_0_bits_last;
  assign sinkVec_validSink_47_bits_last = sinkVec_shifterReg_47_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_47_0_bits_instructionIndex;
  assign sinkVec_validSink_47_bits_instructionIndex = sinkVec_shifterReg_47_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_47 = sinkVec_shifterReg_47_0_valid | sinkVec_validSource_47_valid;
  assign sinkVec_sinkWire_46_ready = sinkVec_23_0_ready;
  assign sinkVec_sinkWire_47_ready = sinkVec_23_1_ready;
  reg          maskUnitFirst_23;
  wire         tryToRead_23 = sinkVec_23_0_valid | sinkVec_23_1_valid;
  wire         sinkWire_23_valid = maskUnitFirst_23 ? sinkVec_23_0_valid : sinkVec_23_1_valid;
  wire [4:0]   sinkWire_23_bits_vd = maskUnitFirst_23 ? sinkVec_23_0_bits_vd : sinkVec_23_1_bits_vd;
  wire [1:0]   sinkWire_23_bits_offset = maskUnitFirst_23 ? sinkVec_23_0_bits_offset : sinkVec_23_1_bits_offset;
  wire [3:0]   sinkWire_23_bits_mask = maskUnitFirst_23 ? sinkVec_23_0_bits_mask : sinkVec_23_1_bits_mask;
  wire [31:0]  sinkWire_23_bits_data = maskUnitFirst_23 ? sinkVec_23_0_bits_data : sinkVec_23_1_bits_data;
  wire         sinkWire_23_bits_last = maskUnitFirst_23 ? sinkVec_23_0_bits_last : sinkVec_23_1_bits_last;
  wire [2:0]   sinkWire_23_bits_instructionIndex = maskUnitFirst_23 ? sinkVec_23_0_bits_instructionIndex : sinkVec_23_1_bits_instructionIndex;
  wire         sinkWire_23_ready;
  assign sinkVec_23_1_ready = sinkWire_23_ready & ~maskUnitFirst_23;
  assign sinkVec_23_0_ready = sinkWire_23_ready & maskUnitFirst_23;
  reg          view__writeRelease_11_pipe_v;
  wire         view__writeRelease_11_pipe_out_valid = view__writeRelease_11_pipe_v;
  reg          pipe_v_33;
  wire         pipe_out_22_valid = pipe_v_33;
  wire         _probeWire_writeQueueEnqVec_11_valid_T = x22_11_0_ready & _maskUnit_exeResp_11_valid;
  reg          instructionFinishedPipe_pipe_v_11;
  wire         instructionFinishedPipe_pipe_out_11_valid = instructionFinishedPipe_pipe_v_11;
  reg  [7:0]   instructionFinishedPipe_pipe_b_11;
  wire [7:0]   instructionFinishedPipe_pipe_out_11_bits = instructionFinishedPipe_pipe_b_11;
  wire         instructionFinished_11_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_11_bits);
  wire         instructionFinished_11_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_11_bits);
  wire         instructionFinished_11_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_11_bits);
  wire         instructionFinished_11_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_11_bits);
  assign vxsatReportVec_11 = _laneVec_11_vxsatReport[3:0];
  reg          pipe_v_34;
  reg  [31:0]  pipe_b_34;
  reg          pipe_pipe_v_11;
  wire         pipe_pipe_out_11_valid = pipe_pipe_v_11;
  reg  [31:0]  pipe_pipe_b_11;
  wire [31:0]  pipe_pipe_out_11_bits = pipe_pipe_b_11;
  reg          view__laneMaskSelect_11_pipe_v;
  reg  [5:0]   view__laneMaskSelect_11_pipe_b;
  reg          view__laneMaskSelect_11_pipe_pipe_v;
  wire         view__laneMaskSelect_11_pipe_pipe_out_valid = view__laneMaskSelect_11_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_11_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_11_pipe_pipe_out_bits = view__laneMaskSelect_11_pipe_pipe_b;
  reg          view__laneMaskSewSelect_11_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_11_pipe_b;
  reg          view__laneMaskSewSelect_11_pipe_pipe_v;
  wire         view__laneMaskSewSelect_11_pipe_pipe_out_valid = view__laneMaskSewSelect_11_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_11_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_11_pipe_pipe_out_bits = view__laneMaskSewSelect_11_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_11;
  wire         lsuLastPipe_pipe_out_11_valid = lsuLastPipe_pipe_v_11;
  reg  [7:0]   lsuLastPipe_pipe_b_11;
  wire [7:0]   lsuLastPipe_pipe_out_11_bits = lsuLastPipe_pipe_b_11;
  reg          maskLastPipe_pipe_v_11;
  wire         maskLastPipe_pipe_out_11_valid = maskLastPipe_pipe_v_11;
  reg  [7:0]   maskLastPipe_pipe_b_11;
  wire [7:0]   maskLastPipe_pipe_out_11_bits = maskLastPipe_pipe_b_11;
  wire [5:0]   writeCounter_11 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h2C};
  reg          pipe_v_35;
  wire         pipe_out_23_valid = pipe_v_35;
  reg  [5:0]   pipe_b_35;
  wire [5:0]   pipe_out_23_bits = pipe_b_35;
  assign laneRequestSinkWire_12_ready = ~laneRequestSinkWire_12_bits_issueInst | _laneVec_12_laneRequest_ready;
  wire         sinkVec_tokenCheck_48;
  wire [4:0]   sinkVec_validSource_48_bits_vs = x13_12_0_bits_vs;
  wire [1:0]   sinkVec_validSource_48_bits_offset = x13_12_0_bits_offset;
  wire [2:0]   sinkVec_validSource_48_bits_instructionIndex = x13_12_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_49;
  wire [4:0]   sinkVec_validSource_49_bits_vs = x13_12_1_bits_vs;
  wire [1:0]   sinkVec_validSource_49_bits_offset = x13_12_1_bits_offset;
  wire [2:0]   sinkVec_validSource_49_bits_instructionIndex = x13_12_1_bits_instructionIndex;
  wire         sinkVec_24_0_ready;
  wire         sinkVec_queue_48_deq_ready = sinkVec_sinkWire_48_ready;
  wire         sinkVec_queue_48_deq_valid;
  wire [4:0]   sinkVec_queue_48_deq_bits_vs;
  wire         sinkVec_24_0_valid = sinkVec_sinkWire_48_valid;
  wire [1:0]   sinkVec_queue_48_deq_bits_readSource;
  wire [4:0]   sinkVec_24_0_bits_vs = sinkVec_sinkWire_48_bits_vs;
  wire [1:0]   sinkVec_queue_48_deq_bits_offset;
  wire [1:0]   sinkVec_24_0_bits_readSource = sinkVec_sinkWire_48_bits_readSource;
  wire [2:0]   sinkVec_queue_48_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_24_0_bits_offset = sinkVec_sinkWire_48_bits_offset;
  wire [2:0]   sinkVec_24_0_bits_instructionIndex = sinkVec_sinkWire_48_bits_instructionIndex;
  wire         sinkVec_validSink_48_valid;
  wire [4:0]   sinkVec_validSink_48_bits_vs;
  wire [1:0]   sinkVec_validSink_48_bits_readSource;
  wire [1:0]   sinkVec_validSink_48_bits_offset;
  wire [2:0]   sinkVec_validSink_48_bits_instructionIndex;
  assign sinkVec_sinkWire_48_valid = sinkVec_queue_48_deq_valid;
  assign sinkVec_sinkWire_48_bits_vs = sinkVec_queue_48_deq_bits_vs;
  assign sinkVec_sinkWire_48_bits_readSource = sinkVec_queue_48_deq_bits_readSource;
  assign sinkVec_sinkWire_48_bits_offset = sinkVec_queue_48_deq_bits_offset;
  assign sinkVec_sinkWire_48_bits_instructionIndex = sinkVec_queue_48_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_48_enq_bits_offset;
  wire [2:0]   sinkVec_queue_48_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_48 = {sinkVec_queue_48_enq_bits_offset, sinkVec_queue_48_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_48_enq_bits_vs;
  wire [1:0]   sinkVec_queue_48_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_48 = {sinkVec_queue_48_enq_bits_vs, sinkVec_queue_48_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_48 = {sinkVec_queue_dataIn_hi_48, sinkVec_queue_dataIn_lo_48};
  wire [2:0]   sinkVec_queue_dataOut_48_instructionIndex = _sinkVec_queue_fifo_48_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_48_offset = _sinkVec_queue_fifo_48_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_48_readSource = _sinkVec_queue_fifo_48_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_48_vs = _sinkVec_queue_fifo_48_data_out[11:7];
  wire         sinkVec_queue_48_enq_ready = ~_sinkVec_queue_fifo_48_full;
  wire         sinkVec_queue_48_enq_valid;
  assign sinkVec_queue_48_deq_valid = ~_sinkVec_queue_fifo_48_empty | sinkVec_queue_48_enq_valid;
  assign sinkVec_queue_48_deq_bits_vs = _sinkVec_queue_fifo_48_empty ? sinkVec_queue_48_enq_bits_vs : sinkVec_queue_dataOut_48_vs;
  assign sinkVec_queue_48_deq_bits_readSource = _sinkVec_queue_fifo_48_empty ? sinkVec_queue_48_enq_bits_readSource : sinkVec_queue_dataOut_48_readSource;
  assign sinkVec_queue_48_deq_bits_offset = _sinkVec_queue_fifo_48_empty ? sinkVec_queue_48_enq_bits_offset : sinkVec_queue_dataOut_48_offset;
  assign sinkVec_queue_48_deq_bits_instructionIndex = _sinkVec_queue_fifo_48_empty ? sinkVec_queue_48_enq_bits_instructionIndex : sinkVec_queue_dataOut_48_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_48;
  wire         sinkVec_releasePipe_pipe_out_48_valid = sinkVec_releasePipe_pipe_v_48;
  wire         x13_12_0_ready;
  wire         x13_12_0_valid;
  wire         sinkVec_validSource_48_valid = x13_12_0_ready & x13_12_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_48;
  wire [2:0]   sinkVec_tokenCheck_counterChange_48 = sinkVec_validSource_48_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_48 = ~(sinkVec_tokenCheck_counter_48[2]);
  assign x13_12_0_ready = sinkVec_tokenCheck_48;
  assign sinkVec_queue_48_enq_valid = sinkVec_validSink_48_valid;
  assign sinkVec_queue_48_enq_bits_vs = sinkVec_validSink_48_bits_vs;
  assign sinkVec_queue_48_enq_bits_readSource = sinkVec_validSink_48_bits_readSource;
  assign sinkVec_queue_48_enq_bits_offset = sinkVec_validSink_48_bits_offset;
  assign sinkVec_queue_48_enq_bits_instructionIndex = sinkVec_validSink_48_bits_instructionIndex;
  reg          sinkVec_shifterReg_48_0_valid;
  assign sinkVec_validSink_48_valid = sinkVec_shifterReg_48_0_valid;
  reg  [4:0]   sinkVec_shifterReg_48_0_bits_vs;
  assign sinkVec_validSink_48_bits_vs = sinkVec_shifterReg_48_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_48_0_bits_readSource;
  assign sinkVec_validSink_48_bits_readSource = sinkVec_shifterReg_48_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_48_0_bits_offset;
  assign sinkVec_validSink_48_bits_offset = sinkVec_shifterReg_48_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_48_0_bits_instructionIndex;
  assign sinkVec_validSink_48_bits_instructionIndex = sinkVec_shifterReg_48_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_48 = sinkVec_shifterReg_48_0_valid | sinkVec_validSource_48_valid;
  wire         sinkVec_24_1_ready;
  wire         sinkVec_queue_49_deq_ready = sinkVec_sinkWire_49_ready;
  wire         sinkVec_queue_49_deq_valid;
  wire [4:0]   sinkVec_queue_49_deq_bits_vs;
  wire         sinkVec_24_1_valid = sinkVec_sinkWire_49_valid;
  wire [1:0]   sinkVec_queue_49_deq_bits_readSource;
  wire [4:0]   sinkVec_24_1_bits_vs = sinkVec_sinkWire_49_bits_vs;
  wire [1:0]   sinkVec_queue_49_deq_bits_offset;
  wire [1:0]   sinkVec_24_1_bits_readSource = sinkVec_sinkWire_49_bits_readSource;
  wire [2:0]   sinkVec_queue_49_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_24_1_bits_offset = sinkVec_sinkWire_49_bits_offset;
  wire [2:0]   sinkVec_24_1_bits_instructionIndex = sinkVec_sinkWire_49_bits_instructionIndex;
  wire         sinkVec_validSink_49_valid;
  wire [4:0]   sinkVec_validSink_49_bits_vs;
  wire [1:0]   sinkVec_validSink_49_bits_readSource;
  wire [1:0]   sinkVec_validSink_49_bits_offset;
  wire [2:0]   sinkVec_validSink_49_bits_instructionIndex;
  assign sinkVec_sinkWire_49_valid = sinkVec_queue_49_deq_valid;
  assign sinkVec_sinkWire_49_bits_vs = sinkVec_queue_49_deq_bits_vs;
  assign sinkVec_sinkWire_49_bits_readSource = sinkVec_queue_49_deq_bits_readSource;
  assign sinkVec_sinkWire_49_bits_offset = sinkVec_queue_49_deq_bits_offset;
  assign sinkVec_sinkWire_49_bits_instructionIndex = sinkVec_queue_49_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_49_enq_bits_offset;
  wire [2:0]   sinkVec_queue_49_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_49 = {sinkVec_queue_49_enq_bits_offset, sinkVec_queue_49_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_49_enq_bits_vs;
  wire [1:0]   sinkVec_queue_49_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_49 = {sinkVec_queue_49_enq_bits_vs, sinkVec_queue_49_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_49 = {sinkVec_queue_dataIn_hi_49, sinkVec_queue_dataIn_lo_49};
  wire [2:0]   sinkVec_queue_dataOut_49_instructionIndex = _sinkVec_queue_fifo_49_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_49_offset = _sinkVec_queue_fifo_49_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_49_readSource = _sinkVec_queue_fifo_49_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_49_vs = _sinkVec_queue_fifo_49_data_out[11:7];
  wire         sinkVec_queue_49_enq_ready = ~_sinkVec_queue_fifo_49_full;
  wire         sinkVec_queue_49_enq_valid;
  assign sinkVec_queue_49_deq_valid = ~_sinkVec_queue_fifo_49_empty | sinkVec_queue_49_enq_valid;
  assign sinkVec_queue_49_deq_bits_vs = _sinkVec_queue_fifo_49_empty ? sinkVec_queue_49_enq_bits_vs : sinkVec_queue_dataOut_49_vs;
  assign sinkVec_queue_49_deq_bits_readSource = _sinkVec_queue_fifo_49_empty ? sinkVec_queue_49_enq_bits_readSource : sinkVec_queue_dataOut_49_readSource;
  assign sinkVec_queue_49_deq_bits_offset = _sinkVec_queue_fifo_49_empty ? sinkVec_queue_49_enq_bits_offset : sinkVec_queue_dataOut_49_offset;
  assign sinkVec_queue_49_deq_bits_instructionIndex = _sinkVec_queue_fifo_49_empty ? sinkVec_queue_49_enq_bits_instructionIndex : sinkVec_queue_dataOut_49_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_49;
  wire         sinkVec_releasePipe_pipe_out_49_valid = sinkVec_releasePipe_pipe_v_49;
  wire         x13_12_1_ready;
  wire         x13_12_1_valid;
  wire         sinkVec_validSource_49_valid = x13_12_1_ready & x13_12_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_49;
  wire [2:0]   sinkVec_tokenCheck_counterChange_49 = sinkVec_validSource_49_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_49 = ~(sinkVec_tokenCheck_counter_49[2]);
  assign x13_12_1_ready = sinkVec_tokenCheck_49;
  assign sinkVec_queue_49_enq_valid = sinkVec_validSink_49_valid;
  assign sinkVec_queue_49_enq_bits_vs = sinkVec_validSink_49_bits_vs;
  assign sinkVec_queue_49_enq_bits_readSource = sinkVec_validSink_49_bits_readSource;
  assign sinkVec_queue_49_enq_bits_offset = sinkVec_validSink_49_bits_offset;
  assign sinkVec_queue_49_enq_bits_instructionIndex = sinkVec_validSink_49_bits_instructionIndex;
  reg          sinkVec_shifterReg_49_0_valid;
  assign sinkVec_validSink_49_valid = sinkVec_shifterReg_49_0_valid;
  reg  [4:0]   sinkVec_shifterReg_49_0_bits_vs;
  assign sinkVec_validSink_49_bits_vs = sinkVec_shifterReg_49_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_49_0_bits_readSource;
  assign sinkVec_validSink_49_bits_readSource = sinkVec_shifterReg_49_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_49_0_bits_offset;
  assign sinkVec_validSink_49_bits_offset = sinkVec_shifterReg_49_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_49_0_bits_instructionIndex;
  assign sinkVec_validSink_49_bits_instructionIndex = sinkVec_shifterReg_49_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_49 = sinkVec_shifterReg_49_0_valid | sinkVec_validSource_49_valid;
  assign sinkVec_sinkWire_48_ready = sinkVec_24_0_ready;
  assign sinkVec_sinkWire_49_ready = sinkVec_24_1_ready;
  reg          maskUnitFirst_24;
  wire         tryToRead_24 = sinkVec_24_0_valid | sinkVec_24_1_valid;
  wire         sinkWire_24_valid = maskUnitFirst_24 ? sinkVec_24_0_valid : sinkVec_24_1_valid;
  wire [4:0]   sinkWire_24_bits_vs = maskUnitFirst_24 ? sinkVec_24_0_bits_vs : sinkVec_24_1_bits_vs;
  wire [1:0]   sinkWire_24_bits_readSource = maskUnitFirst_24 ? sinkVec_24_0_bits_readSource : sinkVec_24_1_bits_readSource;
  wire [1:0]   sinkWire_24_bits_offset = maskUnitFirst_24 ? sinkVec_24_0_bits_offset : sinkVec_24_1_bits_offset;
  wire [2:0]   sinkWire_24_bits_instructionIndex = maskUnitFirst_24 ? sinkVec_24_0_bits_instructionIndex : sinkVec_24_1_bits_instructionIndex;
  wire         sinkWire_24_ready;
  assign sinkVec_24_1_ready = sinkWire_24_ready & ~maskUnitFirst_24;
  assign sinkVec_24_0_ready = sinkWire_24_ready & maskUnitFirst_24;
  reg          accessDataValid_pipe_v_24;
  reg          accessDataValid_pipe_pipe_v_24;
  wire         accessDataValid_pipe_pipe_out_24_valid = accessDataValid_pipe_pipe_v_24;
  wire         accessDataSource_24_valid = accessDataValid_pipe_pipe_out_24_valid;
  reg          shifterReg_40_0_valid;
  reg  [31:0]  shifterReg_40_0_bits;
  wire         shifterValid_40 = shifterReg_40_0_valid | accessDataSource_24_valid;
  reg          accessDataValid_pipe_v_25;
  reg          accessDataValid_pipe_pipe_v_25;
  wire         accessDataValid_pipe_pipe_out_25_valid = accessDataValid_pipe_pipe_v_25;
  wire         accessDataSource_25_valid = accessDataValid_pipe_pipe_out_25_valid;
  reg          shifterReg_41_0_valid;
  reg  [31:0]  shifterReg_41_0_bits;
  wire         shifterValid_41 = shifterReg_41_0_valid | accessDataSource_25_valid;
  wire         sinkVec_tokenCheck_50;
  wire [4:0]   sinkVec_validSource_50_bits_vd = x22_12_0_bits_vd;
  wire [1:0]   sinkVec_validSource_50_bits_offset = x22_12_0_bits_offset;
  wire [3:0]   sinkVec_validSource_50_bits_mask = x22_12_0_bits_mask;
  wire [31:0]  sinkVec_validSource_50_bits_data = x22_12_0_bits_data;
  wire [2:0]   sinkVec_validSource_50_bits_instructionIndex = x22_12_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_51;
  wire [4:0]   sinkVec_validSource_51_bits_vd = x22_12_1_bits_vd;
  wire [1:0]   sinkVec_validSource_51_bits_offset = x22_12_1_bits_offset;
  wire [3:0]   sinkVec_validSource_51_bits_mask = x22_12_1_bits_mask;
  wire [31:0]  sinkVec_validSource_51_bits_data = x22_12_1_bits_data;
  wire         sinkVec_validSource_51_bits_last = x22_12_1_bits_last;
  wire [2:0]   sinkVec_validSource_51_bits_instructionIndex = x22_12_1_bits_instructionIndex;
  wire         sinkVec_25_0_ready;
  wire         sinkVec_queue_50_deq_ready = sinkVec_sinkWire_50_ready;
  wire         sinkVec_queue_50_deq_valid;
  wire [4:0]   sinkVec_queue_50_deq_bits_vd;
  wire         sinkVec_25_0_valid = sinkVec_sinkWire_50_valid;
  wire [1:0]   sinkVec_queue_50_deq_bits_offset;
  wire [4:0]   sinkVec_25_0_bits_vd = sinkVec_sinkWire_50_bits_vd;
  wire [3:0]   sinkVec_queue_50_deq_bits_mask;
  wire [1:0]   sinkVec_25_0_bits_offset = sinkVec_sinkWire_50_bits_offset;
  wire [31:0]  sinkVec_queue_50_deq_bits_data;
  wire [3:0]   sinkVec_25_0_bits_mask = sinkVec_sinkWire_50_bits_mask;
  wire         sinkVec_queue_50_deq_bits_last;
  wire [31:0]  sinkVec_25_0_bits_data = sinkVec_sinkWire_50_bits_data;
  wire [2:0]   sinkVec_queue_50_deq_bits_instructionIndex;
  wire         sinkVec_25_0_bits_last = sinkVec_sinkWire_50_bits_last;
  wire [2:0]   sinkVec_25_0_bits_instructionIndex = sinkVec_sinkWire_50_bits_instructionIndex;
  wire         sinkVec_validSink_50_valid;
  wire [4:0]   sinkVec_validSink_50_bits_vd;
  wire [1:0]   sinkVec_validSink_50_bits_offset;
  wire [3:0]   sinkVec_validSink_50_bits_mask;
  wire [31:0]  sinkVec_validSink_50_bits_data;
  wire [2:0]   sinkVec_validSink_50_bits_instructionIndex;
  assign sinkVec_sinkWire_50_valid = sinkVec_queue_50_deq_valid;
  assign sinkVec_sinkWire_50_bits_vd = sinkVec_queue_50_deq_bits_vd;
  assign sinkVec_sinkWire_50_bits_offset = sinkVec_queue_50_deq_bits_offset;
  assign sinkVec_sinkWire_50_bits_mask = sinkVec_queue_50_deq_bits_mask;
  assign sinkVec_sinkWire_50_bits_data = sinkVec_queue_50_deq_bits_data;
  assign sinkVec_sinkWire_50_bits_last = sinkVec_queue_50_deq_bits_last;
  assign sinkVec_sinkWire_50_bits_instructionIndex = sinkVec_queue_50_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_50_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_24 = {sinkVec_queue_50_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_50_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_50 = {sinkVec_queue_dataIn_lo_hi_24, sinkVec_queue_50_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_50_enq_bits_vd;
  wire [1:0]   sinkVec_queue_50_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_24 = {sinkVec_queue_50_enq_bits_vd, sinkVec_queue_50_enq_bits_offset};
  wire [3:0]   sinkVec_queue_50_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_50 = {sinkVec_queue_dataIn_hi_hi_24, sinkVec_queue_50_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_50 = {sinkVec_queue_dataIn_hi_50, sinkVec_queue_dataIn_lo_50};
  wire [2:0]   sinkVec_queue_dataOut_50_instructionIndex = _sinkVec_queue_fifo_50_data_out[2:0];
  wire         sinkVec_queue_dataOut_50_last = _sinkVec_queue_fifo_50_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_50_data = _sinkVec_queue_fifo_50_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_50_mask = _sinkVec_queue_fifo_50_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_50_offset = _sinkVec_queue_fifo_50_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_50_vd = _sinkVec_queue_fifo_50_data_out[46:42];
  wire         sinkVec_queue_50_enq_ready = ~_sinkVec_queue_fifo_50_full;
  wire         sinkVec_queue_50_enq_valid;
  assign sinkVec_queue_50_deq_valid = ~_sinkVec_queue_fifo_50_empty | sinkVec_queue_50_enq_valid;
  assign sinkVec_queue_50_deq_bits_vd = _sinkVec_queue_fifo_50_empty ? sinkVec_queue_50_enq_bits_vd : sinkVec_queue_dataOut_50_vd;
  assign sinkVec_queue_50_deq_bits_offset = _sinkVec_queue_fifo_50_empty ? sinkVec_queue_50_enq_bits_offset : sinkVec_queue_dataOut_50_offset;
  assign sinkVec_queue_50_deq_bits_mask = _sinkVec_queue_fifo_50_empty ? sinkVec_queue_50_enq_bits_mask : sinkVec_queue_dataOut_50_mask;
  assign sinkVec_queue_50_deq_bits_data = _sinkVec_queue_fifo_50_empty ? sinkVec_queue_50_enq_bits_data : sinkVec_queue_dataOut_50_data;
  assign sinkVec_queue_50_deq_bits_last = ~_sinkVec_queue_fifo_50_empty & sinkVec_queue_dataOut_50_last;
  assign sinkVec_queue_50_deq_bits_instructionIndex = _sinkVec_queue_fifo_50_empty ? sinkVec_queue_50_enq_bits_instructionIndex : sinkVec_queue_dataOut_50_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_50;
  wire         sinkVec_releasePipe_pipe_out_50_valid = sinkVec_releasePipe_pipe_v_50;
  wire         x22_12_0_ready;
  wire         x22_12_0_valid;
  wire         sinkVec_validSource_50_valid = x22_12_0_ready & x22_12_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_50;
  wire [2:0]   sinkVec_tokenCheck_counterChange_50 = sinkVec_validSource_50_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_50 = ~(sinkVec_tokenCheck_counter_50[2]);
  assign x22_12_0_ready = sinkVec_tokenCheck_50;
  assign sinkVec_queue_50_enq_valid = sinkVec_validSink_50_valid;
  assign sinkVec_queue_50_enq_bits_vd = sinkVec_validSink_50_bits_vd;
  assign sinkVec_queue_50_enq_bits_offset = sinkVec_validSink_50_bits_offset;
  assign sinkVec_queue_50_enq_bits_mask = sinkVec_validSink_50_bits_mask;
  assign sinkVec_queue_50_enq_bits_data = sinkVec_validSink_50_bits_data;
  assign sinkVec_queue_50_enq_bits_instructionIndex = sinkVec_validSink_50_bits_instructionIndex;
  reg          sinkVec_shifterReg_50_0_valid;
  assign sinkVec_validSink_50_valid = sinkVec_shifterReg_50_0_valid;
  reg  [4:0]   sinkVec_shifterReg_50_0_bits_vd;
  assign sinkVec_validSink_50_bits_vd = sinkVec_shifterReg_50_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_50_0_bits_offset;
  assign sinkVec_validSink_50_bits_offset = sinkVec_shifterReg_50_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_50_0_bits_mask;
  assign sinkVec_validSink_50_bits_mask = sinkVec_shifterReg_50_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_50_0_bits_data;
  assign sinkVec_validSink_50_bits_data = sinkVec_shifterReg_50_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_50_0_bits_instructionIndex;
  assign sinkVec_validSink_50_bits_instructionIndex = sinkVec_shifterReg_50_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_50 = sinkVec_shifterReg_50_0_valid | sinkVec_validSource_50_valid;
  wire         sinkVec_25_1_ready;
  wire         sinkVec_queue_51_deq_ready = sinkVec_sinkWire_51_ready;
  wire         sinkVec_queue_51_deq_valid;
  wire [4:0]   sinkVec_queue_51_deq_bits_vd;
  wire         sinkVec_25_1_valid = sinkVec_sinkWire_51_valid;
  wire [1:0]   sinkVec_queue_51_deq_bits_offset;
  wire [4:0]   sinkVec_25_1_bits_vd = sinkVec_sinkWire_51_bits_vd;
  wire [3:0]   sinkVec_queue_51_deq_bits_mask;
  wire [1:0]   sinkVec_25_1_bits_offset = sinkVec_sinkWire_51_bits_offset;
  wire [31:0]  sinkVec_queue_51_deq_bits_data;
  wire [3:0]   sinkVec_25_1_bits_mask = sinkVec_sinkWire_51_bits_mask;
  wire         sinkVec_queue_51_deq_bits_last;
  wire [31:0]  sinkVec_25_1_bits_data = sinkVec_sinkWire_51_bits_data;
  wire [2:0]   sinkVec_queue_51_deq_bits_instructionIndex;
  wire         sinkVec_25_1_bits_last = sinkVec_sinkWire_51_bits_last;
  wire [2:0]   sinkVec_25_1_bits_instructionIndex = sinkVec_sinkWire_51_bits_instructionIndex;
  wire         sinkVec_validSink_51_valid;
  wire [4:0]   sinkVec_validSink_51_bits_vd;
  wire [1:0]   sinkVec_validSink_51_bits_offset;
  wire [3:0]   sinkVec_validSink_51_bits_mask;
  wire [31:0]  sinkVec_validSink_51_bits_data;
  wire         sinkVec_validSink_51_bits_last;
  wire [2:0]   sinkVec_validSink_51_bits_instructionIndex;
  assign sinkVec_sinkWire_51_valid = sinkVec_queue_51_deq_valid;
  assign sinkVec_sinkWire_51_bits_vd = sinkVec_queue_51_deq_bits_vd;
  assign sinkVec_sinkWire_51_bits_offset = sinkVec_queue_51_deq_bits_offset;
  assign sinkVec_sinkWire_51_bits_mask = sinkVec_queue_51_deq_bits_mask;
  assign sinkVec_sinkWire_51_bits_data = sinkVec_queue_51_deq_bits_data;
  assign sinkVec_sinkWire_51_bits_last = sinkVec_queue_51_deq_bits_last;
  assign sinkVec_sinkWire_51_bits_instructionIndex = sinkVec_queue_51_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_51_enq_bits_data;
  wire         sinkVec_queue_51_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_25 = {sinkVec_queue_51_enq_bits_data, sinkVec_queue_51_enq_bits_last};
  wire [2:0]   sinkVec_queue_51_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_51 = {sinkVec_queue_dataIn_lo_hi_25, sinkVec_queue_51_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_51_enq_bits_vd;
  wire [1:0]   sinkVec_queue_51_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_25 = {sinkVec_queue_51_enq_bits_vd, sinkVec_queue_51_enq_bits_offset};
  wire [3:0]   sinkVec_queue_51_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_51 = {sinkVec_queue_dataIn_hi_hi_25, sinkVec_queue_51_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_51 = {sinkVec_queue_dataIn_hi_51, sinkVec_queue_dataIn_lo_51};
  wire [2:0]   sinkVec_queue_dataOut_51_instructionIndex = _sinkVec_queue_fifo_51_data_out[2:0];
  wire         sinkVec_queue_dataOut_51_last = _sinkVec_queue_fifo_51_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_51_data = _sinkVec_queue_fifo_51_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_51_mask = _sinkVec_queue_fifo_51_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_51_offset = _sinkVec_queue_fifo_51_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_51_vd = _sinkVec_queue_fifo_51_data_out[46:42];
  wire         sinkVec_queue_51_enq_ready = ~_sinkVec_queue_fifo_51_full;
  wire         sinkVec_queue_51_enq_valid;
  assign sinkVec_queue_51_deq_valid = ~_sinkVec_queue_fifo_51_empty | sinkVec_queue_51_enq_valid;
  assign sinkVec_queue_51_deq_bits_vd = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_vd : sinkVec_queue_dataOut_51_vd;
  assign sinkVec_queue_51_deq_bits_offset = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_offset : sinkVec_queue_dataOut_51_offset;
  assign sinkVec_queue_51_deq_bits_mask = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_mask : sinkVec_queue_dataOut_51_mask;
  assign sinkVec_queue_51_deq_bits_data = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_data : sinkVec_queue_dataOut_51_data;
  assign sinkVec_queue_51_deq_bits_last = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_last : sinkVec_queue_dataOut_51_last;
  assign sinkVec_queue_51_deq_bits_instructionIndex = _sinkVec_queue_fifo_51_empty ? sinkVec_queue_51_enq_bits_instructionIndex : sinkVec_queue_dataOut_51_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_51;
  wire         sinkVec_releasePipe_pipe_out_51_valid = sinkVec_releasePipe_pipe_v_51;
  wire         x22_12_1_ready;
  wire         x22_12_1_valid;
  wire         sinkVec_validSource_51_valid = x22_12_1_ready & x22_12_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_51;
  wire [2:0]   sinkVec_tokenCheck_counterChange_51 = sinkVec_validSource_51_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_51 = ~(sinkVec_tokenCheck_counter_51[2]);
  assign x22_12_1_ready = sinkVec_tokenCheck_51;
  assign sinkVec_queue_51_enq_valid = sinkVec_validSink_51_valid;
  assign sinkVec_queue_51_enq_bits_vd = sinkVec_validSink_51_bits_vd;
  assign sinkVec_queue_51_enq_bits_offset = sinkVec_validSink_51_bits_offset;
  assign sinkVec_queue_51_enq_bits_mask = sinkVec_validSink_51_bits_mask;
  assign sinkVec_queue_51_enq_bits_data = sinkVec_validSink_51_bits_data;
  assign sinkVec_queue_51_enq_bits_last = sinkVec_validSink_51_bits_last;
  assign sinkVec_queue_51_enq_bits_instructionIndex = sinkVec_validSink_51_bits_instructionIndex;
  reg          sinkVec_shifterReg_51_0_valid;
  assign sinkVec_validSink_51_valid = sinkVec_shifterReg_51_0_valid;
  reg  [4:0]   sinkVec_shifterReg_51_0_bits_vd;
  assign sinkVec_validSink_51_bits_vd = sinkVec_shifterReg_51_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_51_0_bits_offset;
  assign sinkVec_validSink_51_bits_offset = sinkVec_shifterReg_51_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_51_0_bits_mask;
  assign sinkVec_validSink_51_bits_mask = sinkVec_shifterReg_51_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_51_0_bits_data;
  assign sinkVec_validSink_51_bits_data = sinkVec_shifterReg_51_0_bits_data;
  reg          sinkVec_shifterReg_51_0_bits_last;
  assign sinkVec_validSink_51_bits_last = sinkVec_shifterReg_51_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_51_0_bits_instructionIndex;
  assign sinkVec_validSink_51_bits_instructionIndex = sinkVec_shifterReg_51_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_51 = sinkVec_shifterReg_51_0_valid | sinkVec_validSource_51_valid;
  assign sinkVec_sinkWire_50_ready = sinkVec_25_0_ready;
  assign sinkVec_sinkWire_51_ready = sinkVec_25_1_ready;
  reg          maskUnitFirst_25;
  wire         tryToRead_25 = sinkVec_25_0_valid | sinkVec_25_1_valid;
  wire         sinkWire_25_valid = maskUnitFirst_25 ? sinkVec_25_0_valid : sinkVec_25_1_valid;
  wire [4:0]   sinkWire_25_bits_vd = maskUnitFirst_25 ? sinkVec_25_0_bits_vd : sinkVec_25_1_bits_vd;
  wire [1:0]   sinkWire_25_bits_offset = maskUnitFirst_25 ? sinkVec_25_0_bits_offset : sinkVec_25_1_bits_offset;
  wire [3:0]   sinkWire_25_bits_mask = maskUnitFirst_25 ? sinkVec_25_0_bits_mask : sinkVec_25_1_bits_mask;
  wire [31:0]  sinkWire_25_bits_data = maskUnitFirst_25 ? sinkVec_25_0_bits_data : sinkVec_25_1_bits_data;
  wire         sinkWire_25_bits_last = maskUnitFirst_25 ? sinkVec_25_0_bits_last : sinkVec_25_1_bits_last;
  wire [2:0]   sinkWire_25_bits_instructionIndex = maskUnitFirst_25 ? sinkVec_25_0_bits_instructionIndex : sinkVec_25_1_bits_instructionIndex;
  wire         sinkWire_25_ready;
  assign sinkVec_25_1_ready = sinkWire_25_ready & ~maskUnitFirst_25;
  assign sinkVec_25_0_ready = sinkWire_25_ready & maskUnitFirst_25;
  reg          view__writeRelease_12_pipe_v;
  wire         view__writeRelease_12_pipe_out_valid = view__writeRelease_12_pipe_v;
  reg          pipe_v_36;
  wire         pipe_out_24_valid = pipe_v_36;
  wire         _probeWire_writeQueueEnqVec_12_valid_T = x22_12_0_ready & _maskUnit_exeResp_12_valid;
  reg          instructionFinishedPipe_pipe_v_12;
  wire         instructionFinishedPipe_pipe_out_12_valid = instructionFinishedPipe_pipe_v_12;
  reg  [7:0]   instructionFinishedPipe_pipe_b_12;
  wire [7:0]   instructionFinishedPipe_pipe_out_12_bits = instructionFinishedPipe_pipe_b_12;
  wire         instructionFinished_12_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_12_bits);
  wire         instructionFinished_12_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_12_bits);
  wire         instructionFinished_12_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_12_bits);
  wire         instructionFinished_12_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_12_bits);
  assign vxsatReportVec_12 = _laneVec_12_vxsatReport[3:0];
  reg          pipe_v_37;
  reg  [31:0]  pipe_b_37;
  reg          pipe_pipe_v_12;
  wire         pipe_pipe_out_12_valid = pipe_pipe_v_12;
  reg  [31:0]  pipe_pipe_b_12;
  wire [31:0]  pipe_pipe_out_12_bits = pipe_pipe_b_12;
  reg          view__laneMaskSelect_12_pipe_v;
  reg  [5:0]   view__laneMaskSelect_12_pipe_b;
  reg          view__laneMaskSelect_12_pipe_pipe_v;
  wire         view__laneMaskSelect_12_pipe_pipe_out_valid = view__laneMaskSelect_12_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_12_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_12_pipe_pipe_out_bits = view__laneMaskSelect_12_pipe_pipe_b;
  reg          view__laneMaskSewSelect_12_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_12_pipe_b;
  reg          view__laneMaskSewSelect_12_pipe_pipe_v;
  wire         view__laneMaskSewSelect_12_pipe_pipe_out_valid = view__laneMaskSewSelect_12_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_12_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_12_pipe_pipe_out_bits = view__laneMaskSewSelect_12_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_12;
  wire         lsuLastPipe_pipe_out_12_valid = lsuLastPipe_pipe_v_12;
  reg  [7:0]   lsuLastPipe_pipe_b_12;
  wire [7:0]   lsuLastPipe_pipe_out_12_bits = lsuLastPipe_pipe_b_12;
  reg          maskLastPipe_pipe_v_12;
  wire         maskLastPipe_pipe_out_12_valid = maskLastPipe_pipe_v_12;
  reg  [7:0]   maskLastPipe_pipe_b_12;
  wire [7:0]   maskLastPipe_pipe_out_12_bits = maskLastPipe_pipe_b_12;
  wire [5:0]   writeCounter_12 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h30};
  reg          pipe_v_38;
  wire         pipe_out_25_valid = pipe_v_38;
  reg  [5:0]   pipe_b_38;
  wire [5:0]   pipe_out_25_bits = pipe_b_38;
  assign laneRequestSinkWire_13_ready = ~laneRequestSinkWire_13_bits_issueInst | _laneVec_13_laneRequest_ready;
  wire         sinkVec_tokenCheck_52;
  wire [4:0]   sinkVec_validSource_52_bits_vs = x13_13_0_bits_vs;
  wire [1:0]   sinkVec_validSource_52_bits_offset = x13_13_0_bits_offset;
  wire [2:0]   sinkVec_validSource_52_bits_instructionIndex = x13_13_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_53;
  wire [4:0]   sinkVec_validSource_53_bits_vs = x13_13_1_bits_vs;
  wire [1:0]   sinkVec_validSource_53_bits_offset = x13_13_1_bits_offset;
  wire [2:0]   sinkVec_validSource_53_bits_instructionIndex = x13_13_1_bits_instructionIndex;
  wire         sinkVec_26_0_ready;
  wire         sinkVec_queue_52_deq_ready = sinkVec_sinkWire_52_ready;
  wire         sinkVec_queue_52_deq_valid;
  wire [4:0]   sinkVec_queue_52_deq_bits_vs;
  wire         sinkVec_26_0_valid = sinkVec_sinkWire_52_valid;
  wire [1:0]   sinkVec_queue_52_deq_bits_readSource;
  wire [4:0]   sinkVec_26_0_bits_vs = sinkVec_sinkWire_52_bits_vs;
  wire [1:0]   sinkVec_queue_52_deq_bits_offset;
  wire [1:0]   sinkVec_26_0_bits_readSource = sinkVec_sinkWire_52_bits_readSource;
  wire [2:0]   sinkVec_queue_52_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_26_0_bits_offset = sinkVec_sinkWire_52_bits_offset;
  wire [2:0]   sinkVec_26_0_bits_instructionIndex = sinkVec_sinkWire_52_bits_instructionIndex;
  wire         sinkVec_validSink_52_valid;
  wire [4:0]   sinkVec_validSink_52_bits_vs;
  wire [1:0]   sinkVec_validSink_52_bits_readSource;
  wire [1:0]   sinkVec_validSink_52_bits_offset;
  wire [2:0]   sinkVec_validSink_52_bits_instructionIndex;
  assign sinkVec_sinkWire_52_valid = sinkVec_queue_52_deq_valid;
  assign sinkVec_sinkWire_52_bits_vs = sinkVec_queue_52_deq_bits_vs;
  assign sinkVec_sinkWire_52_bits_readSource = sinkVec_queue_52_deq_bits_readSource;
  assign sinkVec_sinkWire_52_bits_offset = sinkVec_queue_52_deq_bits_offset;
  assign sinkVec_sinkWire_52_bits_instructionIndex = sinkVec_queue_52_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_52_enq_bits_offset;
  wire [2:0]   sinkVec_queue_52_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_52 = {sinkVec_queue_52_enq_bits_offset, sinkVec_queue_52_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_52_enq_bits_vs;
  wire [1:0]   sinkVec_queue_52_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_52 = {sinkVec_queue_52_enq_bits_vs, sinkVec_queue_52_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_52 = {sinkVec_queue_dataIn_hi_52, sinkVec_queue_dataIn_lo_52};
  wire [2:0]   sinkVec_queue_dataOut_52_instructionIndex = _sinkVec_queue_fifo_52_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_52_offset = _sinkVec_queue_fifo_52_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_52_readSource = _sinkVec_queue_fifo_52_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_52_vs = _sinkVec_queue_fifo_52_data_out[11:7];
  wire         sinkVec_queue_52_enq_ready = ~_sinkVec_queue_fifo_52_full;
  wire         sinkVec_queue_52_enq_valid;
  assign sinkVec_queue_52_deq_valid = ~_sinkVec_queue_fifo_52_empty | sinkVec_queue_52_enq_valid;
  assign sinkVec_queue_52_deq_bits_vs = _sinkVec_queue_fifo_52_empty ? sinkVec_queue_52_enq_bits_vs : sinkVec_queue_dataOut_52_vs;
  assign sinkVec_queue_52_deq_bits_readSource = _sinkVec_queue_fifo_52_empty ? sinkVec_queue_52_enq_bits_readSource : sinkVec_queue_dataOut_52_readSource;
  assign sinkVec_queue_52_deq_bits_offset = _sinkVec_queue_fifo_52_empty ? sinkVec_queue_52_enq_bits_offset : sinkVec_queue_dataOut_52_offset;
  assign sinkVec_queue_52_deq_bits_instructionIndex = _sinkVec_queue_fifo_52_empty ? sinkVec_queue_52_enq_bits_instructionIndex : sinkVec_queue_dataOut_52_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_52;
  wire         sinkVec_releasePipe_pipe_out_52_valid = sinkVec_releasePipe_pipe_v_52;
  wire         x13_13_0_ready;
  wire         x13_13_0_valid;
  wire         sinkVec_validSource_52_valid = x13_13_0_ready & x13_13_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_52;
  wire [2:0]   sinkVec_tokenCheck_counterChange_52 = sinkVec_validSource_52_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_52 = ~(sinkVec_tokenCheck_counter_52[2]);
  assign x13_13_0_ready = sinkVec_tokenCheck_52;
  assign sinkVec_queue_52_enq_valid = sinkVec_validSink_52_valid;
  assign sinkVec_queue_52_enq_bits_vs = sinkVec_validSink_52_bits_vs;
  assign sinkVec_queue_52_enq_bits_readSource = sinkVec_validSink_52_bits_readSource;
  assign sinkVec_queue_52_enq_bits_offset = sinkVec_validSink_52_bits_offset;
  assign sinkVec_queue_52_enq_bits_instructionIndex = sinkVec_validSink_52_bits_instructionIndex;
  reg          sinkVec_shifterReg_52_0_valid;
  assign sinkVec_validSink_52_valid = sinkVec_shifterReg_52_0_valid;
  reg  [4:0]   sinkVec_shifterReg_52_0_bits_vs;
  assign sinkVec_validSink_52_bits_vs = sinkVec_shifterReg_52_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_52_0_bits_readSource;
  assign sinkVec_validSink_52_bits_readSource = sinkVec_shifterReg_52_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_52_0_bits_offset;
  assign sinkVec_validSink_52_bits_offset = sinkVec_shifterReg_52_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_52_0_bits_instructionIndex;
  assign sinkVec_validSink_52_bits_instructionIndex = sinkVec_shifterReg_52_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_52 = sinkVec_shifterReg_52_0_valid | sinkVec_validSource_52_valid;
  wire         sinkVec_26_1_ready;
  wire         sinkVec_queue_53_deq_ready = sinkVec_sinkWire_53_ready;
  wire         sinkVec_queue_53_deq_valid;
  wire [4:0]   sinkVec_queue_53_deq_bits_vs;
  wire         sinkVec_26_1_valid = sinkVec_sinkWire_53_valid;
  wire [1:0]   sinkVec_queue_53_deq_bits_readSource;
  wire [4:0]   sinkVec_26_1_bits_vs = sinkVec_sinkWire_53_bits_vs;
  wire [1:0]   sinkVec_queue_53_deq_bits_offset;
  wire [1:0]   sinkVec_26_1_bits_readSource = sinkVec_sinkWire_53_bits_readSource;
  wire [2:0]   sinkVec_queue_53_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_26_1_bits_offset = sinkVec_sinkWire_53_bits_offset;
  wire [2:0]   sinkVec_26_1_bits_instructionIndex = sinkVec_sinkWire_53_bits_instructionIndex;
  wire         sinkVec_validSink_53_valid;
  wire [4:0]   sinkVec_validSink_53_bits_vs;
  wire [1:0]   sinkVec_validSink_53_bits_readSource;
  wire [1:0]   sinkVec_validSink_53_bits_offset;
  wire [2:0]   sinkVec_validSink_53_bits_instructionIndex;
  assign sinkVec_sinkWire_53_valid = sinkVec_queue_53_deq_valid;
  assign sinkVec_sinkWire_53_bits_vs = sinkVec_queue_53_deq_bits_vs;
  assign sinkVec_sinkWire_53_bits_readSource = sinkVec_queue_53_deq_bits_readSource;
  assign sinkVec_sinkWire_53_bits_offset = sinkVec_queue_53_deq_bits_offset;
  assign sinkVec_sinkWire_53_bits_instructionIndex = sinkVec_queue_53_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_53_enq_bits_offset;
  wire [2:0]   sinkVec_queue_53_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_53 = {sinkVec_queue_53_enq_bits_offset, sinkVec_queue_53_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_53_enq_bits_vs;
  wire [1:0]   sinkVec_queue_53_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_53 = {sinkVec_queue_53_enq_bits_vs, sinkVec_queue_53_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_53 = {sinkVec_queue_dataIn_hi_53, sinkVec_queue_dataIn_lo_53};
  wire [2:0]   sinkVec_queue_dataOut_53_instructionIndex = _sinkVec_queue_fifo_53_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_53_offset = _sinkVec_queue_fifo_53_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_53_readSource = _sinkVec_queue_fifo_53_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_53_vs = _sinkVec_queue_fifo_53_data_out[11:7];
  wire         sinkVec_queue_53_enq_ready = ~_sinkVec_queue_fifo_53_full;
  wire         sinkVec_queue_53_enq_valid;
  assign sinkVec_queue_53_deq_valid = ~_sinkVec_queue_fifo_53_empty | sinkVec_queue_53_enq_valid;
  assign sinkVec_queue_53_deq_bits_vs = _sinkVec_queue_fifo_53_empty ? sinkVec_queue_53_enq_bits_vs : sinkVec_queue_dataOut_53_vs;
  assign sinkVec_queue_53_deq_bits_readSource = _sinkVec_queue_fifo_53_empty ? sinkVec_queue_53_enq_bits_readSource : sinkVec_queue_dataOut_53_readSource;
  assign sinkVec_queue_53_deq_bits_offset = _sinkVec_queue_fifo_53_empty ? sinkVec_queue_53_enq_bits_offset : sinkVec_queue_dataOut_53_offset;
  assign sinkVec_queue_53_deq_bits_instructionIndex = _sinkVec_queue_fifo_53_empty ? sinkVec_queue_53_enq_bits_instructionIndex : sinkVec_queue_dataOut_53_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_53;
  wire         sinkVec_releasePipe_pipe_out_53_valid = sinkVec_releasePipe_pipe_v_53;
  wire         x13_13_1_ready;
  wire         x13_13_1_valid;
  wire         sinkVec_validSource_53_valid = x13_13_1_ready & x13_13_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_53;
  wire [2:0]   sinkVec_tokenCheck_counterChange_53 = sinkVec_validSource_53_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_53 = ~(sinkVec_tokenCheck_counter_53[2]);
  assign x13_13_1_ready = sinkVec_tokenCheck_53;
  assign sinkVec_queue_53_enq_valid = sinkVec_validSink_53_valid;
  assign sinkVec_queue_53_enq_bits_vs = sinkVec_validSink_53_bits_vs;
  assign sinkVec_queue_53_enq_bits_readSource = sinkVec_validSink_53_bits_readSource;
  assign sinkVec_queue_53_enq_bits_offset = sinkVec_validSink_53_bits_offset;
  assign sinkVec_queue_53_enq_bits_instructionIndex = sinkVec_validSink_53_bits_instructionIndex;
  reg          sinkVec_shifterReg_53_0_valid;
  assign sinkVec_validSink_53_valid = sinkVec_shifterReg_53_0_valid;
  reg  [4:0]   sinkVec_shifterReg_53_0_bits_vs;
  assign sinkVec_validSink_53_bits_vs = sinkVec_shifterReg_53_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_53_0_bits_readSource;
  assign sinkVec_validSink_53_bits_readSource = sinkVec_shifterReg_53_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_53_0_bits_offset;
  assign sinkVec_validSink_53_bits_offset = sinkVec_shifterReg_53_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_53_0_bits_instructionIndex;
  assign sinkVec_validSink_53_bits_instructionIndex = sinkVec_shifterReg_53_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_53 = sinkVec_shifterReg_53_0_valid | sinkVec_validSource_53_valid;
  assign sinkVec_sinkWire_52_ready = sinkVec_26_0_ready;
  assign sinkVec_sinkWire_53_ready = sinkVec_26_1_ready;
  reg          maskUnitFirst_26;
  wire         tryToRead_26 = sinkVec_26_0_valid | sinkVec_26_1_valid;
  wire         sinkWire_26_valid = maskUnitFirst_26 ? sinkVec_26_0_valid : sinkVec_26_1_valid;
  wire [4:0]   sinkWire_26_bits_vs = maskUnitFirst_26 ? sinkVec_26_0_bits_vs : sinkVec_26_1_bits_vs;
  wire [1:0]   sinkWire_26_bits_readSource = maskUnitFirst_26 ? sinkVec_26_0_bits_readSource : sinkVec_26_1_bits_readSource;
  wire [1:0]   sinkWire_26_bits_offset = maskUnitFirst_26 ? sinkVec_26_0_bits_offset : sinkVec_26_1_bits_offset;
  wire [2:0]   sinkWire_26_bits_instructionIndex = maskUnitFirst_26 ? sinkVec_26_0_bits_instructionIndex : sinkVec_26_1_bits_instructionIndex;
  wire         sinkWire_26_ready;
  assign sinkVec_26_1_ready = sinkWire_26_ready & ~maskUnitFirst_26;
  assign sinkVec_26_0_ready = sinkWire_26_ready & maskUnitFirst_26;
  reg          accessDataValid_pipe_v_26;
  reg          accessDataValid_pipe_pipe_v_26;
  wire         accessDataValid_pipe_pipe_out_26_valid = accessDataValid_pipe_pipe_v_26;
  wire         accessDataSource_26_valid = accessDataValid_pipe_pipe_out_26_valid;
  reg          shifterReg_42_0_valid;
  reg  [31:0]  shifterReg_42_0_bits;
  wire         shifterValid_42 = shifterReg_42_0_valid | accessDataSource_26_valid;
  reg          accessDataValid_pipe_v_27;
  reg          accessDataValid_pipe_pipe_v_27;
  wire         accessDataValid_pipe_pipe_out_27_valid = accessDataValid_pipe_pipe_v_27;
  wire         accessDataSource_27_valid = accessDataValid_pipe_pipe_out_27_valid;
  reg          shifterReg_43_0_valid;
  reg  [31:0]  shifterReg_43_0_bits;
  wire         shifterValid_43 = shifterReg_43_0_valid | accessDataSource_27_valid;
  wire         sinkVec_tokenCheck_54;
  wire [4:0]   sinkVec_validSource_54_bits_vd = x22_13_0_bits_vd;
  wire [1:0]   sinkVec_validSource_54_bits_offset = x22_13_0_bits_offset;
  wire [3:0]   sinkVec_validSource_54_bits_mask = x22_13_0_bits_mask;
  wire [31:0]  sinkVec_validSource_54_bits_data = x22_13_0_bits_data;
  wire [2:0]   sinkVec_validSource_54_bits_instructionIndex = x22_13_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_55;
  wire [4:0]   sinkVec_validSource_55_bits_vd = x22_13_1_bits_vd;
  wire [1:0]   sinkVec_validSource_55_bits_offset = x22_13_1_bits_offset;
  wire [3:0]   sinkVec_validSource_55_bits_mask = x22_13_1_bits_mask;
  wire [31:0]  sinkVec_validSource_55_bits_data = x22_13_1_bits_data;
  wire         sinkVec_validSource_55_bits_last = x22_13_1_bits_last;
  wire [2:0]   sinkVec_validSource_55_bits_instructionIndex = x22_13_1_bits_instructionIndex;
  wire         sinkVec_27_0_ready;
  wire         sinkVec_queue_54_deq_ready = sinkVec_sinkWire_54_ready;
  wire         sinkVec_queue_54_deq_valid;
  wire [4:0]   sinkVec_queue_54_deq_bits_vd;
  wire         sinkVec_27_0_valid = sinkVec_sinkWire_54_valid;
  wire [1:0]   sinkVec_queue_54_deq_bits_offset;
  wire [4:0]   sinkVec_27_0_bits_vd = sinkVec_sinkWire_54_bits_vd;
  wire [3:0]   sinkVec_queue_54_deq_bits_mask;
  wire [1:0]   sinkVec_27_0_bits_offset = sinkVec_sinkWire_54_bits_offset;
  wire [31:0]  sinkVec_queue_54_deq_bits_data;
  wire [3:0]   sinkVec_27_0_bits_mask = sinkVec_sinkWire_54_bits_mask;
  wire         sinkVec_queue_54_deq_bits_last;
  wire [31:0]  sinkVec_27_0_bits_data = sinkVec_sinkWire_54_bits_data;
  wire [2:0]   sinkVec_queue_54_deq_bits_instructionIndex;
  wire         sinkVec_27_0_bits_last = sinkVec_sinkWire_54_bits_last;
  wire [2:0]   sinkVec_27_0_bits_instructionIndex = sinkVec_sinkWire_54_bits_instructionIndex;
  wire         sinkVec_validSink_54_valid;
  wire [4:0]   sinkVec_validSink_54_bits_vd;
  wire [1:0]   sinkVec_validSink_54_bits_offset;
  wire [3:0]   sinkVec_validSink_54_bits_mask;
  wire [31:0]  sinkVec_validSink_54_bits_data;
  wire [2:0]   sinkVec_validSink_54_bits_instructionIndex;
  assign sinkVec_sinkWire_54_valid = sinkVec_queue_54_deq_valid;
  assign sinkVec_sinkWire_54_bits_vd = sinkVec_queue_54_deq_bits_vd;
  assign sinkVec_sinkWire_54_bits_offset = sinkVec_queue_54_deq_bits_offset;
  assign sinkVec_sinkWire_54_bits_mask = sinkVec_queue_54_deq_bits_mask;
  assign sinkVec_sinkWire_54_bits_data = sinkVec_queue_54_deq_bits_data;
  assign sinkVec_sinkWire_54_bits_last = sinkVec_queue_54_deq_bits_last;
  assign sinkVec_sinkWire_54_bits_instructionIndex = sinkVec_queue_54_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_54_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_26 = {sinkVec_queue_54_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_54_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_54 = {sinkVec_queue_dataIn_lo_hi_26, sinkVec_queue_54_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_54_enq_bits_vd;
  wire [1:0]   sinkVec_queue_54_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_26 = {sinkVec_queue_54_enq_bits_vd, sinkVec_queue_54_enq_bits_offset};
  wire [3:0]   sinkVec_queue_54_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_54 = {sinkVec_queue_dataIn_hi_hi_26, sinkVec_queue_54_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_54 = {sinkVec_queue_dataIn_hi_54, sinkVec_queue_dataIn_lo_54};
  wire [2:0]   sinkVec_queue_dataOut_54_instructionIndex = _sinkVec_queue_fifo_54_data_out[2:0];
  wire         sinkVec_queue_dataOut_54_last = _sinkVec_queue_fifo_54_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_54_data = _sinkVec_queue_fifo_54_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_54_mask = _sinkVec_queue_fifo_54_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_54_offset = _sinkVec_queue_fifo_54_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_54_vd = _sinkVec_queue_fifo_54_data_out[46:42];
  wire         sinkVec_queue_54_enq_ready = ~_sinkVec_queue_fifo_54_full;
  wire         sinkVec_queue_54_enq_valid;
  assign sinkVec_queue_54_deq_valid = ~_sinkVec_queue_fifo_54_empty | sinkVec_queue_54_enq_valid;
  assign sinkVec_queue_54_deq_bits_vd = _sinkVec_queue_fifo_54_empty ? sinkVec_queue_54_enq_bits_vd : sinkVec_queue_dataOut_54_vd;
  assign sinkVec_queue_54_deq_bits_offset = _sinkVec_queue_fifo_54_empty ? sinkVec_queue_54_enq_bits_offset : sinkVec_queue_dataOut_54_offset;
  assign sinkVec_queue_54_deq_bits_mask = _sinkVec_queue_fifo_54_empty ? sinkVec_queue_54_enq_bits_mask : sinkVec_queue_dataOut_54_mask;
  assign sinkVec_queue_54_deq_bits_data = _sinkVec_queue_fifo_54_empty ? sinkVec_queue_54_enq_bits_data : sinkVec_queue_dataOut_54_data;
  assign sinkVec_queue_54_deq_bits_last = ~_sinkVec_queue_fifo_54_empty & sinkVec_queue_dataOut_54_last;
  assign sinkVec_queue_54_deq_bits_instructionIndex = _sinkVec_queue_fifo_54_empty ? sinkVec_queue_54_enq_bits_instructionIndex : sinkVec_queue_dataOut_54_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_54;
  wire         sinkVec_releasePipe_pipe_out_54_valid = sinkVec_releasePipe_pipe_v_54;
  wire         x22_13_0_ready;
  wire         x22_13_0_valid;
  wire         sinkVec_validSource_54_valid = x22_13_0_ready & x22_13_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_54;
  wire [2:0]   sinkVec_tokenCheck_counterChange_54 = sinkVec_validSource_54_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_54 = ~(sinkVec_tokenCheck_counter_54[2]);
  assign x22_13_0_ready = sinkVec_tokenCheck_54;
  assign sinkVec_queue_54_enq_valid = sinkVec_validSink_54_valid;
  assign sinkVec_queue_54_enq_bits_vd = sinkVec_validSink_54_bits_vd;
  assign sinkVec_queue_54_enq_bits_offset = sinkVec_validSink_54_bits_offset;
  assign sinkVec_queue_54_enq_bits_mask = sinkVec_validSink_54_bits_mask;
  assign sinkVec_queue_54_enq_bits_data = sinkVec_validSink_54_bits_data;
  assign sinkVec_queue_54_enq_bits_instructionIndex = sinkVec_validSink_54_bits_instructionIndex;
  reg          sinkVec_shifterReg_54_0_valid;
  assign sinkVec_validSink_54_valid = sinkVec_shifterReg_54_0_valid;
  reg  [4:0]   sinkVec_shifterReg_54_0_bits_vd;
  assign sinkVec_validSink_54_bits_vd = sinkVec_shifterReg_54_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_54_0_bits_offset;
  assign sinkVec_validSink_54_bits_offset = sinkVec_shifterReg_54_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_54_0_bits_mask;
  assign sinkVec_validSink_54_bits_mask = sinkVec_shifterReg_54_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_54_0_bits_data;
  assign sinkVec_validSink_54_bits_data = sinkVec_shifterReg_54_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_54_0_bits_instructionIndex;
  assign sinkVec_validSink_54_bits_instructionIndex = sinkVec_shifterReg_54_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_54 = sinkVec_shifterReg_54_0_valid | sinkVec_validSource_54_valid;
  wire         sinkVec_27_1_ready;
  wire         sinkVec_queue_55_deq_ready = sinkVec_sinkWire_55_ready;
  wire         sinkVec_queue_55_deq_valid;
  wire [4:0]   sinkVec_queue_55_deq_bits_vd;
  wire         sinkVec_27_1_valid = sinkVec_sinkWire_55_valid;
  wire [1:0]   sinkVec_queue_55_deq_bits_offset;
  wire [4:0]   sinkVec_27_1_bits_vd = sinkVec_sinkWire_55_bits_vd;
  wire [3:0]   sinkVec_queue_55_deq_bits_mask;
  wire [1:0]   sinkVec_27_1_bits_offset = sinkVec_sinkWire_55_bits_offset;
  wire [31:0]  sinkVec_queue_55_deq_bits_data;
  wire [3:0]   sinkVec_27_1_bits_mask = sinkVec_sinkWire_55_bits_mask;
  wire         sinkVec_queue_55_deq_bits_last;
  wire [31:0]  sinkVec_27_1_bits_data = sinkVec_sinkWire_55_bits_data;
  wire [2:0]   sinkVec_queue_55_deq_bits_instructionIndex;
  wire         sinkVec_27_1_bits_last = sinkVec_sinkWire_55_bits_last;
  wire [2:0]   sinkVec_27_1_bits_instructionIndex = sinkVec_sinkWire_55_bits_instructionIndex;
  wire         sinkVec_validSink_55_valid;
  wire [4:0]   sinkVec_validSink_55_bits_vd;
  wire [1:0]   sinkVec_validSink_55_bits_offset;
  wire [3:0]   sinkVec_validSink_55_bits_mask;
  wire [31:0]  sinkVec_validSink_55_bits_data;
  wire         sinkVec_validSink_55_bits_last;
  wire [2:0]   sinkVec_validSink_55_bits_instructionIndex;
  assign sinkVec_sinkWire_55_valid = sinkVec_queue_55_deq_valid;
  assign sinkVec_sinkWire_55_bits_vd = sinkVec_queue_55_deq_bits_vd;
  assign sinkVec_sinkWire_55_bits_offset = sinkVec_queue_55_deq_bits_offset;
  assign sinkVec_sinkWire_55_bits_mask = sinkVec_queue_55_deq_bits_mask;
  assign sinkVec_sinkWire_55_bits_data = sinkVec_queue_55_deq_bits_data;
  assign sinkVec_sinkWire_55_bits_last = sinkVec_queue_55_deq_bits_last;
  assign sinkVec_sinkWire_55_bits_instructionIndex = sinkVec_queue_55_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_55_enq_bits_data;
  wire         sinkVec_queue_55_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_27 = {sinkVec_queue_55_enq_bits_data, sinkVec_queue_55_enq_bits_last};
  wire [2:0]   sinkVec_queue_55_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_55 = {sinkVec_queue_dataIn_lo_hi_27, sinkVec_queue_55_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_55_enq_bits_vd;
  wire [1:0]   sinkVec_queue_55_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_27 = {sinkVec_queue_55_enq_bits_vd, sinkVec_queue_55_enq_bits_offset};
  wire [3:0]   sinkVec_queue_55_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_55 = {sinkVec_queue_dataIn_hi_hi_27, sinkVec_queue_55_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_55 = {sinkVec_queue_dataIn_hi_55, sinkVec_queue_dataIn_lo_55};
  wire [2:0]   sinkVec_queue_dataOut_55_instructionIndex = _sinkVec_queue_fifo_55_data_out[2:0];
  wire         sinkVec_queue_dataOut_55_last = _sinkVec_queue_fifo_55_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_55_data = _sinkVec_queue_fifo_55_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_55_mask = _sinkVec_queue_fifo_55_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_55_offset = _sinkVec_queue_fifo_55_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_55_vd = _sinkVec_queue_fifo_55_data_out[46:42];
  wire         sinkVec_queue_55_enq_ready = ~_sinkVec_queue_fifo_55_full;
  wire         sinkVec_queue_55_enq_valid;
  assign sinkVec_queue_55_deq_valid = ~_sinkVec_queue_fifo_55_empty | sinkVec_queue_55_enq_valid;
  assign sinkVec_queue_55_deq_bits_vd = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_vd : sinkVec_queue_dataOut_55_vd;
  assign sinkVec_queue_55_deq_bits_offset = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_offset : sinkVec_queue_dataOut_55_offset;
  assign sinkVec_queue_55_deq_bits_mask = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_mask : sinkVec_queue_dataOut_55_mask;
  assign sinkVec_queue_55_deq_bits_data = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_data : sinkVec_queue_dataOut_55_data;
  assign sinkVec_queue_55_deq_bits_last = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_last : sinkVec_queue_dataOut_55_last;
  assign sinkVec_queue_55_deq_bits_instructionIndex = _sinkVec_queue_fifo_55_empty ? sinkVec_queue_55_enq_bits_instructionIndex : sinkVec_queue_dataOut_55_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_55;
  wire         sinkVec_releasePipe_pipe_out_55_valid = sinkVec_releasePipe_pipe_v_55;
  wire         x22_13_1_ready;
  wire         x22_13_1_valid;
  wire         sinkVec_validSource_55_valid = x22_13_1_ready & x22_13_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_55;
  wire [2:0]   sinkVec_tokenCheck_counterChange_55 = sinkVec_validSource_55_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_55 = ~(sinkVec_tokenCheck_counter_55[2]);
  assign x22_13_1_ready = sinkVec_tokenCheck_55;
  assign sinkVec_queue_55_enq_valid = sinkVec_validSink_55_valid;
  assign sinkVec_queue_55_enq_bits_vd = sinkVec_validSink_55_bits_vd;
  assign sinkVec_queue_55_enq_bits_offset = sinkVec_validSink_55_bits_offset;
  assign sinkVec_queue_55_enq_bits_mask = sinkVec_validSink_55_bits_mask;
  assign sinkVec_queue_55_enq_bits_data = sinkVec_validSink_55_bits_data;
  assign sinkVec_queue_55_enq_bits_last = sinkVec_validSink_55_bits_last;
  assign sinkVec_queue_55_enq_bits_instructionIndex = sinkVec_validSink_55_bits_instructionIndex;
  reg          sinkVec_shifterReg_55_0_valid;
  assign sinkVec_validSink_55_valid = sinkVec_shifterReg_55_0_valid;
  reg  [4:0]   sinkVec_shifterReg_55_0_bits_vd;
  assign sinkVec_validSink_55_bits_vd = sinkVec_shifterReg_55_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_55_0_bits_offset;
  assign sinkVec_validSink_55_bits_offset = sinkVec_shifterReg_55_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_55_0_bits_mask;
  assign sinkVec_validSink_55_bits_mask = sinkVec_shifterReg_55_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_55_0_bits_data;
  assign sinkVec_validSink_55_bits_data = sinkVec_shifterReg_55_0_bits_data;
  reg          sinkVec_shifterReg_55_0_bits_last;
  assign sinkVec_validSink_55_bits_last = sinkVec_shifterReg_55_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_55_0_bits_instructionIndex;
  assign sinkVec_validSink_55_bits_instructionIndex = sinkVec_shifterReg_55_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_55 = sinkVec_shifterReg_55_0_valid | sinkVec_validSource_55_valid;
  assign sinkVec_sinkWire_54_ready = sinkVec_27_0_ready;
  assign sinkVec_sinkWire_55_ready = sinkVec_27_1_ready;
  reg          maskUnitFirst_27;
  wire         tryToRead_27 = sinkVec_27_0_valid | sinkVec_27_1_valid;
  wire         sinkWire_27_valid = maskUnitFirst_27 ? sinkVec_27_0_valid : sinkVec_27_1_valid;
  wire [4:0]   sinkWire_27_bits_vd = maskUnitFirst_27 ? sinkVec_27_0_bits_vd : sinkVec_27_1_bits_vd;
  wire [1:0]   sinkWire_27_bits_offset = maskUnitFirst_27 ? sinkVec_27_0_bits_offset : sinkVec_27_1_bits_offset;
  wire [3:0]   sinkWire_27_bits_mask = maskUnitFirst_27 ? sinkVec_27_0_bits_mask : sinkVec_27_1_bits_mask;
  wire [31:0]  sinkWire_27_bits_data = maskUnitFirst_27 ? sinkVec_27_0_bits_data : sinkVec_27_1_bits_data;
  wire         sinkWire_27_bits_last = maskUnitFirst_27 ? sinkVec_27_0_bits_last : sinkVec_27_1_bits_last;
  wire [2:0]   sinkWire_27_bits_instructionIndex = maskUnitFirst_27 ? sinkVec_27_0_bits_instructionIndex : sinkVec_27_1_bits_instructionIndex;
  wire         sinkWire_27_ready;
  assign sinkVec_27_1_ready = sinkWire_27_ready & ~maskUnitFirst_27;
  assign sinkVec_27_0_ready = sinkWire_27_ready & maskUnitFirst_27;
  reg          view__writeRelease_13_pipe_v;
  wire         view__writeRelease_13_pipe_out_valid = view__writeRelease_13_pipe_v;
  reg          pipe_v_39;
  wire         pipe_out_26_valid = pipe_v_39;
  wire         _probeWire_writeQueueEnqVec_13_valid_T = x22_13_0_ready & _maskUnit_exeResp_13_valid;
  reg          instructionFinishedPipe_pipe_v_13;
  wire         instructionFinishedPipe_pipe_out_13_valid = instructionFinishedPipe_pipe_v_13;
  reg  [7:0]   instructionFinishedPipe_pipe_b_13;
  wire [7:0]   instructionFinishedPipe_pipe_out_13_bits = instructionFinishedPipe_pipe_b_13;
  wire         instructionFinished_13_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_13_bits);
  wire         instructionFinished_13_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_13_bits);
  wire         instructionFinished_13_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_13_bits);
  wire         instructionFinished_13_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_13_bits);
  assign vxsatReportVec_13 = _laneVec_13_vxsatReport[3:0];
  reg          pipe_v_40;
  reg  [31:0]  pipe_b_40;
  reg          pipe_pipe_v_13;
  wire         pipe_pipe_out_13_valid = pipe_pipe_v_13;
  reg  [31:0]  pipe_pipe_b_13;
  wire [31:0]  pipe_pipe_out_13_bits = pipe_pipe_b_13;
  reg          view__laneMaskSelect_13_pipe_v;
  reg  [5:0]   view__laneMaskSelect_13_pipe_b;
  reg          view__laneMaskSelect_13_pipe_pipe_v;
  wire         view__laneMaskSelect_13_pipe_pipe_out_valid = view__laneMaskSelect_13_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_13_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_13_pipe_pipe_out_bits = view__laneMaskSelect_13_pipe_pipe_b;
  reg          view__laneMaskSewSelect_13_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_13_pipe_b;
  reg          view__laneMaskSewSelect_13_pipe_pipe_v;
  wire         view__laneMaskSewSelect_13_pipe_pipe_out_valid = view__laneMaskSewSelect_13_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_13_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_13_pipe_pipe_out_bits = view__laneMaskSewSelect_13_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_13;
  wire         lsuLastPipe_pipe_out_13_valid = lsuLastPipe_pipe_v_13;
  reg  [7:0]   lsuLastPipe_pipe_b_13;
  wire [7:0]   lsuLastPipe_pipe_out_13_bits = lsuLastPipe_pipe_b_13;
  reg          maskLastPipe_pipe_v_13;
  wire         maskLastPipe_pipe_out_13_valid = maskLastPipe_pipe_v_13;
  reg  [7:0]   maskLastPipe_pipe_b_13;
  wire [7:0]   maskLastPipe_pipe_out_13_bits = maskLastPipe_pipe_b_13;
  wire [5:0]   writeCounter_13 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h34};
  reg          pipe_v_41;
  wire         pipe_out_27_valid = pipe_v_41;
  reg  [5:0]   pipe_b_41;
  wire [5:0]   pipe_out_27_bits = pipe_b_41;
  assign laneRequestSinkWire_14_ready = ~laneRequestSinkWire_14_bits_issueInst | _laneVec_14_laneRequest_ready;
  wire         sinkVec_tokenCheck_56;
  wire [4:0]   sinkVec_validSource_56_bits_vs = x13_14_0_bits_vs;
  wire [1:0]   sinkVec_validSource_56_bits_offset = x13_14_0_bits_offset;
  wire [2:0]   sinkVec_validSource_56_bits_instructionIndex = x13_14_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_57;
  wire [4:0]   sinkVec_validSource_57_bits_vs = x13_14_1_bits_vs;
  wire [1:0]   sinkVec_validSource_57_bits_offset = x13_14_1_bits_offset;
  wire [2:0]   sinkVec_validSource_57_bits_instructionIndex = x13_14_1_bits_instructionIndex;
  wire         sinkVec_28_0_ready;
  wire         sinkVec_queue_56_deq_ready = sinkVec_sinkWire_56_ready;
  wire         sinkVec_queue_56_deq_valid;
  wire [4:0]   sinkVec_queue_56_deq_bits_vs;
  wire         sinkVec_28_0_valid = sinkVec_sinkWire_56_valid;
  wire [1:0]   sinkVec_queue_56_deq_bits_readSource;
  wire [4:0]   sinkVec_28_0_bits_vs = sinkVec_sinkWire_56_bits_vs;
  wire [1:0]   sinkVec_queue_56_deq_bits_offset;
  wire [1:0]   sinkVec_28_0_bits_readSource = sinkVec_sinkWire_56_bits_readSource;
  wire [2:0]   sinkVec_queue_56_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_28_0_bits_offset = sinkVec_sinkWire_56_bits_offset;
  wire [2:0]   sinkVec_28_0_bits_instructionIndex = sinkVec_sinkWire_56_bits_instructionIndex;
  wire         sinkVec_validSink_56_valid;
  wire [4:0]   sinkVec_validSink_56_bits_vs;
  wire [1:0]   sinkVec_validSink_56_bits_readSource;
  wire [1:0]   sinkVec_validSink_56_bits_offset;
  wire [2:0]   sinkVec_validSink_56_bits_instructionIndex;
  assign sinkVec_sinkWire_56_valid = sinkVec_queue_56_deq_valid;
  assign sinkVec_sinkWire_56_bits_vs = sinkVec_queue_56_deq_bits_vs;
  assign sinkVec_sinkWire_56_bits_readSource = sinkVec_queue_56_deq_bits_readSource;
  assign sinkVec_sinkWire_56_bits_offset = sinkVec_queue_56_deq_bits_offset;
  assign sinkVec_sinkWire_56_bits_instructionIndex = sinkVec_queue_56_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_56_enq_bits_offset;
  wire [2:0]   sinkVec_queue_56_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_56 = {sinkVec_queue_56_enq_bits_offset, sinkVec_queue_56_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_56_enq_bits_vs;
  wire [1:0]   sinkVec_queue_56_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_56 = {sinkVec_queue_56_enq_bits_vs, sinkVec_queue_56_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_56 = {sinkVec_queue_dataIn_hi_56, sinkVec_queue_dataIn_lo_56};
  wire [2:0]   sinkVec_queue_dataOut_56_instructionIndex = _sinkVec_queue_fifo_56_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_56_offset = _sinkVec_queue_fifo_56_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_56_readSource = _sinkVec_queue_fifo_56_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_56_vs = _sinkVec_queue_fifo_56_data_out[11:7];
  wire         sinkVec_queue_56_enq_ready = ~_sinkVec_queue_fifo_56_full;
  wire         sinkVec_queue_56_enq_valid;
  assign sinkVec_queue_56_deq_valid = ~_sinkVec_queue_fifo_56_empty | sinkVec_queue_56_enq_valid;
  assign sinkVec_queue_56_deq_bits_vs = _sinkVec_queue_fifo_56_empty ? sinkVec_queue_56_enq_bits_vs : sinkVec_queue_dataOut_56_vs;
  assign sinkVec_queue_56_deq_bits_readSource = _sinkVec_queue_fifo_56_empty ? sinkVec_queue_56_enq_bits_readSource : sinkVec_queue_dataOut_56_readSource;
  assign sinkVec_queue_56_deq_bits_offset = _sinkVec_queue_fifo_56_empty ? sinkVec_queue_56_enq_bits_offset : sinkVec_queue_dataOut_56_offset;
  assign sinkVec_queue_56_deq_bits_instructionIndex = _sinkVec_queue_fifo_56_empty ? sinkVec_queue_56_enq_bits_instructionIndex : sinkVec_queue_dataOut_56_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_56;
  wire         sinkVec_releasePipe_pipe_out_56_valid = sinkVec_releasePipe_pipe_v_56;
  wire         x13_14_0_ready;
  wire         x13_14_0_valid;
  wire         sinkVec_validSource_56_valid = x13_14_0_ready & x13_14_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_56;
  wire [2:0]   sinkVec_tokenCheck_counterChange_56 = sinkVec_validSource_56_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_56 = ~(sinkVec_tokenCheck_counter_56[2]);
  assign x13_14_0_ready = sinkVec_tokenCheck_56;
  assign sinkVec_queue_56_enq_valid = sinkVec_validSink_56_valid;
  assign sinkVec_queue_56_enq_bits_vs = sinkVec_validSink_56_bits_vs;
  assign sinkVec_queue_56_enq_bits_readSource = sinkVec_validSink_56_bits_readSource;
  assign sinkVec_queue_56_enq_bits_offset = sinkVec_validSink_56_bits_offset;
  assign sinkVec_queue_56_enq_bits_instructionIndex = sinkVec_validSink_56_bits_instructionIndex;
  reg          sinkVec_shifterReg_56_0_valid;
  assign sinkVec_validSink_56_valid = sinkVec_shifterReg_56_0_valid;
  reg  [4:0]   sinkVec_shifterReg_56_0_bits_vs;
  assign sinkVec_validSink_56_bits_vs = sinkVec_shifterReg_56_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_56_0_bits_readSource;
  assign sinkVec_validSink_56_bits_readSource = sinkVec_shifterReg_56_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_56_0_bits_offset;
  assign sinkVec_validSink_56_bits_offset = sinkVec_shifterReg_56_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_56_0_bits_instructionIndex;
  assign sinkVec_validSink_56_bits_instructionIndex = sinkVec_shifterReg_56_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_56 = sinkVec_shifterReg_56_0_valid | sinkVec_validSource_56_valid;
  wire         sinkVec_28_1_ready;
  wire         sinkVec_queue_57_deq_ready = sinkVec_sinkWire_57_ready;
  wire         sinkVec_queue_57_deq_valid;
  wire [4:0]   sinkVec_queue_57_deq_bits_vs;
  wire         sinkVec_28_1_valid = sinkVec_sinkWire_57_valid;
  wire [1:0]   sinkVec_queue_57_deq_bits_readSource;
  wire [4:0]   sinkVec_28_1_bits_vs = sinkVec_sinkWire_57_bits_vs;
  wire [1:0]   sinkVec_queue_57_deq_bits_offset;
  wire [1:0]   sinkVec_28_1_bits_readSource = sinkVec_sinkWire_57_bits_readSource;
  wire [2:0]   sinkVec_queue_57_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_28_1_bits_offset = sinkVec_sinkWire_57_bits_offset;
  wire [2:0]   sinkVec_28_1_bits_instructionIndex = sinkVec_sinkWire_57_bits_instructionIndex;
  wire         sinkVec_validSink_57_valid;
  wire [4:0]   sinkVec_validSink_57_bits_vs;
  wire [1:0]   sinkVec_validSink_57_bits_readSource;
  wire [1:0]   sinkVec_validSink_57_bits_offset;
  wire [2:0]   sinkVec_validSink_57_bits_instructionIndex;
  assign sinkVec_sinkWire_57_valid = sinkVec_queue_57_deq_valid;
  assign sinkVec_sinkWire_57_bits_vs = sinkVec_queue_57_deq_bits_vs;
  assign sinkVec_sinkWire_57_bits_readSource = sinkVec_queue_57_deq_bits_readSource;
  assign sinkVec_sinkWire_57_bits_offset = sinkVec_queue_57_deq_bits_offset;
  assign sinkVec_sinkWire_57_bits_instructionIndex = sinkVec_queue_57_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_57_enq_bits_offset;
  wire [2:0]   sinkVec_queue_57_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_57 = {sinkVec_queue_57_enq_bits_offset, sinkVec_queue_57_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_57_enq_bits_vs;
  wire [1:0]   sinkVec_queue_57_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_57 = {sinkVec_queue_57_enq_bits_vs, sinkVec_queue_57_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_57 = {sinkVec_queue_dataIn_hi_57, sinkVec_queue_dataIn_lo_57};
  wire [2:0]   sinkVec_queue_dataOut_57_instructionIndex = _sinkVec_queue_fifo_57_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_57_offset = _sinkVec_queue_fifo_57_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_57_readSource = _sinkVec_queue_fifo_57_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_57_vs = _sinkVec_queue_fifo_57_data_out[11:7];
  wire         sinkVec_queue_57_enq_ready = ~_sinkVec_queue_fifo_57_full;
  wire         sinkVec_queue_57_enq_valid;
  assign sinkVec_queue_57_deq_valid = ~_sinkVec_queue_fifo_57_empty | sinkVec_queue_57_enq_valid;
  assign sinkVec_queue_57_deq_bits_vs = _sinkVec_queue_fifo_57_empty ? sinkVec_queue_57_enq_bits_vs : sinkVec_queue_dataOut_57_vs;
  assign sinkVec_queue_57_deq_bits_readSource = _sinkVec_queue_fifo_57_empty ? sinkVec_queue_57_enq_bits_readSource : sinkVec_queue_dataOut_57_readSource;
  assign sinkVec_queue_57_deq_bits_offset = _sinkVec_queue_fifo_57_empty ? sinkVec_queue_57_enq_bits_offset : sinkVec_queue_dataOut_57_offset;
  assign sinkVec_queue_57_deq_bits_instructionIndex = _sinkVec_queue_fifo_57_empty ? sinkVec_queue_57_enq_bits_instructionIndex : sinkVec_queue_dataOut_57_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_57;
  wire         sinkVec_releasePipe_pipe_out_57_valid = sinkVec_releasePipe_pipe_v_57;
  wire         x13_14_1_ready;
  wire         x13_14_1_valid;
  wire         sinkVec_validSource_57_valid = x13_14_1_ready & x13_14_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_57;
  wire [2:0]   sinkVec_tokenCheck_counterChange_57 = sinkVec_validSource_57_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_57 = ~(sinkVec_tokenCheck_counter_57[2]);
  assign x13_14_1_ready = sinkVec_tokenCheck_57;
  assign sinkVec_queue_57_enq_valid = sinkVec_validSink_57_valid;
  assign sinkVec_queue_57_enq_bits_vs = sinkVec_validSink_57_bits_vs;
  assign sinkVec_queue_57_enq_bits_readSource = sinkVec_validSink_57_bits_readSource;
  assign sinkVec_queue_57_enq_bits_offset = sinkVec_validSink_57_bits_offset;
  assign sinkVec_queue_57_enq_bits_instructionIndex = sinkVec_validSink_57_bits_instructionIndex;
  reg          sinkVec_shifterReg_57_0_valid;
  assign sinkVec_validSink_57_valid = sinkVec_shifterReg_57_0_valid;
  reg  [4:0]   sinkVec_shifterReg_57_0_bits_vs;
  assign sinkVec_validSink_57_bits_vs = sinkVec_shifterReg_57_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_57_0_bits_readSource;
  assign sinkVec_validSink_57_bits_readSource = sinkVec_shifterReg_57_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_57_0_bits_offset;
  assign sinkVec_validSink_57_bits_offset = sinkVec_shifterReg_57_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_57_0_bits_instructionIndex;
  assign sinkVec_validSink_57_bits_instructionIndex = sinkVec_shifterReg_57_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_57 = sinkVec_shifterReg_57_0_valid | sinkVec_validSource_57_valid;
  assign sinkVec_sinkWire_56_ready = sinkVec_28_0_ready;
  assign sinkVec_sinkWire_57_ready = sinkVec_28_1_ready;
  reg          maskUnitFirst_28;
  wire         tryToRead_28 = sinkVec_28_0_valid | sinkVec_28_1_valid;
  wire         sinkWire_28_valid = maskUnitFirst_28 ? sinkVec_28_0_valid : sinkVec_28_1_valid;
  wire [4:0]   sinkWire_28_bits_vs = maskUnitFirst_28 ? sinkVec_28_0_bits_vs : sinkVec_28_1_bits_vs;
  wire [1:0]   sinkWire_28_bits_readSource = maskUnitFirst_28 ? sinkVec_28_0_bits_readSource : sinkVec_28_1_bits_readSource;
  wire [1:0]   sinkWire_28_bits_offset = maskUnitFirst_28 ? sinkVec_28_0_bits_offset : sinkVec_28_1_bits_offset;
  wire [2:0]   sinkWire_28_bits_instructionIndex = maskUnitFirst_28 ? sinkVec_28_0_bits_instructionIndex : sinkVec_28_1_bits_instructionIndex;
  wire         sinkWire_28_ready;
  assign sinkVec_28_1_ready = sinkWire_28_ready & ~maskUnitFirst_28;
  assign sinkVec_28_0_ready = sinkWire_28_ready & maskUnitFirst_28;
  reg          accessDataValid_pipe_v_28;
  reg          accessDataValid_pipe_pipe_v_28;
  wire         accessDataValid_pipe_pipe_out_28_valid = accessDataValid_pipe_pipe_v_28;
  wire         accessDataSource_28_valid = accessDataValid_pipe_pipe_out_28_valid;
  reg          shifterReg_44_0_valid;
  reg  [31:0]  shifterReg_44_0_bits;
  wire         shifterValid_44 = shifterReg_44_0_valid | accessDataSource_28_valid;
  reg          accessDataValid_pipe_v_29;
  reg          accessDataValid_pipe_pipe_v_29;
  wire         accessDataValid_pipe_pipe_out_29_valid = accessDataValid_pipe_pipe_v_29;
  wire         accessDataSource_29_valid = accessDataValid_pipe_pipe_out_29_valid;
  reg          shifterReg_45_0_valid;
  reg  [31:0]  shifterReg_45_0_bits;
  wire         shifterValid_45 = shifterReg_45_0_valid | accessDataSource_29_valid;
  wire         sinkVec_tokenCheck_58;
  wire [4:0]   sinkVec_validSource_58_bits_vd = x22_14_0_bits_vd;
  wire [1:0]   sinkVec_validSource_58_bits_offset = x22_14_0_bits_offset;
  wire [3:0]   sinkVec_validSource_58_bits_mask = x22_14_0_bits_mask;
  wire [31:0]  sinkVec_validSource_58_bits_data = x22_14_0_bits_data;
  wire [2:0]   sinkVec_validSource_58_bits_instructionIndex = x22_14_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_59;
  wire [4:0]   sinkVec_validSource_59_bits_vd = x22_14_1_bits_vd;
  wire [1:0]   sinkVec_validSource_59_bits_offset = x22_14_1_bits_offset;
  wire [3:0]   sinkVec_validSource_59_bits_mask = x22_14_1_bits_mask;
  wire [31:0]  sinkVec_validSource_59_bits_data = x22_14_1_bits_data;
  wire         sinkVec_validSource_59_bits_last = x22_14_1_bits_last;
  wire [2:0]   sinkVec_validSource_59_bits_instructionIndex = x22_14_1_bits_instructionIndex;
  wire         sinkVec_29_0_ready;
  wire         sinkVec_queue_58_deq_ready = sinkVec_sinkWire_58_ready;
  wire         sinkVec_queue_58_deq_valid;
  wire [4:0]   sinkVec_queue_58_deq_bits_vd;
  wire         sinkVec_29_0_valid = sinkVec_sinkWire_58_valid;
  wire [1:0]   sinkVec_queue_58_deq_bits_offset;
  wire [4:0]   sinkVec_29_0_bits_vd = sinkVec_sinkWire_58_bits_vd;
  wire [3:0]   sinkVec_queue_58_deq_bits_mask;
  wire [1:0]   sinkVec_29_0_bits_offset = sinkVec_sinkWire_58_bits_offset;
  wire [31:0]  sinkVec_queue_58_deq_bits_data;
  wire [3:0]   sinkVec_29_0_bits_mask = sinkVec_sinkWire_58_bits_mask;
  wire         sinkVec_queue_58_deq_bits_last;
  wire [31:0]  sinkVec_29_0_bits_data = sinkVec_sinkWire_58_bits_data;
  wire [2:0]   sinkVec_queue_58_deq_bits_instructionIndex;
  wire         sinkVec_29_0_bits_last = sinkVec_sinkWire_58_bits_last;
  wire [2:0]   sinkVec_29_0_bits_instructionIndex = sinkVec_sinkWire_58_bits_instructionIndex;
  wire         sinkVec_validSink_58_valid;
  wire [4:0]   sinkVec_validSink_58_bits_vd;
  wire [1:0]   sinkVec_validSink_58_bits_offset;
  wire [3:0]   sinkVec_validSink_58_bits_mask;
  wire [31:0]  sinkVec_validSink_58_bits_data;
  wire [2:0]   sinkVec_validSink_58_bits_instructionIndex;
  assign sinkVec_sinkWire_58_valid = sinkVec_queue_58_deq_valid;
  assign sinkVec_sinkWire_58_bits_vd = sinkVec_queue_58_deq_bits_vd;
  assign sinkVec_sinkWire_58_bits_offset = sinkVec_queue_58_deq_bits_offset;
  assign sinkVec_sinkWire_58_bits_mask = sinkVec_queue_58_deq_bits_mask;
  assign sinkVec_sinkWire_58_bits_data = sinkVec_queue_58_deq_bits_data;
  assign sinkVec_sinkWire_58_bits_last = sinkVec_queue_58_deq_bits_last;
  assign sinkVec_sinkWire_58_bits_instructionIndex = sinkVec_queue_58_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_58_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_28 = {sinkVec_queue_58_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_58_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_58 = {sinkVec_queue_dataIn_lo_hi_28, sinkVec_queue_58_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_58_enq_bits_vd;
  wire [1:0]   sinkVec_queue_58_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_28 = {sinkVec_queue_58_enq_bits_vd, sinkVec_queue_58_enq_bits_offset};
  wire [3:0]   sinkVec_queue_58_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_58 = {sinkVec_queue_dataIn_hi_hi_28, sinkVec_queue_58_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_58 = {sinkVec_queue_dataIn_hi_58, sinkVec_queue_dataIn_lo_58};
  wire [2:0]   sinkVec_queue_dataOut_58_instructionIndex = _sinkVec_queue_fifo_58_data_out[2:0];
  wire         sinkVec_queue_dataOut_58_last = _sinkVec_queue_fifo_58_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_58_data = _sinkVec_queue_fifo_58_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_58_mask = _sinkVec_queue_fifo_58_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_58_offset = _sinkVec_queue_fifo_58_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_58_vd = _sinkVec_queue_fifo_58_data_out[46:42];
  wire         sinkVec_queue_58_enq_ready = ~_sinkVec_queue_fifo_58_full;
  wire         sinkVec_queue_58_enq_valid;
  assign sinkVec_queue_58_deq_valid = ~_sinkVec_queue_fifo_58_empty | sinkVec_queue_58_enq_valid;
  assign sinkVec_queue_58_deq_bits_vd = _sinkVec_queue_fifo_58_empty ? sinkVec_queue_58_enq_bits_vd : sinkVec_queue_dataOut_58_vd;
  assign sinkVec_queue_58_deq_bits_offset = _sinkVec_queue_fifo_58_empty ? sinkVec_queue_58_enq_bits_offset : sinkVec_queue_dataOut_58_offset;
  assign sinkVec_queue_58_deq_bits_mask = _sinkVec_queue_fifo_58_empty ? sinkVec_queue_58_enq_bits_mask : sinkVec_queue_dataOut_58_mask;
  assign sinkVec_queue_58_deq_bits_data = _sinkVec_queue_fifo_58_empty ? sinkVec_queue_58_enq_bits_data : sinkVec_queue_dataOut_58_data;
  assign sinkVec_queue_58_deq_bits_last = ~_sinkVec_queue_fifo_58_empty & sinkVec_queue_dataOut_58_last;
  assign sinkVec_queue_58_deq_bits_instructionIndex = _sinkVec_queue_fifo_58_empty ? sinkVec_queue_58_enq_bits_instructionIndex : sinkVec_queue_dataOut_58_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_58;
  wire         sinkVec_releasePipe_pipe_out_58_valid = sinkVec_releasePipe_pipe_v_58;
  wire         x22_14_0_ready;
  wire         x22_14_0_valid;
  wire         sinkVec_validSource_58_valid = x22_14_0_ready & x22_14_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_58;
  wire [2:0]   sinkVec_tokenCheck_counterChange_58 = sinkVec_validSource_58_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_58 = ~(sinkVec_tokenCheck_counter_58[2]);
  assign x22_14_0_ready = sinkVec_tokenCheck_58;
  assign sinkVec_queue_58_enq_valid = sinkVec_validSink_58_valid;
  assign sinkVec_queue_58_enq_bits_vd = sinkVec_validSink_58_bits_vd;
  assign sinkVec_queue_58_enq_bits_offset = sinkVec_validSink_58_bits_offset;
  assign sinkVec_queue_58_enq_bits_mask = sinkVec_validSink_58_bits_mask;
  assign sinkVec_queue_58_enq_bits_data = sinkVec_validSink_58_bits_data;
  assign sinkVec_queue_58_enq_bits_instructionIndex = sinkVec_validSink_58_bits_instructionIndex;
  reg          sinkVec_shifterReg_58_0_valid;
  assign sinkVec_validSink_58_valid = sinkVec_shifterReg_58_0_valid;
  reg  [4:0]   sinkVec_shifterReg_58_0_bits_vd;
  assign sinkVec_validSink_58_bits_vd = sinkVec_shifterReg_58_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_58_0_bits_offset;
  assign sinkVec_validSink_58_bits_offset = sinkVec_shifterReg_58_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_58_0_bits_mask;
  assign sinkVec_validSink_58_bits_mask = sinkVec_shifterReg_58_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_58_0_bits_data;
  assign sinkVec_validSink_58_bits_data = sinkVec_shifterReg_58_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_58_0_bits_instructionIndex;
  assign sinkVec_validSink_58_bits_instructionIndex = sinkVec_shifterReg_58_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_58 = sinkVec_shifterReg_58_0_valid | sinkVec_validSource_58_valid;
  wire         sinkVec_29_1_ready;
  wire         sinkVec_queue_59_deq_ready = sinkVec_sinkWire_59_ready;
  wire         sinkVec_queue_59_deq_valid;
  wire [4:0]   sinkVec_queue_59_deq_bits_vd;
  wire         sinkVec_29_1_valid = sinkVec_sinkWire_59_valid;
  wire [1:0]   sinkVec_queue_59_deq_bits_offset;
  wire [4:0]   sinkVec_29_1_bits_vd = sinkVec_sinkWire_59_bits_vd;
  wire [3:0]   sinkVec_queue_59_deq_bits_mask;
  wire [1:0]   sinkVec_29_1_bits_offset = sinkVec_sinkWire_59_bits_offset;
  wire [31:0]  sinkVec_queue_59_deq_bits_data;
  wire [3:0]   sinkVec_29_1_bits_mask = sinkVec_sinkWire_59_bits_mask;
  wire         sinkVec_queue_59_deq_bits_last;
  wire [31:0]  sinkVec_29_1_bits_data = sinkVec_sinkWire_59_bits_data;
  wire [2:0]   sinkVec_queue_59_deq_bits_instructionIndex;
  wire         sinkVec_29_1_bits_last = sinkVec_sinkWire_59_bits_last;
  wire [2:0]   sinkVec_29_1_bits_instructionIndex = sinkVec_sinkWire_59_bits_instructionIndex;
  wire         sinkVec_validSink_59_valid;
  wire [4:0]   sinkVec_validSink_59_bits_vd;
  wire [1:0]   sinkVec_validSink_59_bits_offset;
  wire [3:0]   sinkVec_validSink_59_bits_mask;
  wire [31:0]  sinkVec_validSink_59_bits_data;
  wire         sinkVec_validSink_59_bits_last;
  wire [2:0]   sinkVec_validSink_59_bits_instructionIndex;
  assign sinkVec_sinkWire_59_valid = sinkVec_queue_59_deq_valid;
  assign sinkVec_sinkWire_59_bits_vd = sinkVec_queue_59_deq_bits_vd;
  assign sinkVec_sinkWire_59_bits_offset = sinkVec_queue_59_deq_bits_offset;
  assign sinkVec_sinkWire_59_bits_mask = sinkVec_queue_59_deq_bits_mask;
  assign sinkVec_sinkWire_59_bits_data = sinkVec_queue_59_deq_bits_data;
  assign sinkVec_sinkWire_59_bits_last = sinkVec_queue_59_deq_bits_last;
  assign sinkVec_sinkWire_59_bits_instructionIndex = sinkVec_queue_59_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_59_enq_bits_data;
  wire         sinkVec_queue_59_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_29 = {sinkVec_queue_59_enq_bits_data, sinkVec_queue_59_enq_bits_last};
  wire [2:0]   sinkVec_queue_59_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_59 = {sinkVec_queue_dataIn_lo_hi_29, sinkVec_queue_59_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_59_enq_bits_vd;
  wire [1:0]   sinkVec_queue_59_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_29 = {sinkVec_queue_59_enq_bits_vd, sinkVec_queue_59_enq_bits_offset};
  wire [3:0]   sinkVec_queue_59_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_59 = {sinkVec_queue_dataIn_hi_hi_29, sinkVec_queue_59_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_59 = {sinkVec_queue_dataIn_hi_59, sinkVec_queue_dataIn_lo_59};
  wire [2:0]   sinkVec_queue_dataOut_59_instructionIndex = _sinkVec_queue_fifo_59_data_out[2:0];
  wire         sinkVec_queue_dataOut_59_last = _sinkVec_queue_fifo_59_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_59_data = _sinkVec_queue_fifo_59_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_59_mask = _sinkVec_queue_fifo_59_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_59_offset = _sinkVec_queue_fifo_59_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_59_vd = _sinkVec_queue_fifo_59_data_out[46:42];
  wire         sinkVec_queue_59_enq_ready = ~_sinkVec_queue_fifo_59_full;
  wire         sinkVec_queue_59_enq_valid;
  assign sinkVec_queue_59_deq_valid = ~_sinkVec_queue_fifo_59_empty | sinkVec_queue_59_enq_valid;
  assign sinkVec_queue_59_deq_bits_vd = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_vd : sinkVec_queue_dataOut_59_vd;
  assign sinkVec_queue_59_deq_bits_offset = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_offset : sinkVec_queue_dataOut_59_offset;
  assign sinkVec_queue_59_deq_bits_mask = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_mask : sinkVec_queue_dataOut_59_mask;
  assign sinkVec_queue_59_deq_bits_data = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_data : sinkVec_queue_dataOut_59_data;
  assign sinkVec_queue_59_deq_bits_last = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_last : sinkVec_queue_dataOut_59_last;
  assign sinkVec_queue_59_deq_bits_instructionIndex = _sinkVec_queue_fifo_59_empty ? sinkVec_queue_59_enq_bits_instructionIndex : sinkVec_queue_dataOut_59_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_59;
  wire         sinkVec_releasePipe_pipe_out_59_valid = sinkVec_releasePipe_pipe_v_59;
  wire         x22_14_1_ready;
  wire         x22_14_1_valid;
  wire         sinkVec_validSource_59_valid = x22_14_1_ready & x22_14_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_59;
  wire [2:0]   sinkVec_tokenCheck_counterChange_59 = sinkVec_validSource_59_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_59 = ~(sinkVec_tokenCheck_counter_59[2]);
  assign x22_14_1_ready = sinkVec_tokenCheck_59;
  assign sinkVec_queue_59_enq_valid = sinkVec_validSink_59_valid;
  assign sinkVec_queue_59_enq_bits_vd = sinkVec_validSink_59_bits_vd;
  assign sinkVec_queue_59_enq_bits_offset = sinkVec_validSink_59_bits_offset;
  assign sinkVec_queue_59_enq_bits_mask = sinkVec_validSink_59_bits_mask;
  assign sinkVec_queue_59_enq_bits_data = sinkVec_validSink_59_bits_data;
  assign sinkVec_queue_59_enq_bits_last = sinkVec_validSink_59_bits_last;
  assign sinkVec_queue_59_enq_bits_instructionIndex = sinkVec_validSink_59_bits_instructionIndex;
  reg          sinkVec_shifterReg_59_0_valid;
  assign sinkVec_validSink_59_valid = sinkVec_shifterReg_59_0_valid;
  reg  [4:0]   sinkVec_shifterReg_59_0_bits_vd;
  assign sinkVec_validSink_59_bits_vd = sinkVec_shifterReg_59_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_59_0_bits_offset;
  assign sinkVec_validSink_59_bits_offset = sinkVec_shifterReg_59_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_59_0_bits_mask;
  assign sinkVec_validSink_59_bits_mask = sinkVec_shifterReg_59_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_59_0_bits_data;
  assign sinkVec_validSink_59_bits_data = sinkVec_shifterReg_59_0_bits_data;
  reg          sinkVec_shifterReg_59_0_bits_last;
  assign sinkVec_validSink_59_bits_last = sinkVec_shifterReg_59_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_59_0_bits_instructionIndex;
  assign sinkVec_validSink_59_bits_instructionIndex = sinkVec_shifterReg_59_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_59 = sinkVec_shifterReg_59_0_valid | sinkVec_validSource_59_valid;
  assign sinkVec_sinkWire_58_ready = sinkVec_29_0_ready;
  assign sinkVec_sinkWire_59_ready = sinkVec_29_1_ready;
  reg          maskUnitFirst_29;
  wire         tryToRead_29 = sinkVec_29_0_valid | sinkVec_29_1_valid;
  wire         sinkWire_29_valid = maskUnitFirst_29 ? sinkVec_29_0_valid : sinkVec_29_1_valid;
  wire [4:0]   sinkWire_29_bits_vd = maskUnitFirst_29 ? sinkVec_29_0_bits_vd : sinkVec_29_1_bits_vd;
  wire [1:0]   sinkWire_29_bits_offset = maskUnitFirst_29 ? sinkVec_29_0_bits_offset : sinkVec_29_1_bits_offset;
  wire [3:0]   sinkWire_29_bits_mask = maskUnitFirst_29 ? sinkVec_29_0_bits_mask : sinkVec_29_1_bits_mask;
  wire [31:0]  sinkWire_29_bits_data = maskUnitFirst_29 ? sinkVec_29_0_bits_data : sinkVec_29_1_bits_data;
  wire         sinkWire_29_bits_last = maskUnitFirst_29 ? sinkVec_29_0_bits_last : sinkVec_29_1_bits_last;
  wire [2:0]   sinkWire_29_bits_instructionIndex = maskUnitFirst_29 ? sinkVec_29_0_bits_instructionIndex : sinkVec_29_1_bits_instructionIndex;
  wire         sinkWire_29_ready;
  assign sinkVec_29_1_ready = sinkWire_29_ready & ~maskUnitFirst_29;
  assign sinkVec_29_0_ready = sinkWire_29_ready & maskUnitFirst_29;
  reg          view__writeRelease_14_pipe_v;
  wire         view__writeRelease_14_pipe_out_valid = view__writeRelease_14_pipe_v;
  reg          pipe_v_42;
  wire         pipe_out_28_valid = pipe_v_42;
  wire         _probeWire_writeQueueEnqVec_14_valid_T = x22_14_0_ready & _maskUnit_exeResp_14_valid;
  reg          instructionFinishedPipe_pipe_v_14;
  wire         instructionFinishedPipe_pipe_out_14_valid = instructionFinishedPipe_pipe_v_14;
  reg  [7:0]   instructionFinishedPipe_pipe_b_14;
  wire [7:0]   instructionFinishedPipe_pipe_out_14_bits = instructionFinishedPipe_pipe_b_14;
  wire         instructionFinished_14_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_14_bits);
  wire         instructionFinished_14_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_14_bits);
  wire         instructionFinished_14_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_14_bits);
  wire         instructionFinished_14_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_14_bits);
  assign vxsatReportVec_14 = _laneVec_14_vxsatReport[3:0];
  reg          pipe_v_43;
  reg  [31:0]  pipe_b_43;
  reg          pipe_pipe_v_14;
  wire         pipe_pipe_out_14_valid = pipe_pipe_v_14;
  reg  [31:0]  pipe_pipe_b_14;
  wire [31:0]  pipe_pipe_out_14_bits = pipe_pipe_b_14;
  reg          view__laneMaskSelect_14_pipe_v;
  reg  [5:0]   view__laneMaskSelect_14_pipe_b;
  reg          view__laneMaskSelect_14_pipe_pipe_v;
  wire         view__laneMaskSelect_14_pipe_pipe_out_valid = view__laneMaskSelect_14_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_14_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_14_pipe_pipe_out_bits = view__laneMaskSelect_14_pipe_pipe_b;
  reg          view__laneMaskSewSelect_14_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_14_pipe_b;
  reg          view__laneMaskSewSelect_14_pipe_pipe_v;
  wire         view__laneMaskSewSelect_14_pipe_pipe_out_valid = view__laneMaskSewSelect_14_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_14_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_14_pipe_pipe_out_bits = view__laneMaskSewSelect_14_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_14;
  wire         lsuLastPipe_pipe_out_14_valid = lsuLastPipe_pipe_v_14;
  reg  [7:0]   lsuLastPipe_pipe_b_14;
  wire [7:0]   lsuLastPipe_pipe_out_14_bits = lsuLastPipe_pipe_b_14;
  reg          maskLastPipe_pipe_v_14;
  wire         maskLastPipe_pipe_out_14_valid = maskLastPipe_pipe_v_14;
  reg  [7:0]   maskLastPipe_pipe_b_14;
  wire [7:0]   maskLastPipe_pipe_out_14_bits = maskLastPipe_pipe_b_14;
  wire [5:0]   writeCounter_14 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h38};
  reg          pipe_v_44;
  wire         pipe_out_29_valid = pipe_v_44;
  reg  [5:0]   pipe_b_44;
  wire [5:0]   pipe_out_29_bits = pipe_b_44;
  assign laneRequestSinkWire_15_ready = ~laneRequestSinkWire_15_bits_issueInst | _laneVec_15_laneRequest_ready;
  wire         sinkVec_tokenCheck_60;
  wire [4:0]   sinkVec_validSource_60_bits_vs = x13_15_0_bits_vs;
  wire [1:0]   sinkVec_validSource_60_bits_offset = x13_15_0_bits_offset;
  wire [2:0]   sinkVec_validSource_60_bits_instructionIndex = x13_15_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_61;
  wire [4:0]   sinkVec_validSource_61_bits_vs = x13_15_1_bits_vs;
  wire [1:0]   sinkVec_validSource_61_bits_offset = x13_15_1_bits_offset;
  wire [2:0]   sinkVec_validSource_61_bits_instructionIndex = x13_15_1_bits_instructionIndex;
  wire         sinkVec_30_0_ready;
  wire         sinkVec_queue_60_deq_ready = sinkVec_sinkWire_60_ready;
  wire         sinkVec_queue_60_deq_valid;
  wire [4:0]   sinkVec_queue_60_deq_bits_vs;
  wire         sinkVec_30_0_valid = sinkVec_sinkWire_60_valid;
  wire [1:0]   sinkVec_queue_60_deq_bits_readSource;
  wire [4:0]   sinkVec_30_0_bits_vs = sinkVec_sinkWire_60_bits_vs;
  wire [1:0]   sinkVec_queue_60_deq_bits_offset;
  wire [1:0]   sinkVec_30_0_bits_readSource = sinkVec_sinkWire_60_bits_readSource;
  wire [2:0]   sinkVec_queue_60_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_30_0_bits_offset = sinkVec_sinkWire_60_bits_offset;
  wire [2:0]   sinkVec_30_0_bits_instructionIndex = sinkVec_sinkWire_60_bits_instructionIndex;
  wire         sinkVec_validSink_60_valid;
  wire [4:0]   sinkVec_validSink_60_bits_vs;
  wire [1:0]   sinkVec_validSink_60_bits_readSource;
  wire [1:0]   sinkVec_validSink_60_bits_offset;
  wire [2:0]   sinkVec_validSink_60_bits_instructionIndex;
  assign sinkVec_sinkWire_60_valid = sinkVec_queue_60_deq_valid;
  assign sinkVec_sinkWire_60_bits_vs = sinkVec_queue_60_deq_bits_vs;
  assign sinkVec_sinkWire_60_bits_readSource = sinkVec_queue_60_deq_bits_readSource;
  assign sinkVec_sinkWire_60_bits_offset = sinkVec_queue_60_deq_bits_offset;
  assign sinkVec_sinkWire_60_bits_instructionIndex = sinkVec_queue_60_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_60_enq_bits_offset;
  wire [2:0]   sinkVec_queue_60_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_60 = {sinkVec_queue_60_enq_bits_offset, sinkVec_queue_60_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_60_enq_bits_vs;
  wire [1:0]   sinkVec_queue_60_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_60 = {sinkVec_queue_60_enq_bits_vs, sinkVec_queue_60_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_60 = {sinkVec_queue_dataIn_hi_60, sinkVec_queue_dataIn_lo_60};
  wire [2:0]   sinkVec_queue_dataOut_60_instructionIndex = _sinkVec_queue_fifo_60_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_60_offset = _sinkVec_queue_fifo_60_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_60_readSource = _sinkVec_queue_fifo_60_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_60_vs = _sinkVec_queue_fifo_60_data_out[11:7];
  wire         sinkVec_queue_60_enq_ready = ~_sinkVec_queue_fifo_60_full;
  wire         sinkVec_queue_60_enq_valid;
  assign sinkVec_queue_60_deq_valid = ~_sinkVec_queue_fifo_60_empty | sinkVec_queue_60_enq_valid;
  assign sinkVec_queue_60_deq_bits_vs = _sinkVec_queue_fifo_60_empty ? sinkVec_queue_60_enq_bits_vs : sinkVec_queue_dataOut_60_vs;
  assign sinkVec_queue_60_deq_bits_readSource = _sinkVec_queue_fifo_60_empty ? sinkVec_queue_60_enq_bits_readSource : sinkVec_queue_dataOut_60_readSource;
  assign sinkVec_queue_60_deq_bits_offset = _sinkVec_queue_fifo_60_empty ? sinkVec_queue_60_enq_bits_offset : sinkVec_queue_dataOut_60_offset;
  assign sinkVec_queue_60_deq_bits_instructionIndex = _sinkVec_queue_fifo_60_empty ? sinkVec_queue_60_enq_bits_instructionIndex : sinkVec_queue_dataOut_60_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_60;
  wire         sinkVec_releasePipe_pipe_out_60_valid = sinkVec_releasePipe_pipe_v_60;
  wire         x13_15_0_ready;
  wire         x13_15_0_valid;
  wire         sinkVec_validSource_60_valid = x13_15_0_ready & x13_15_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_60;
  wire [2:0]   sinkVec_tokenCheck_counterChange_60 = sinkVec_validSource_60_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_60 = ~(sinkVec_tokenCheck_counter_60[2]);
  assign x13_15_0_ready = sinkVec_tokenCheck_60;
  assign sinkVec_queue_60_enq_valid = sinkVec_validSink_60_valid;
  assign sinkVec_queue_60_enq_bits_vs = sinkVec_validSink_60_bits_vs;
  assign sinkVec_queue_60_enq_bits_readSource = sinkVec_validSink_60_bits_readSource;
  assign sinkVec_queue_60_enq_bits_offset = sinkVec_validSink_60_bits_offset;
  assign sinkVec_queue_60_enq_bits_instructionIndex = sinkVec_validSink_60_bits_instructionIndex;
  reg          sinkVec_shifterReg_60_0_valid;
  assign sinkVec_validSink_60_valid = sinkVec_shifterReg_60_0_valid;
  reg  [4:0]   sinkVec_shifterReg_60_0_bits_vs;
  assign sinkVec_validSink_60_bits_vs = sinkVec_shifterReg_60_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_60_0_bits_readSource;
  assign sinkVec_validSink_60_bits_readSource = sinkVec_shifterReg_60_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_60_0_bits_offset;
  assign sinkVec_validSink_60_bits_offset = sinkVec_shifterReg_60_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_60_0_bits_instructionIndex;
  assign sinkVec_validSink_60_bits_instructionIndex = sinkVec_shifterReg_60_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_60 = sinkVec_shifterReg_60_0_valid | sinkVec_validSource_60_valid;
  wire         sinkVec_30_1_ready;
  wire         sinkVec_queue_61_deq_ready = sinkVec_sinkWire_61_ready;
  wire         sinkVec_queue_61_deq_valid;
  wire [4:0]   sinkVec_queue_61_deq_bits_vs;
  wire         sinkVec_30_1_valid = sinkVec_sinkWire_61_valid;
  wire [1:0]   sinkVec_queue_61_deq_bits_readSource;
  wire [4:0]   sinkVec_30_1_bits_vs = sinkVec_sinkWire_61_bits_vs;
  wire [1:0]   sinkVec_queue_61_deq_bits_offset;
  wire [1:0]   sinkVec_30_1_bits_readSource = sinkVec_sinkWire_61_bits_readSource;
  wire [2:0]   sinkVec_queue_61_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_30_1_bits_offset = sinkVec_sinkWire_61_bits_offset;
  wire [2:0]   sinkVec_30_1_bits_instructionIndex = sinkVec_sinkWire_61_bits_instructionIndex;
  wire         sinkVec_validSink_61_valid;
  wire [4:0]   sinkVec_validSink_61_bits_vs;
  wire [1:0]   sinkVec_validSink_61_bits_readSource;
  wire [1:0]   sinkVec_validSink_61_bits_offset;
  wire [2:0]   sinkVec_validSink_61_bits_instructionIndex;
  assign sinkVec_sinkWire_61_valid = sinkVec_queue_61_deq_valid;
  assign sinkVec_sinkWire_61_bits_vs = sinkVec_queue_61_deq_bits_vs;
  assign sinkVec_sinkWire_61_bits_readSource = sinkVec_queue_61_deq_bits_readSource;
  assign sinkVec_sinkWire_61_bits_offset = sinkVec_queue_61_deq_bits_offset;
  assign sinkVec_sinkWire_61_bits_instructionIndex = sinkVec_queue_61_deq_bits_instructionIndex;
  wire [1:0]   sinkVec_queue_61_enq_bits_offset;
  wire [2:0]   sinkVec_queue_61_enq_bits_instructionIndex;
  wire [4:0]   sinkVec_queue_dataIn_lo_61 = {sinkVec_queue_61_enq_bits_offset, sinkVec_queue_61_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_61_enq_bits_vs;
  wire [1:0]   sinkVec_queue_61_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_61 = {sinkVec_queue_61_enq_bits_vs, sinkVec_queue_61_enq_bits_readSource};
  wire [11:0]  sinkVec_queue_dataIn_61 = {sinkVec_queue_dataIn_hi_61, sinkVec_queue_dataIn_lo_61};
  wire [2:0]   sinkVec_queue_dataOut_61_instructionIndex = _sinkVec_queue_fifo_61_data_out[2:0];
  wire [1:0]   sinkVec_queue_dataOut_61_offset = _sinkVec_queue_fifo_61_data_out[4:3];
  wire [1:0]   sinkVec_queue_dataOut_61_readSource = _sinkVec_queue_fifo_61_data_out[6:5];
  wire [4:0]   sinkVec_queue_dataOut_61_vs = _sinkVec_queue_fifo_61_data_out[11:7];
  wire         sinkVec_queue_61_enq_ready = ~_sinkVec_queue_fifo_61_full;
  wire         sinkVec_queue_61_enq_valid;
  assign sinkVec_queue_61_deq_valid = ~_sinkVec_queue_fifo_61_empty | sinkVec_queue_61_enq_valid;
  assign sinkVec_queue_61_deq_bits_vs = _sinkVec_queue_fifo_61_empty ? sinkVec_queue_61_enq_bits_vs : sinkVec_queue_dataOut_61_vs;
  assign sinkVec_queue_61_deq_bits_readSource = _sinkVec_queue_fifo_61_empty ? sinkVec_queue_61_enq_bits_readSource : sinkVec_queue_dataOut_61_readSource;
  assign sinkVec_queue_61_deq_bits_offset = _sinkVec_queue_fifo_61_empty ? sinkVec_queue_61_enq_bits_offset : sinkVec_queue_dataOut_61_offset;
  assign sinkVec_queue_61_deq_bits_instructionIndex = _sinkVec_queue_fifo_61_empty ? sinkVec_queue_61_enq_bits_instructionIndex : sinkVec_queue_dataOut_61_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_61;
  wire         sinkVec_releasePipe_pipe_out_61_valid = sinkVec_releasePipe_pipe_v_61;
  wire         x13_15_1_ready;
  wire         x13_15_1_valid;
  wire         sinkVec_validSource_61_valid = x13_15_1_ready & x13_15_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_61;
  wire [2:0]   sinkVec_tokenCheck_counterChange_61 = sinkVec_validSource_61_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_61 = ~(sinkVec_tokenCheck_counter_61[2]);
  assign x13_15_1_ready = sinkVec_tokenCheck_61;
  assign sinkVec_queue_61_enq_valid = sinkVec_validSink_61_valid;
  assign sinkVec_queue_61_enq_bits_vs = sinkVec_validSink_61_bits_vs;
  assign sinkVec_queue_61_enq_bits_readSource = sinkVec_validSink_61_bits_readSource;
  assign sinkVec_queue_61_enq_bits_offset = sinkVec_validSink_61_bits_offset;
  assign sinkVec_queue_61_enq_bits_instructionIndex = sinkVec_validSink_61_bits_instructionIndex;
  reg          sinkVec_shifterReg_61_0_valid;
  assign sinkVec_validSink_61_valid = sinkVec_shifterReg_61_0_valid;
  reg  [4:0]   sinkVec_shifterReg_61_0_bits_vs;
  assign sinkVec_validSink_61_bits_vs = sinkVec_shifterReg_61_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_61_0_bits_readSource;
  assign sinkVec_validSink_61_bits_readSource = sinkVec_shifterReg_61_0_bits_readSource;
  reg  [1:0]   sinkVec_shifterReg_61_0_bits_offset;
  assign sinkVec_validSink_61_bits_offset = sinkVec_shifterReg_61_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_61_0_bits_instructionIndex;
  assign sinkVec_validSink_61_bits_instructionIndex = sinkVec_shifterReg_61_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_61 = sinkVec_shifterReg_61_0_valid | sinkVec_validSource_61_valid;
  assign sinkVec_sinkWire_60_ready = sinkVec_30_0_ready;
  assign sinkVec_sinkWire_61_ready = sinkVec_30_1_ready;
  reg          maskUnitFirst_30;
  wire         tryToRead_30 = sinkVec_30_0_valid | sinkVec_30_1_valid;
  wire         sinkWire_30_valid = maskUnitFirst_30 ? sinkVec_30_0_valid : sinkVec_30_1_valid;
  wire [4:0]   sinkWire_30_bits_vs = maskUnitFirst_30 ? sinkVec_30_0_bits_vs : sinkVec_30_1_bits_vs;
  wire [1:0]   sinkWire_30_bits_readSource = maskUnitFirst_30 ? sinkVec_30_0_bits_readSource : sinkVec_30_1_bits_readSource;
  wire [1:0]   sinkWire_30_bits_offset = maskUnitFirst_30 ? sinkVec_30_0_bits_offset : sinkVec_30_1_bits_offset;
  wire [2:0]   sinkWire_30_bits_instructionIndex = maskUnitFirst_30 ? sinkVec_30_0_bits_instructionIndex : sinkVec_30_1_bits_instructionIndex;
  wire         sinkWire_30_ready;
  assign sinkVec_30_1_ready = sinkWire_30_ready & ~maskUnitFirst_30;
  assign sinkVec_30_0_ready = sinkWire_30_ready & maskUnitFirst_30;
  reg          accessDataValid_pipe_v_30;
  reg          accessDataValid_pipe_pipe_v_30;
  wire         accessDataValid_pipe_pipe_out_30_valid = accessDataValid_pipe_pipe_v_30;
  wire         accessDataSource_30_valid = accessDataValid_pipe_pipe_out_30_valid;
  reg          shifterReg_46_0_valid;
  reg  [31:0]  shifterReg_46_0_bits;
  wire         shifterValid_46 = shifterReg_46_0_valid | accessDataSource_30_valid;
  reg          accessDataValid_pipe_v_31;
  reg          accessDataValid_pipe_pipe_v_31;
  wire         accessDataValid_pipe_pipe_out_31_valid = accessDataValid_pipe_pipe_v_31;
  wire         accessDataSource_31_valid = accessDataValid_pipe_pipe_out_31_valid;
  reg          shifterReg_47_0_valid;
  reg  [31:0]  shifterReg_47_0_bits;
  wire         shifterValid_47 = shifterReg_47_0_valid | accessDataSource_31_valid;
  wire         sinkVec_tokenCheck_62;
  wire [4:0]   sinkVec_validSource_62_bits_vd = x22_15_0_bits_vd;
  wire [1:0]   sinkVec_validSource_62_bits_offset = x22_15_0_bits_offset;
  wire [3:0]   sinkVec_validSource_62_bits_mask = x22_15_0_bits_mask;
  wire [31:0]  sinkVec_validSource_62_bits_data = x22_15_0_bits_data;
  wire [2:0]   sinkVec_validSource_62_bits_instructionIndex = x22_15_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_63;
  wire [4:0]   sinkVec_validSource_63_bits_vd = x22_15_1_bits_vd;
  wire [1:0]   sinkVec_validSource_63_bits_offset = x22_15_1_bits_offset;
  wire [3:0]   sinkVec_validSource_63_bits_mask = x22_15_1_bits_mask;
  wire [31:0]  sinkVec_validSource_63_bits_data = x22_15_1_bits_data;
  wire         sinkVec_validSource_63_bits_last = x22_15_1_bits_last;
  wire [2:0]   sinkVec_validSource_63_bits_instructionIndex = x22_15_1_bits_instructionIndex;
  wire         sinkVec_31_0_ready;
  wire         sinkVec_queue_62_deq_ready = sinkVec_sinkWire_62_ready;
  wire         sinkVec_queue_62_deq_valid;
  wire [4:0]   sinkVec_queue_62_deq_bits_vd;
  wire         sinkVec_31_0_valid = sinkVec_sinkWire_62_valid;
  wire [1:0]   sinkVec_queue_62_deq_bits_offset;
  wire [4:0]   sinkVec_31_0_bits_vd = sinkVec_sinkWire_62_bits_vd;
  wire [3:0]   sinkVec_queue_62_deq_bits_mask;
  wire [1:0]   sinkVec_31_0_bits_offset = sinkVec_sinkWire_62_bits_offset;
  wire [31:0]  sinkVec_queue_62_deq_bits_data;
  wire [3:0]   sinkVec_31_0_bits_mask = sinkVec_sinkWire_62_bits_mask;
  wire         sinkVec_queue_62_deq_bits_last;
  wire [31:0]  sinkVec_31_0_bits_data = sinkVec_sinkWire_62_bits_data;
  wire [2:0]   sinkVec_queue_62_deq_bits_instructionIndex;
  wire         sinkVec_31_0_bits_last = sinkVec_sinkWire_62_bits_last;
  wire [2:0]   sinkVec_31_0_bits_instructionIndex = sinkVec_sinkWire_62_bits_instructionIndex;
  wire         sinkVec_validSink_62_valid;
  wire [4:0]   sinkVec_validSink_62_bits_vd;
  wire [1:0]   sinkVec_validSink_62_bits_offset;
  wire [3:0]   sinkVec_validSink_62_bits_mask;
  wire [31:0]  sinkVec_validSink_62_bits_data;
  wire [2:0]   sinkVec_validSink_62_bits_instructionIndex;
  assign sinkVec_sinkWire_62_valid = sinkVec_queue_62_deq_valid;
  assign sinkVec_sinkWire_62_bits_vd = sinkVec_queue_62_deq_bits_vd;
  assign sinkVec_sinkWire_62_bits_offset = sinkVec_queue_62_deq_bits_offset;
  assign sinkVec_sinkWire_62_bits_mask = sinkVec_queue_62_deq_bits_mask;
  assign sinkVec_sinkWire_62_bits_data = sinkVec_queue_62_deq_bits_data;
  assign sinkVec_sinkWire_62_bits_last = sinkVec_queue_62_deq_bits_last;
  assign sinkVec_sinkWire_62_bits_instructionIndex = sinkVec_queue_62_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_62_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_30 = {sinkVec_queue_62_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_62_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_62 = {sinkVec_queue_dataIn_lo_hi_30, sinkVec_queue_62_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_62_enq_bits_vd;
  wire [1:0]   sinkVec_queue_62_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_30 = {sinkVec_queue_62_enq_bits_vd, sinkVec_queue_62_enq_bits_offset};
  wire [3:0]   sinkVec_queue_62_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_62 = {sinkVec_queue_dataIn_hi_hi_30, sinkVec_queue_62_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_62 = {sinkVec_queue_dataIn_hi_62, sinkVec_queue_dataIn_lo_62};
  wire [2:0]   sinkVec_queue_dataOut_62_instructionIndex = _sinkVec_queue_fifo_62_data_out[2:0];
  wire         sinkVec_queue_dataOut_62_last = _sinkVec_queue_fifo_62_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_62_data = _sinkVec_queue_fifo_62_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_62_mask = _sinkVec_queue_fifo_62_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_62_offset = _sinkVec_queue_fifo_62_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_62_vd = _sinkVec_queue_fifo_62_data_out[46:42];
  wire         sinkVec_queue_62_enq_ready = ~_sinkVec_queue_fifo_62_full;
  wire         sinkVec_queue_62_enq_valid;
  assign sinkVec_queue_62_deq_valid = ~_sinkVec_queue_fifo_62_empty | sinkVec_queue_62_enq_valid;
  assign sinkVec_queue_62_deq_bits_vd = _sinkVec_queue_fifo_62_empty ? sinkVec_queue_62_enq_bits_vd : sinkVec_queue_dataOut_62_vd;
  assign sinkVec_queue_62_deq_bits_offset = _sinkVec_queue_fifo_62_empty ? sinkVec_queue_62_enq_bits_offset : sinkVec_queue_dataOut_62_offset;
  assign sinkVec_queue_62_deq_bits_mask = _sinkVec_queue_fifo_62_empty ? sinkVec_queue_62_enq_bits_mask : sinkVec_queue_dataOut_62_mask;
  assign sinkVec_queue_62_deq_bits_data = _sinkVec_queue_fifo_62_empty ? sinkVec_queue_62_enq_bits_data : sinkVec_queue_dataOut_62_data;
  assign sinkVec_queue_62_deq_bits_last = ~_sinkVec_queue_fifo_62_empty & sinkVec_queue_dataOut_62_last;
  assign sinkVec_queue_62_deq_bits_instructionIndex = _sinkVec_queue_fifo_62_empty ? sinkVec_queue_62_enq_bits_instructionIndex : sinkVec_queue_dataOut_62_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_62;
  wire         sinkVec_releasePipe_pipe_out_62_valid = sinkVec_releasePipe_pipe_v_62;
  wire         x22_15_0_ready;
  wire         x22_15_0_valid;
  wire         sinkVec_validSource_62_valid = x22_15_0_ready & x22_15_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_62;
  wire [2:0]   sinkVec_tokenCheck_counterChange_62 = sinkVec_validSource_62_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_62 = ~(sinkVec_tokenCheck_counter_62[2]);
  assign x22_15_0_ready = sinkVec_tokenCheck_62;
  assign sinkVec_queue_62_enq_valid = sinkVec_validSink_62_valid;
  assign sinkVec_queue_62_enq_bits_vd = sinkVec_validSink_62_bits_vd;
  assign sinkVec_queue_62_enq_bits_offset = sinkVec_validSink_62_bits_offset;
  assign sinkVec_queue_62_enq_bits_mask = sinkVec_validSink_62_bits_mask;
  assign sinkVec_queue_62_enq_bits_data = sinkVec_validSink_62_bits_data;
  assign sinkVec_queue_62_enq_bits_instructionIndex = sinkVec_validSink_62_bits_instructionIndex;
  reg          sinkVec_shifterReg_62_0_valid;
  assign sinkVec_validSink_62_valid = sinkVec_shifterReg_62_0_valid;
  reg  [4:0]   sinkVec_shifterReg_62_0_bits_vd;
  assign sinkVec_validSink_62_bits_vd = sinkVec_shifterReg_62_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_62_0_bits_offset;
  assign sinkVec_validSink_62_bits_offset = sinkVec_shifterReg_62_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_62_0_bits_mask;
  assign sinkVec_validSink_62_bits_mask = sinkVec_shifterReg_62_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_62_0_bits_data;
  assign sinkVec_validSink_62_bits_data = sinkVec_shifterReg_62_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_62_0_bits_instructionIndex;
  assign sinkVec_validSink_62_bits_instructionIndex = sinkVec_shifterReg_62_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_62 = sinkVec_shifterReg_62_0_valid | sinkVec_validSource_62_valid;
  wire         sinkVec_31_1_ready;
  wire         sinkVec_queue_63_deq_ready = sinkVec_sinkWire_63_ready;
  wire         sinkVec_queue_63_deq_valid;
  wire [4:0]   sinkVec_queue_63_deq_bits_vd;
  wire         sinkVec_31_1_valid = sinkVec_sinkWire_63_valid;
  wire [1:0]   sinkVec_queue_63_deq_bits_offset;
  wire [4:0]   sinkVec_31_1_bits_vd = sinkVec_sinkWire_63_bits_vd;
  wire [3:0]   sinkVec_queue_63_deq_bits_mask;
  wire [1:0]   sinkVec_31_1_bits_offset = sinkVec_sinkWire_63_bits_offset;
  wire [31:0]  sinkVec_queue_63_deq_bits_data;
  wire [3:0]   sinkVec_31_1_bits_mask = sinkVec_sinkWire_63_bits_mask;
  wire         sinkVec_queue_63_deq_bits_last;
  wire [31:0]  sinkVec_31_1_bits_data = sinkVec_sinkWire_63_bits_data;
  wire [2:0]   sinkVec_queue_63_deq_bits_instructionIndex;
  wire         sinkVec_31_1_bits_last = sinkVec_sinkWire_63_bits_last;
  wire [2:0]   sinkVec_31_1_bits_instructionIndex = sinkVec_sinkWire_63_bits_instructionIndex;
  wire         sinkVec_validSink_63_valid;
  wire [4:0]   sinkVec_validSink_63_bits_vd;
  wire [1:0]   sinkVec_validSink_63_bits_offset;
  wire [3:0]   sinkVec_validSink_63_bits_mask;
  wire [31:0]  sinkVec_validSink_63_bits_data;
  wire         sinkVec_validSink_63_bits_last;
  wire [2:0]   sinkVec_validSink_63_bits_instructionIndex;
  assign sinkVec_sinkWire_63_valid = sinkVec_queue_63_deq_valid;
  assign sinkVec_sinkWire_63_bits_vd = sinkVec_queue_63_deq_bits_vd;
  assign sinkVec_sinkWire_63_bits_offset = sinkVec_queue_63_deq_bits_offset;
  assign sinkVec_sinkWire_63_bits_mask = sinkVec_queue_63_deq_bits_mask;
  assign sinkVec_sinkWire_63_bits_data = sinkVec_queue_63_deq_bits_data;
  assign sinkVec_sinkWire_63_bits_last = sinkVec_queue_63_deq_bits_last;
  assign sinkVec_sinkWire_63_bits_instructionIndex = sinkVec_queue_63_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_63_enq_bits_data;
  wire         sinkVec_queue_63_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_31 = {sinkVec_queue_63_enq_bits_data, sinkVec_queue_63_enq_bits_last};
  wire [2:0]   sinkVec_queue_63_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_63 = {sinkVec_queue_dataIn_lo_hi_31, sinkVec_queue_63_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_63_enq_bits_vd;
  wire [1:0]   sinkVec_queue_63_enq_bits_offset;
  wire [6:0]   sinkVec_queue_dataIn_hi_hi_31 = {sinkVec_queue_63_enq_bits_vd, sinkVec_queue_63_enq_bits_offset};
  wire [3:0]   sinkVec_queue_63_enq_bits_mask;
  wire [10:0]  sinkVec_queue_dataIn_hi_63 = {sinkVec_queue_dataIn_hi_hi_31, sinkVec_queue_63_enq_bits_mask};
  wire [46:0]  sinkVec_queue_dataIn_63 = {sinkVec_queue_dataIn_hi_63, sinkVec_queue_dataIn_lo_63};
  wire [2:0]   sinkVec_queue_dataOut_63_instructionIndex = _sinkVec_queue_fifo_63_data_out[2:0];
  wire         sinkVec_queue_dataOut_63_last = _sinkVec_queue_fifo_63_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_63_data = _sinkVec_queue_fifo_63_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_63_mask = _sinkVec_queue_fifo_63_data_out[39:36];
  wire [1:0]   sinkVec_queue_dataOut_63_offset = _sinkVec_queue_fifo_63_data_out[41:40];
  wire [4:0]   sinkVec_queue_dataOut_63_vd = _sinkVec_queue_fifo_63_data_out[46:42];
  wire         sinkVec_queue_63_enq_ready = ~_sinkVec_queue_fifo_63_full;
  wire         sinkVec_queue_63_enq_valid;
  assign sinkVec_queue_63_deq_valid = ~_sinkVec_queue_fifo_63_empty | sinkVec_queue_63_enq_valid;
  assign sinkVec_queue_63_deq_bits_vd = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_vd : sinkVec_queue_dataOut_63_vd;
  assign sinkVec_queue_63_deq_bits_offset = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_offset : sinkVec_queue_dataOut_63_offset;
  assign sinkVec_queue_63_deq_bits_mask = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_mask : sinkVec_queue_dataOut_63_mask;
  assign sinkVec_queue_63_deq_bits_data = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_data : sinkVec_queue_dataOut_63_data;
  assign sinkVec_queue_63_deq_bits_last = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_last : sinkVec_queue_dataOut_63_last;
  assign sinkVec_queue_63_deq_bits_instructionIndex = _sinkVec_queue_fifo_63_empty ? sinkVec_queue_63_enq_bits_instructionIndex : sinkVec_queue_dataOut_63_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_63;
  wire         sinkVec_releasePipe_pipe_out_63_valid = sinkVec_releasePipe_pipe_v_63;
  wire         x22_15_1_ready;
  wire         x22_15_1_valid;
  wire         sinkVec_validSource_63_valid = x22_15_1_ready & x22_15_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_63;
  wire [2:0]   sinkVec_tokenCheck_counterChange_63 = sinkVec_validSource_63_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_63 = ~(sinkVec_tokenCheck_counter_63[2]);
  assign x22_15_1_ready = sinkVec_tokenCheck_63;
  assign sinkVec_queue_63_enq_valid = sinkVec_validSink_63_valid;
  assign sinkVec_queue_63_enq_bits_vd = sinkVec_validSink_63_bits_vd;
  assign sinkVec_queue_63_enq_bits_offset = sinkVec_validSink_63_bits_offset;
  assign sinkVec_queue_63_enq_bits_mask = sinkVec_validSink_63_bits_mask;
  assign sinkVec_queue_63_enq_bits_data = sinkVec_validSink_63_bits_data;
  assign sinkVec_queue_63_enq_bits_last = sinkVec_validSink_63_bits_last;
  assign sinkVec_queue_63_enq_bits_instructionIndex = sinkVec_validSink_63_bits_instructionIndex;
  reg          sinkVec_shifterReg_63_0_valid;
  assign sinkVec_validSink_63_valid = sinkVec_shifterReg_63_0_valid;
  reg  [4:0]   sinkVec_shifterReg_63_0_bits_vd;
  assign sinkVec_validSink_63_bits_vd = sinkVec_shifterReg_63_0_bits_vd;
  reg  [1:0]   sinkVec_shifterReg_63_0_bits_offset;
  assign sinkVec_validSink_63_bits_offset = sinkVec_shifterReg_63_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_63_0_bits_mask;
  assign sinkVec_validSink_63_bits_mask = sinkVec_shifterReg_63_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_63_0_bits_data;
  assign sinkVec_validSink_63_bits_data = sinkVec_shifterReg_63_0_bits_data;
  reg          sinkVec_shifterReg_63_0_bits_last;
  assign sinkVec_validSink_63_bits_last = sinkVec_shifterReg_63_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_63_0_bits_instructionIndex;
  assign sinkVec_validSink_63_bits_instructionIndex = sinkVec_shifterReg_63_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_63 = sinkVec_shifterReg_63_0_valid | sinkVec_validSource_63_valid;
  assign sinkVec_sinkWire_62_ready = sinkVec_31_0_ready;
  assign sinkVec_sinkWire_63_ready = sinkVec_31_1_ready;
  reg          maskUnitFirst_31;
  wire         tryToRead_31 = sinkVec_31_0_valid | sinkVec_31_1_valid;
  wire         sinkWire_31_valid = maskUnitFirst_31 ? sinkVec_31_0_valid : sinkVec_31_1_valid;
  wire [4:0]   sinkWire_31_bits_vd = maskUnitFirst_31 ? sinkVec_31_0_bits_vd : sinkVec_31_1_bits_vd;
  wire [1:0]   sinkWire_31_bits_offset = maskUnitFirst_31 ? sinkVec_31_0_bits_offset : sinkVec_31_1_bits_offset;
  wire [3:0]   sinkWire_31_bits_mask = maskUnitFirst_31 ? sinkVec_31_0_bits_mask : sinkVec_31_1_bits_mask;
  wire [31:0]  sinkWire_31_bits_data = maskUnitFirst_31 ? sinkVec_31_0_bits_data : sinkVec_31_1_bits_data;
  wire         sinkWire_31_bits_last = maskUnitFirst_31 ? sinkVec_31_0_bits_last : sinkVec_31_1_bits_last;
  wire [2:0]   sinkWire_31_bits_instructionIndex = maskUnitFirst_31 ? sinkVec_31_0_bits_instructionIndex : sinkVec_31_1_bits_instructionIndex;
  wire         sinkWire_31_ready;
  assign sinkVec_31_1_ready = sinkWire_31_ready & ~maskUnitFirst_31;
  assign sinkVec_31_0_ready = sinkWire_31_ready & maskUnitFirst_31;
  reg          view__writeRelease_15_pipe_v;
  wire         view__writeRelease_15_pipe_out_valid = view__writeRelease_15_pipe_v;
  reg          pipe_v_45;
  wire         pipe_out_30_valid = pipe_v_45;
  wire         _probeWire_writeQueueEnqVec_15_valid_T = x22_15_0_ready & _maskUnit_exeResp_15_valid;
  reg          instructionFinishedPipe_pipe_v_15;
  wire         instructionFinishedPipe_pipe_out_15_valid = instructionFinishedPipe_pipe_v_15;
  reg  [7:0]   instructionFinishedPipe_pipe_b_15;
  wire [7:0]   instructionFinishedPipe_pipe_out_15_bits = instructionFinishedPipe_pipe_b_15;
  wire         instructionFinished_15_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_15_bits);
  wire         instructionFinished_15_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_15_bits);
  wire         instructionFinished_15_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_15_bits);
  wire         instructionFinished_15_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_15_bits);
  assign vxsatReportVec_15 = _laneVec_15_vxsatReport[3:0];
  reg          pipe_v_46;
  reg  [31:0]  pipe_b_46;
  reg          pipe_pipe_v_15;
  wire         pipe_pipe_out_15_valid = pipe_pipe_v_15;
  reg  [31:0]  pipe_pipe_b_15;
  wire [31:0]  pipe_pipe_out_15_bits = pipe_pipe_b_15;
  reg          view__laneMaskSelect_15_pipe_v;
  reg  [5:0]   view__laneMaskSelect_15_pipe_b;
  reg          view__laneMaskSelect_15_pipe_pipe_v;
  wire         view__laneMaskSelect_15_pipe_pipe_out_valid = view__laneMaskSelect_15_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_15_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_15_pipe_pipe_out_bits = view__laneMaskSelect_15_pipe_pipe_b;
  reg          view__laneMaskSewSelect_15_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_15_pipe_b;
  reg          view__laneMaskSewSelect_15_pipe_pipe_v;
  wire         view__laneMaskSewSelect_15_pipe_pipe_out_valid = view__laneMaskSewSelect_15_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_15_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_15_pipe_pipe_out_bits = view__laneMaskSewSelect_15_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_15;
  wire         lsuLastPipe_pipe_out_15_valid = lsuLastPipe_pipe_v_15;
  reg  [7:0]   lsuLastPipe_pipe_b_15;
  wire [7:0]   lsuLastPipe_pipe_out_15_bits = lsuLastPipe_pipe_b_15;
  reg          maskLastPipe_pipe_v_15;
  wire         maskLastPipe_pipe_out_15_valid = maskLastPipe_pipe_v_15;
  reg  [7:0]   maskLastPipe_pipe_b_15;
  wire [7:0]   maskLastPipe_pipe_out_15_bits = maskLastPipe_pipe_b_15;
  wire [5:0]   writeCounter_15 = requestReg_bits_writeByte[11:6] + {5'h0, requestReg_bits_writeByte[5:0] > 6'h3C};
  reg          pipe_v_47;
  wire         pipe_out_31_valid = pipe_v_47;
  reg  [5:0]   pipe_b_47;
  wire [5:0]   pipe_out_31_bits = pipe_b_47;
  reg          pipe_v_48;
  wire         pipe_out_32_valid = pipe_v_48;
  reg          shifterReg_48_0_valid;
  reg  [31:0]  shifterReg_48_0_bits_data;
  wire         shifterValid_48 = shifterReg_48_0_valid | _laneVec_0_readBusPort_0_deq_valid;
  reg          pipe_v_49;
  wire         pipe_out_33_valid = pipe_v_49;
  reg          shifterReg_49_0_valid;
  reg  [31:0]  shifterReg_49_0_bits_data;
  reg  [1:0]   shifterReg_49_0_bits_mask;
  reg  [2:0]   shifterReg_49_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_49_0_bits_counter;
  wire         shifterValid_49 = shifterReg_49_0_valid | _laneVec_0_writeBusPort_0_deq_valid;
  reg          pipe_v_50;
  wire         pipe_out_34_valid = pipe_v_50;
  reg          shifterReg_50_0_valid;
  reg  [31:0]  shifterReg_50_0_bits_data;
  wire         shifterValid_50 = shifterReg_50_0_valid | _laneVec_1_readBusPort_0_deq_valid;
  reg          pipe_v_51;
  wire         pipe_out_35_valid = pipe_v_51;
  reg          shifterReg_51_0_valid;
  reg  [31:0]  shifterReg_51_0_bits_data;
  reg  [1:0]   shifterReg_51_0_bits_mask;
  reg  [2:0]   shifterReg_51_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_51_0_bits_counter;
  wire         shifterValid_51 = shifterReg_51_0_valid | _laneVec_0_writeBusPort_1_deq_valid;
  reg          pipe_v_52;
  wire         pipe_out_36_valid = pipe_v_52;
  reg          shifterReg_52_0_valid;
  reg  [31:0]  shifterReg_52_0_bits_data;
  wire         shifterValid_52 = shifterReg_52_0_valid | _laneVec_2_readBusPort_0_deq_valid;
  reg          pipe_v_53;
  wire         pipe_out_37_valid = pipe_v_53;
  reg          shifterReg_53_0_valid;
  reg  [31:0]  shifterReg_53_0_bits_data;
  reg  [1:0]   shifterReg_53_0_bits_mask;
  reg  [2:0]   shifterReg_53_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_53_0_bits_counter;
  wire         shifterValid_53 = shifterReg_53_0_valid | _laneVec_1_writeBusPort_0_deq_valid;
  reg          pipe_v_54;
  wire         pipe_out_38_valid = pipe_v_54;
  reg          shifterReg_54_0_valid;
  reg  [31:0]  shifterReg_54_0_bits_data;
  wire         shifterValid_54 = shifterReg_54_0_valid | _laneVec_3_readBusPort_0_deq_valid;
  reg          pipe_v_55;
  wire         pipe_out_39_valid = pipe_v_55;
  reg          shifterReg_55_0_valid;
  reg  [31:0]  shifterReg_55_0_bits_data;
  reg  [1:0]   shifterReg_55_0_bits_mask;
  reg  [2:0]   shifterReg_55_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_55_0_bits_counter;
  wire         shifterValid_55 = shifterReg_55_0_valid | _laneVec_1_writeBusPort_1_deq_valid;
  reg          pipe_v_56;
  wire         pipe_out_40_valid = pipe_v_56;
  reg          shifterReg_56_0_valid;
  reg  [31:0]  shifterReg_56_0_bits_data;
  wire         shifterValid_56 = shifterReg_56_0_valid | _laneVec_4_readBusPort_0_deq_valid;
  reg          pipe_v_57;
  wire         pipe_out_41_valid = pipe_v_57;
  reg          shifterReg_57_0_valid;
  reg  [31:0]  shifterReg_57_0_bits_data;
  reg  [1:0]   shifterReg_57_0_bits_mask;
  reg  [2:0]   shifterReg_57_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_57_0_bits_counter;
  wire         shifterValid_57 = shifterReg_57_0_valid | _laneVec_2_writeBusPort_0_deq_valid;
  reg          pipe_v_58;
  wire         pipe_out_42_valid = pipe_v_58;
  reg          shifterReg_58_0_valid;
  reg  [31:0]  shifterReg_58_0_bits_data;
  wire         shifterValid_58 = shifterReg_58_0_valid | _laneVec_5_readBusPort_0_deq_valid;
  reg          pipe_v_59;
  wire         pipe_out_43_valid = pipe_v_59;
  reg          shifterReg_59_0_valid;
  reg  [31:0]  shifterReg_59_0_bits_data;
  reg  [1:0]   shifterReg_59_0_bits_mask;
  reg  [2:0]   shifterReg_59_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_59_0_bits_counter;
  wire         shifterValid_59 = shifterReg_59_0_valid | _laneVec_2_writeBusPort_1_deq_valid;
  reg          pipe_v_60;
  wire         pipe_out_44_valid = pipe_v_60;
  reg          shifterReg_60_0_valid;
  reg  [31:0]  shifterReg_60_0_bits_data;
  wire         shifterValid_60 = shifterReg_60_0_valid | _laneVec_6_readBusPort_0_deq_valid;
  reg          pipe_v_61;
  wire         pipe_out_45_valid = pipe_v_61;
  reg          shifterReg_61_0_valid;
  reg  [31:0]  shifterReg_61_0_bits_data;
  reg  [1:0]   shifterReg_61_0_bits_mask;
  reg  [2:0]   shifterReg_61_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_61_0_bits_counter;
  wire         shifterValid_61 = shifterReg_61_0_valid | _laneVec_3_writeBusPort_0_deq_valid;
  reg          pipe_v_62;
  wire         pipe_out_46_valid = pipe_v_62;
  reg          shifterReg_62_0_valid;
  reg  [31:0]  shifterReg_62_0_bits_data;
  wire         shifterValid_62 = shifterReg_62_0_valid | _laneVec_7_readBusPort_0_deq_valid;
  reg          pipe_v_63;
  wire         pipe_out_47_valid = pipe_v_63;
  reg          shifterReg_63_0_valid;
  reg  [31:0]  shifterReg_63_0_bits_data;
  reg  [1:0]   shifterReg_63_0_bits_mask;
  reg  [2:0]   shifterReg_63_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_63_0_bits_counter;
  wire         shifterValid_63 = shifterReg_63_0_valid | _laneVec_3_writeBusPort_1_deq_valid;
  reg          pipe_v_64;
  wire         pipe_out_48_valid = pipe_v_64;
  reg          shifterReg_64_0_valid;
  reg  [31:0]  shifterReg_64_0_bits_data;
  wire         shifterValid_64 = shifterReg_64_0_valid | _laneVec_8_readBusPort_0_deq_valid;
  reg          pipe_v_65;
  wire         pipe_out_49_valid = pipe_v_65;
  reg          shifterReg_65_0_valid;
  reg  [31:0]  shifterReg_65_0_bits_data;
  reg  [1:0]   shifterReg_65_0_bits_mask;
  reg  [2:0]   shifterReg_65_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_65_0_bits_counter;
  wire         shifterValid_65 = shifterReg_65_0_valid | _laneVec_4_writeBusPort_0_deq_valid;
  reg          pipe_v_66;
  wire         pipe_out_50_valid = pipe_v_66;
  reg          shifterReg_66_0_valid;
  reg  [31:0]  shifterReg_66_0_bits_data;
  wire         shifterValid_66 = shifterReg_66_0_valid | _laneVec_9_readBusPort_0_deq_valid;
  reg          pipe_v_67;
  wire         pipe_out_51_valid = pipe_v_67;
  reg          shifterReg_67_0_valid;
  reg  [31:0]  shifterReg_67_0_bits_data;
  reg  [1:0]   shifterReg_67_0_bits_mask;
  reg  [2:0]   shifterReg_67_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_67_0_bits_counter;
  wire         shifterValid_67 = shifterReg_67_0_valid | _laneVec_4_writeBusPort_1_deq_valid;
  reg          pipe_v_68;
  wire         pipe_out_52_valid = pipe_v_68;
  reg          shifterReg_68_0_valid;
  reg  [31:0]  shifterReg_68_0_bits_data;
  wire         shifterValid_68 = shifterReg_68_0_valid | _laneVec_10_readBusPort_0_deq_valid;
  reg          pipe_v_69;
  wire         pipe_out_53_valid = pipe_v_69;
  reg          shifterReg_69_0_valid;
  reg  [31:0]  shifterReg_69_0_bits_data;
  reg  [1:0]   shifterReg_69_0_bits_mask;
  reg  [2:0]   shifterReg_69_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_69_0_bits_counter;
  wire         shifterValid_69 = shifterReg_69_0_valid | _laneVec_5_writeBusPort_0_deq_valid;
  reg          pipe_v_70;
  wire         pipe_out_54_valid = pipe_v_70;
  reg          shifterReg_70_0_valid;
  reg  [31:0]  shifterReg_70_0_bits_data;
  wire         shifterValid_70 = shifterReg_70_0_valid | _laneVec_11_readBusPort_0_deq_valid;
  reg          pipe_v_71;
  wire         pipe_out_55_valid = pipe_v_71;
  reg          shifterReg_71_0_valid;
  reg  [31:0]  shifterReg_71_0_bits_data;
  reg  [1:0]   shifterReg_71_0_bits_mask;
  reg  [2:0]   shifterReg_71_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_71_0_bits_counter;
  wire         shifterValid_71 = shifterReg_71_0_valid | _laneVec_5_writeBusPort_1_deq_valid;
  reg          pipe_v_72;
  wire         pipe_out_56_valid = pipe_v_72;
  reg          shifterReg_72_0_valid;
  reg  [31:0]  shifterReg_72_0_bits_data;
  wire         shifterValid_72 = shifterReg_72_0_valid | _laneVec_12_readBusPort_0_deq_valid;
  reg          pipe_v_73;
  wire         pipe_out_57_valid = pipe_v_73;
  reg          shifterReg_73_0_valid;
  reg  [31:0]  shifterReg_73_0_bits_data;
  reg  [1:0]   shifterReg_73_0_bits_mask;
  reg  [2:0]   shifterReg_73_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_73_0_bits_counter;
  wire         shifterValid_73 = shifterReg_73_0_valid | _laneVec_6_writeBusPort_0_deq_valid;
  reg          pipe_v_74;
  wire         pipe_out_58_valid = pipe_v_74;
  reg          shifterReg_74_0_valid;
  reg  [31:0]  shifterReg_74_0_bits_data;
  wire         shifterValid_74 = shifterReg_74_0_valid | _laneVec_13_readBusPort_0_deq_valid;
  reg          pipe_v_75;
  wire         pipe_out_59_valid = pipe_v_75;
  reg          shifterReg_75_0_valid;
  reg  [31:0]  shifterReg_75_0_bits_data;
  reg  [1:0]   shifterReg_75_0_bits_mask;
  reg  [2:0]   shifterReg_75_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_75_0_bits_counter;
  wire         shifterValid_75 = shifterReg_75_0_valid | _laneVec_6_writeBusPort_1_deq_valid;
  reg          pipe_v_76;
  wire         pipe_out_60_valid = pipe_v_76;
  reg          shifterReg_76_0_valid;
  reg  [31:0]  shifterReg_76_0_bits_data;
  wire         shifterValid_76 = shifterReg_76_0_valid | _laneVec_14_readBusPort_0_deq_valid;
  reg          pipe_v_77;
  wire         pipe_out_61_valid = pipe_v_77;
  reg          shifterReg_77_0_valid;
  reg  [31:0]  shifterReg_77_0_bits_data;
  reg  [1:0]   shifterReg_77_0_bits_mask;
  reg  [2:0]   shifterReg_77_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_77_0_bits_counter;
  wire         shifterValid_77 = shifterReg_77_0_valid | _laneVec_7_writeBusPort_0_deq_valid;
  reg          pipe_v_78;
  wire         pipe_out_62_valid = pipe_v_78;
  reg          shifterReg_78_0_valid;
  reg  [31:0]  shifterReg_78_0_bits_data;
  wire         shifterValid_78 = shifterReg_78_0_valid | _laneVec_15_readBusPort_0_deq_valid;
  reg          pipe_v_79;
  wire         pipe_out_63_valid = pipe_v_79;
  reg          shifterReg_79_0_valid;
  reg  [31:0]  shifterReg_79_0_bits_data;
  reg  [1:0]   shifterReg_79_0_bits_mask;
  reg  [2:0]   shifterReg_79_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_79_0_bits_counter;
  wire         shifterValid_79 = shifterReg_79_0_valid | _laneVec_7_writeBusPort_1_deq_valid;
  reg          pipe_v_80;
  wire         pipe_out_64_valid = pipe_v_80;
  reg          shifterReg_80_0_valid;
  reg  [31:0]  shifterReg_80_0_bits_data;
  wire         shifterValid_80 = shifterReg_80_0_valid | _laneVec_0_readBusPort_1_deq_valid;
  reg          pipe_v_81;
  wire         pipe_out_65_valid = pipe_v_81;
  reg          shifterReg_81_0_valid;
  reg  [31:0]  shifterReg_81_0_bits_data;
  reg  [1:0]   shifterReg_81_0_bits_mask;
  reg  [2:0]   shifterReg_81_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_81_0_bits_counter;
  wire         shifterValid_81 = shifterReg_81_0_valid | _laneVec_8_writeBusPort_0_deq_valid;
  reg          pipe_v_82;
  wire         pipe_out_66_valid = pipe_v_82;
  reg          shifterReg_82_0_valid;
  reg  [31:0]  shifterReg_82_0_bits_data;
  wire         shifterValid_82 = shifterReg_82_0_valid | _laneVec_1_readBusPort_1_deq_valid;
  reg          pipe_v_83;
  wire         pipe_out_67_valid = pipe_v_83;
  reg          shifterReg_83_0_valid;
  reg  [31:0]  shifterReg_83_0_bits_data;
  reg  [1:0]   shifterReg_83_0_bits_mask;
  reg  [2:0]   shifterReg_83_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_83_0_bits_counter;
  wire         shifterValid_83 = shifterReg_83_0_valid | _laneVec_8_writeBusPort_1_deq_valid;
  reg          pipe_v_84;
  wire         pipe_out_68_valid = pipe_v_84;
  reg          shifterReg_84_0_valid;
  reg  [31:0]  shifterReg_84_0_bits_data;
  wire         shifterValid_84 = shifterReg_84_0_valid | _laneVec_2_readBusPort_1_deq_valid;
  reg          pipe_v_85;
  wire         pipe_out_69_valid = pipe_v_85;
  reg          shifterReg_85_0_valid;
  reg  [31:0]  shifterReg_85_0_bits_data;
  reg  [1:0]   shifterReg_85_0_bits_mask;
  reg  [2:0]   shifterReg_85_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_85_0_bits_counter;
  wire         shifterValid_85 = shifterReg_85_0_valid | _laneVec_9_writeBusPort_0_deq_valid;
  reg          pipe_v_86;
  wire         pipe_out_70_valid = pipe_v_86;
  reg          shifterReg_86_0_valid;
  reg  [31:0]  shifterReg_86_0_bits_data;
  wire         shifterValid_86 = shifterReg_86_0_valid | _laneVec_3_readBusPort_1_deq_valid;
  reg          pipe_v_87;
  wire         pipe_out_71_valid = pipe_v_87;
  reg          shifterReg_87_0_valid;
  reg  [31:0]  shifterReg_87_0_bits_data;
  reg  [1:0]   shifterReg_87_0_bits_mask;
  reg  [2:0]   shifterReg_87_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_87_0_bits_counter;
  wire         shifterValid_87 = shifterReg_87_0_valid | _laneVec_9_writeBusPort_1_deq_valid;
  reg          pipe_v_88;
  wire         pipe_out_72_valid = pipe_v_88;
  reg          shifterReg_88_0_valid;
  reg  [31:0]  shifterReg_88_0_bits_data;
  wire         shifterValid_88 = shifterReg_88_0_valid | _laneVec_4_readBusPort_1_deq_valid;
  reg          pipe_v_89;
  wire         pipe_out_73_valid = pipe_v_89;
  reg          shifterReg_89_0_valid;
  reg  [31:0]  shifterReg_89_0_bits_data;
  reg  [1:0]   shifterReg_89_0_bits_mask;
  reg  [2:0]   shifterReg_89_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_89_0_bits_counter;
  wire         shifterValid_89 = shifterReg_89_0_valid | _laneVec_10_writeBusPort_0_deq_valid;
  reg          pipe_v_90;
  wire         pipe_out_74_valid = pipe_v_90;
  reg          shifterReg_90_0_valid;
  reg  [31:0]  shifterReg_90_0_bits_data;
  wire         shifterValid_90 = shifterReg_90_0_valid | _laneVec_5_readBusPort_1_deq_valid;
  reg          pipe_v_91;
  wire         pipe_out_75_valid = pipe_v_91;
  reg          shifterReg_91_0_valid;
  reg  [31:0]  shifterReg_91_0_bits_data;
  reg  [1:0]   shifterReg_91_0_bits_mask;
  reg  [2:0]   shifterReg_91_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_91_0_bits_counter;
  wire         shifterValid_91 = shifterReg_91_0_valid | _laneVec_10_writeBusPort_1_deq_valid;
  reg          pipe_v_92;
  wire         pipe_out_76_valid = pipe_v_92;
  reg          shifterReg_92_0_valid;
  reg  [31:0]  shifterReg_92_0_bits_data;
  wire         shifterValid_92 = shifterReg_92_0_valid | _laneVec_6_readBusPort_1_deq_valid;
  reg          pipe_v_93;
  wire         pipe_out_77_valid = pipe_v_93;
  reg          shifterReg_93_0_valid;
  reg  [31:0]  shifterReg_93_0_bits_data;
  reg  [1:0]   shifterReg_93_0_bits_mask;
  reg  [2:0]   shifterReg_93_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_93_0_bits_counter;
  wire         shifterValid_93 = shifterReg_93_0_valid | _laneVec_11_writeBusPort_0_deq_valid;
  reg          pipe_v_94;
  wire         pipe_out_78_valid = pipe_v_94;
  reg          shifterReg_94_0_valid;
  reg  [31:0]  shifterReg_94_0_bits_data;
  wire         shifterValid_94 = shifterReg_94_0_valid | _laneVec_7_readBusPort_1_deq_valid;
  reg          pipe_v_95;
  wire         pipe_out_79_valid = pipe_v_95;
  reg          shifterReg_95_0_valid;
  reg  [31:0]  shifterReg_95_0_bits_data;
  reg  [1:0]   shifterReg_95_0_bits_mask;
  reg  [2:0]   shifterReg_95_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_95_0_bits_counter;
  wire         shifterValid_95 = shifterReg_95_0_valid | _laneVec_11_writeBusPort_1_deq_valid;
  reg          pipe_v_96;
  wire         pipe_out_80_valid = pipe_v_96;
  reg          shifterReg_96_0_valid;
  reg  [31:0]  shifterReg_96_0_bits_data;
  wire         shifterValid_96 = shifterReg_96_0_valid | _laneVec_8_readBusPort_1_deq_valid;
  reg          pipe_v_97;
  wire         pipe_out_81_valid = pipe_v_97;
  reg          shifterReg_97_0_valid;
  reg  [31:0]  shifterReg_97_0_bits_data;
  reg  [1:0]   shifterReg_97_0_bits_mask;
  reg  [2:0]   shifterReg_97_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_97_0_bits_counter;
  wire         shifterValid_97 = shifterReg_97_0_valid | _laneVec_12_writeBusPort_0_deq_valid;
  reg          pipe_v_98;
  wire         pipe_out_82_valid = pipe_v_98;
  reg          shifterReg_98_0_valid;
  reg  [31:0]  shifterReg_98_0_bits_data;
  wire         shifterValid_98 = shifterReg_98_0_valid | _laneVec_9_readBusPort_1_deq_valid;
  reg          pipe_v_99;
  wire         pipe_out_83_valid = pipe_v_99;
  reg          shifterReg_99_0_valid;
  reg  [31:0]  shifterReg_99_0_bits_data;
  reg  [1:0]   shifterReg_99_0_bits_mask;
  reg  [2:0]   shifterReg_99_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_99_0_bits_counter;
  wire         shifterValid_99 = shifterReg_99_0_valid | _laneVec_12_writeBusPort_1_deq_valid;
  reg          pipe_v_100;
  wire         pipe_out_84_valid = pipe_v_100;
  reg          shifterReg_100_0_valid;
  reg  [31:0]  shifterReg_100_0_bits_data;
  wire         shifterValid_100 = shifterReg_100_0_valid | _laneVec_10_readBusPort_1_deq_valid;
  reg          pipe_v_101;
  wire         pipe_out_85_valid = pipe_v_101;
  reg          shifterReg_101_0_valid;
  reg  [31:0]  shifterReg_101_0_bits_data;
  reg  [1:0]   shifterReg_101_0_bits_mask;
  reg  [2:0]   shifterReg_101_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_101_0_bits_counter;
  wire         shifterValid_101 = shifterReg_101_0_valid | _laneVec_13_writeBusPort_0_deq_valid;
  reg          pipe_v_102;
  wire         pipe_out_86_valid = pipe_v_102;
  reg          shifterReg_102_0_valid;
  reg  [31:0]  shifterReg_102_0_bits_data;
  wire         shifterValid_102 = shifterReg_102_0_valid | _laneVec_11_readBusPort_1_deq_valid;
  reg          pipe_v_103;
  wire         pipe_out_87_valid = pipe_v_103;
  reg          shifterReg_103_0_valid;
  reg  [31:0]  shifterReg_103_0_bits_data;
  reg  [1:0]   shifterReg_103_0_bits_mask;
  reg  [2:0]   shifterReg_103_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_103_0_bits_counter;
  wire         shifterValid_103 = shifterReg_103_0_valid | _laneVec_13_writeBusPort_1_deq_valid;
  reg          pipe_v_104;
  wire         pipe_out_88_valid = pipe_v_104;
  reg          shifterReg_104_0_valid;
  reg  [31:0]  shifterReg_104_0_bits_data;
  wire         shifterValid_104 = shifterReg_104_0_valid | _laneVec_12_readBusPort_1_deq_valid;
  reg          pipe_v_105;
  wire         pipe_out_89_valid = pipe_v_105;
  reg          shifterReg_105_0_valid;
  reg  [31:0]  shifterReg_105_0_bits_data;
  reg  [1:0]   shifterReg_105_0_bits_mask;
  reg  [2:0]   shifterReg_105_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_105_0_bits_counter;
  wire         shifterValid_105 = shifterReg_105_0_valid | _laneVec_14_writeBusPort_0_deq_valid;
  reg          pipe_v_106;
  wire         pipe_out_90_valid = pipe_v_106;
  reg          shifterReg_106_0_valid;
  reg  [31:0]  shifterReg_106_0_bits_data;
  wire         shifterValid_106 = shifterReg_106_0_valid | _laneVec_13_readBusPort_1_deq_valid;
  reg          pipe_v_107;
  wire         pipe_out_91_valid = pipe_v_107;
  reg          shifterReg_107_0_valid;
  reg  [31:0]  shifterReg_107_0_bits_data;
  reg  [1:0]   shifterReg_107_0_bits_mask;
  reg  [2:0]   shifterReg_107_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_107_0_bits_counter;
  wire         shifterValid_107 = shifterReg_107_0_valid | _laneVec_14_writeBusPort_1_deq_valid;
  reg          pipe_v_108;
  wire         pipe_out_92_valid = pipe_v_108;
  reg          shifterReg_108_0_valid;
  reg  [31:0]  shifterReg_108_0_bits_data;
  wire         shifterValid_108 = shifterReg_108_0_valid | _laneVec_14_readBusPort_1_deq_valid;
  reg          pipe_v_109;
  wire         pipe_out_93_valid = pipe_v_109;
  reg          shifterReg_109_0_valid;
  reg  [31:0]  shifterReg_109_0_bits_data;
  reg  [1:0]   shifterReg_109_0_bits_mask;
  reg  [2:0]   shifterReg_109_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_109_0_bits_counter;
  wire         shifterValid_109 = shifterReg_109_0_valid | _laneVec_15_writeBusPort_0_deq_valid;
  reg          pipe_v_110;
  wire         pipe_out_94_valid = pipe_v_110;
  reg          shifterReg_110_0_valid;
  reg  [31:0]  shifterReg_110_0_bits_data;
  wire         shifterValid_110 = shifterReg_110_0_valid | _laneVec_15_readBusPort_1_deq_valid;
  reg          pipe_v_111;
  wire         pipe_out_95_valid = pipe_v_111;
  reg          shifterReg_111_0_valid;
  reg  [31:0]  shifterReg_111_0_bits_data;
  reg  [1:0]   shifterReg_111_0_bits_mask;
  reg  [2:0]   shifterReg_111_0_bits_instructionIndex;
  reg  [5:0]   shifterReg_111_0_bits_counter;
  wire         shifterValid_111 = shifterReg_111_0_valid | _laneVec_15_writeBusPort_1_deq_valid;
  wire [3:0]   free = {free_hi, free_lo};
  wire         allSlotFree = &free;
  wire [1:0]   existMaskType_lo = {~slots_1_state_idle & slots_1_record_maskType, ~slots_0_state_idle & slots_0_record_maskType};
  wire [1:0]   existMaskType_hi = {~slots_3_state_idle & slots_3_record_maskType, ~slots_2_state_idle & slots_2_record_maskType};
  wire         existMaskType = |{existMaskType_hi, existMaskType_lo};
  wire [2:0]   _free1H_T_2 = free[2:0] | {free[1:0], 1'h0};
  wire [3:0]   free1H = {~(_free1H_T_2 | {_free1H_T_2[0], 2'h0}), 1'h1} & free;
  wire [3:0]   slotToEnqueue = specialInstruction ? 4'h8 : free1H;
  wire         instructionIndexFree =
    (slots_0_state_idle | slots_0_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]) & (slots_1_state_idle | slots_1_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0])
    & (slots_2_state_idle | slots_2_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]) & (slots_3_state_idle | slots_3_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]);
  wire         executionReady = (~isLoadStoreType | _lsu_request_ready) & (noOffsetReadLoadStore | allLaneReady);
  assign requestRegDequeue_ready = executionReady & slotReady & (~gatherNeedRead | _maskUnit_gatherData_valid) & _tokenManager_issueAllow & instructionIndexFree & olderCheck;
  wire [3:0]   instructionToSlotOH = maskUnit_gatherData_ready ? slotToEnqueue : 4'h0;
  wire         slotCommit_0 = slots_0_state_wMaskUnitLast & slots_0_state_wLast & slots_0_state_wVRFWrite & ~slots_0_state_sCommit & slots_0_record_instructionIndex == responseCounter;
  wire         slotCommit_1 = slots_1_state_wMaskUnitLast & slots_1_state_wLast & slots_1_state_wVRFWrite & ~slots_1_state_sCommit & slots_1_record_instructionIndex == responseCounter;
  wire         slotCommit_2 = slots_2_state_wMaskUnitLast & slots_2_state_wLast & slots_2_state_wVRFWrite & ~slots_2_state_sCommit & slots_2_record_instructionIndex == responseCounter;
  assign slotCommit_3 = slots_3_state_wMaskUnitLast & slots_3_state_wLast & slots_3_state_wVRFWrite & ~slots_3_state_sCommit & slots_3_record_instructionIndex == responseCounter;
  assign lastSlotCommit = slotCommit_3;
  wire [1:0]   _GEN_5 = {slotCommit_1, slotCommit_0};
  wire [1:0]   retire_lo;
  assign retire_lo = _GEN_5;
  wire [1:0]   view__retire_csr_bits_vxsat_lo;
  assign view__retire_csr_bits_vxsat_lo = _GEN_5;
  wire [1:0]   view__retire_mem_valid_lo;
  assign view__retire_mem_valid_lo = _GEN_5;
  wire [1:0]   _GEN_6 = {slotCommit_3, slotCommit_2};
  wire [1:0]   retire_hi;
  assign retire_hi = _GEN_6;
  wire [1:0]   view__retire_csr_bits_vxsat_hi;
  assign view__retire_csr_bits_vxsat_hi = _GEN_6;
  wire [1:0]   view__retire_mem_valid_hi;
  assign view__retire_mem_valid_hi = _GEN_6;
  wire         retire_1 = |{retire_hi, retire_lo};
  wire [1:0]   view__retire_csr_bits_vxsat_lo_1 = {slots_1_vxsat, slots_0_vxsat};
  wire [1:0]   view__retire_csr_bits_vxsat_hi_1 = {slots_3_vxsat, slots_2_vxsat};
  wire [31:0]  retire_csr_bits_vxsat_0 = {31'h0, |({view__retire_csr_bits_vxsat_hi, view__retire_csr_bits_vxsat_lo} & {view__retire_csr_bits_vxsat_hi_1, view__retire_csr_bits_vxsat_lo_1})};
  wire [1:0]   view__retire_mem_valid_lo_1 = {slots_1_record_isLoadStore, slots_0_record_isLoadStore};
  wire [1:0]   view__retire_mem_valid_hi_1 = {slots_3_record_isLoadStore, slots_2_record_isLoadStore};
  wire         retire_mem_valid_0 = |({view__retire_mem_valid_hi, view__retire_mem_valid_lo} & {view__retire_mem_valid_hi_1, view__retire_mem_valid_lo_1});
  wire [31:0]  accessDataSource_bits;
  wire [31:0]  accessDataSource_1_bits;
  wire [31:0]  accessDataSource_2_bits;
  wire [31:0]  accessDataSource_3_bits;
  wire [31:0]  accessDataSource_4_bits;
  wire [31:0]  accessDataSource_5_bits;
  wire [31:0]  accessDataSource_6_bits;
  wire [31:0]  accessDataSource_7_bits;
  wire [31:0]  accessDataSource_8_bits;
  wire [31:0]  accessDataSource_9_bits;
  wire [31:0]  accessDataSource_10_bits;
  wire [31:0]  accessDataSource_11_bits;
  wire [31:0]  accessDataSource_12_bits;
  wire [31:0]  accessDataSource_13_bits;
  wire [31:0]  accessDataSource_14_bits;
  wire [31:0]  accessDataSource_15_bits;
  wire [31:0]  accessDataSource_16_bits;
  wire [31:0]  accessDataSource_17_bits;
  wire [31:0]  accessDataSource_18_bits;
  wire [31:0]  accessDataSource_19_bits;
  wire [31:0]  accessDataSource_20_bits;
  wire [31:0]  accessDataSource_21_bits;
  wire [31:0]  accessDataSource_22_bits;
  wire [31:0]  accessDataSource_23_bits;
  wire [31:0]  accessDataSource_24_bits;
  wire [31:0]  accessDataSource_25_bits;
  wire [31:0]  accessDataSource_26_bits;
  wire [31:0]  accessDataSource_27_bits;
  wire [31:0]  accessDataSource_28_bits;
  wire [31:0]  accessDataSource_29_bits;
  wire [31:0]  accessDataSource_30_bits;
  wire [31:0]  accessDataSource_31_bits;
  always @(posedge clock) begin
    if (reset) begin
      instructionCounter <= 3'h0;
      responseCounter <= 3'h0;
      requestReg_valid <= 1'h0;
      requestReg_bits_issue_instruction <= 32'h0;
      requestReg_bits_issue_rs1Data <= 32'h0;
      requestReg_bits_issue_rs2Data <= 32'h0;
      requestReg_bits_issue_vtype <= 32'h0;
      requestReg_bits_issue_vl <= 32'h0;
      requestReg_bits_issue_vstart <= 32'h0;
      requestReg_bits_issue_vcsr <= 32'h0;
      requestReg_bits_decodeResult_orderReduce <= 1'h0;
      requestReg_bits_decodeResult_floatMul <= 1'h0;
      requestReg_bits_decodeResult_fpExecutionType <= 2'h0;
      requestReg_bits_decodeResult_float <= 1'h0;
      requestReg_bits_decodeResult_specialSlot <= 1'h0;
      requestReg_bits_decodeResult_topUop <= 5'h0;
      requestReg_bits_decodeResult_popCount <= 1'h0;
      requestReg_bits_decodeResult_ffo <= 1'h0;
      requestReg_bits_decodeResult_average <= 1'h0;
      requestReg_bits_decodeResult_reverse <= 1'h0;
      requestReg_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      requestReg_bits_decodeResult_scheduler <= 1'h0;
      requestReg_bits_decodeResult_sReadVD <= 1'h0;
      requestReg_bits_decodeResult_vtype <= 1'h0;
      requestReg_bits_decodeResult_sWrite <= 1'h0;
      requestReg_bits_decodeResult_crossRead <= 1'h0;
      requestReg_bits_decodeResult_crossWrite <= 1'h0;
      requestReg_bits_decodeResult_maskUnit <= 1'h0;
      requestReg_bits_decodeResult_special <= 1'h0;
      requestReg_bits_decodeResult_saturate <= 1'h0;
      requestReg_bits_decodeResult_vwmacc <= 1'h0;
      requestReg_bits_decodeResult_readOnly <= 1'h0;
      requestReg_bits_decodeResult_maskSource <= 1'h0;
      requestReg_bits_decodeResult_maskDestination <= 1'h0;
      requestReg_bits_decodeResult_maskLogic <= 1'h0;
      requestReg_bits_decodeResult_uop <= 4'h0;
      requestReg_bits_decodeResult_iota <= 1'h0;
      requestReg_bits_decodeResult_mv <= 1'h0;
      requestReg_bits_decodeResult_extend <= 1'h0;
      requestReg_bits_decodeResult_unOrderWrite <= 1'h0;
      requestReg_bits_decodeResult_compress <= 1'h0;
      requestReg_bits_decodeResult_gather16 <= 1'h0;
      requestReg_bits_decodeResult_gather <= 1'h0;
      requestReg_bits_decodeResult_slid <= 1'h0;
      requestReg_bits_decodeResult_targetRd <= 1'h0;
      requestReg_bits_decodeResult_widenReduce <= 1'h0;
      requestReg_bits_decodeResult_red <= 1'h0;
      requestReg_bits_decodeResult_nr <= 1'h0;
      requestReg_bits_decodeResult_itype <= 1'h0;
      requestReg_bits_decodeResult_unsigned1 <= 1'h0;
      requestReg_bits_decodeResult_unsigned0 <= 1'h0;
      requestReg_bits_decodeResult_other <= 1'h0;
      requestReg_bits_decodeResult_multiCycle <= 1'h0;
      requestReg_bits_decodeResult_divider <= 1'h0;
      requestReg_bits_decodeResult_multiplier <= 1'h0;
      requestReg_bits_decodeResult_shift <= 1'h0;
      requestReg_bits_decodeResult_adder <= 1'h0;
      requestReg_bits_decodeResult_logic <= 1'h0;
      requestReg_bits_instructionIndex <= 3'h0;
      requestReg_bits_vdIsV0 <= 1'h0;
      requestReg_bits_writeByte <= 12'h0;
      slots_0_record_instructionIndex <= 3'h7;
      slots_0_record_isLoadStore <= 1'h1;
      slots_0_record_maskType <= 1'h1;
      slots_0_state_wLast <= 1'h1;
      slots_0_state_idle <= 1'h1;
      slots_0_state_wMaskUnitLast <= 1'h1;
      slots_0_state_wVRFWrite <= 1'h1;
      slots_0_state_sCommit <= 1'h1;
      slots_0_endTag_0 <= 1'h1;
      slots_0_endTag_1 <= 1'h1;
      slots_0_endTag_2 <= 1'h1;
      slots_0_endTag_3 <= 1'h1;
      slots_0_endTag_4 <= 1'h1;
      slots_0_endTag_5 <= 1'h1;
      slots_0_endTag_6 <= 1'h1;
      slots_0_endTag_7 <= 1'h1;
      slots_0_endTag_8 <= 1'h1;
      slots_0_endTag_9 <= 1'h1;
      slots_0_endTag_10 <= 1'h1;
      slots_0_endTag_11 <= 1'h1;
      slots_0_endTag_12 <= 1'h1;
      slots_0_endTag_13 <= 1'h1;
      slots_0_endTag_14 <= 1'h1;
      slots_0_endTag_15 <= 1'h1;
      slots_0_endTag_16 <= 1'h1;
      slots_0_vxsat <= 1'h1;
      slots_1_record_instructionIndex <= 3'h7;
      slots_1_record_isLoadStore <= 1'h1;
      slots_1_record_maskType <= 1'h1;
      slots_1_state_wLast <= 1'h1;
      slots_1_state_idle <= 1'h1;
      slots_1_state_wMaskUnitLast <= 1'h1;
      slots_1_state_wVRFWrite <= 1'h1;
      slots_1_state_sCommit <= 1'h1;
      slots_1_endTag_0 <= 1'h1;
      slots_1_endTag_1 <= 1'h1;
      slots_1_endTag_2 <= 1'h1;
      slots_1_endTag_3 <= 1'h1;
      slots_1_endTag_4 <= 1'h1;
      slots_1_endTag_5 <= 1'h1;
      slots_1_endTag_6 <= 1'h1;
      slots_1_endTag_7 <= 1'h1;
      slots_1_endTag_8 <= 1'h1;
      slots_1_endTag_9 <= 1'h1;
      slots_1_endTag_10 <= 1'h1;
      slots_1_endTag_11 <= 1'h1;
      slots_1_endTag_12 <= 1'h1;
      slots_1_endTag_13 <= 1'h1;
      slots_1_endTag_14 <= 1'h1;
      slots_1_endTag_15 <= 1'h1;
      slots_1_endTag_16 <= 1'h1;
      slots_1_vxsat <= 1'h1;
      slots_2_record_instructionIndex <= 3'h7;
      slots_2_record_isLoadStore <= 1'h1;
      slots_2_record_maskType <= 1'h1;
      slots_2_state_wLast <= 1'h1;
      slots_2_state_idle <= 1'h1;
      slots_2_state_wMaskUnitLast <= 1'h1;
      slots_2_state_wVRFWrite <= 1'h1;
      slots_2_state_sCommit <= 1'h1;
      slots_2_endTag_0 <= 1'h1;
      slots_2_endTag_1 <= 1'h1;
      slots_2_endTag_2 <= 1'h1;
      slots_2_endTag_3 <= 1'h1;
      slots_2_endTag_4 <= 1'h1;
      slots_2_endTag_5 <= 1'h1;
      slots_2_endTag_6 <= 1'h1;
      slots_2_endTag_7 <= 1'h1;
      slots_2_endTag_8 <= 1'h1;
      slots_2_endTag_9 <= 1'h1;
      slots_2_endTag_10 <= 1'h1;
      slots_2_endTag_11 <= 1'h1;
      slots_2_endTag_12 <= 1'h1;
      slots_2_endTag_13 <= 1'h1;
      slots_2_endTag_14 <= 1'h1;
      slots_2_endTag_15 <= 1'h1;
      slots_2_endTag_16 <= 1'h1;
      slots_2_vxsat <= 1'h1;
      slots_3_record_instructionIndex <= 3'h7;
      slots_3_record_isLoadStore <= 1'h1;
      slots_3_record_maskType <= 1'h1;
      slots_3_state_wLast <= 1'h1;
      slots_3_state_idle <= 1'h1;
      slots_3_state_wMaskUnitLast <= 1'h1;
      slots_3_state_wVRFWrite <= 1'h1;
      slots_3_state_sCommit <= 1'h1;
      slots_3_endTag_0 <= 1'h1;
      slots_3_endTag_1 <= 1'h1;
      slots_3_endTag_2 <= 1'h1;
      slots_3_endTag_3 <= 1'h1;
      slots_3_endTag_4 <= 1'h1;
      slots_3_endTag_5 <= 1'h1;
      slots_3_endTag_6 <= 1'h1;
      slots_3_endTag_7 <= 1'h1;
      slots_3_endTag_8 <= 1'h1;
      slots_3_endTag_9 <= 1'h1;
      slots_3_endTag_10 <= 1'h1;
      slots_3_endTag_11 <= 1'h1;
      slots_3_endTag_12 <= 1'h1;
      slots_3_endTag_13 <= 1'h1;
      slots_3_endTag_14 <= 1'h1;
      slots_3_endTag_15 <= 1'h1;
      slots_3_endTag_16 <= 1'h1;
      slots_3_vxsat <= 1'h1;
      slots_writeRD <= 1'h0;
      slots_float <= 1'h0;
      slots_vd <= 5'h0;
      releasePipe_pipe_v <= 1'h0;
      tokenCheck_counter <= 3'h0;
      shifterReg_0_valid <= 1'h0;
      shifterReg_0_bits_instructionIndex <= 3'h0;
      shifterReg_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_0_bits_decodeResult_float <= 1'h0;
      shifterReg_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_0_bits_decodeResult_average <= 1'h0;
      shifterReg_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_0_bits_decodeResult_special <= 1'h0;
      shifterReg_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_0_bits_decodeResult_red <= 1'h0;
      shifterReg_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_0_bits_decodeResult_other <= 1'h0;
      shifterReg_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_0_bits_loadStore <= 1'h0;
      shifterReg_0_bits_issueInst <= 1'h0;
      shifterReg_0_bits_store <= 1'h0;
      shifterReg_0_bits_special <= 1'h0;
      shifterReg_0_bits_lsWholeReg <= 1'h0;
      shifterReg_0_bits_vs1 <= 5'h0;
      shifterReg_0_bits_vs2 <= 5'h0;
      shifterReg_0_bits_vd <= 5'h0;
      shifterReg_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_0_bits_mask <= 1'h0;
      shifterReg_0_bits_segment <= 3'h0;
      shifterReg_0_bits_readFromScalar <= 32'h0;
      shifterReg_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_1 <= 1'h0;
      tokenCheck_counter_1 <= 3'h0;
      shifterReg_1_0_valid <= 1'h0;
      shifterReg_1_0_bits_instructionIndex <= 3'h0;
      shifterReg_1_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_1_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_1_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_1_0_bits_decodeResult_float <= 1'h0;
      shifterReg_1_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_1_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_1_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_1_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_1_0_bits_decodeResult_average <= 1'h0;
      shifterReg_1_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_1_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_1_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_1_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_1_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_1_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_1_0_bits_decodeResult_special <= 1'h0;
      shifterReg_1_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_1_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_1_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_1_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_1_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_1_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_1_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_1_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_1_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_1_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_1_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_1_0_bits_decodeResult_red <= 1'h0;
      shifterReg_1_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_1_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_other <= 1'h0;
      shifterReg_1_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_1_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_1_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_1_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_1_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_1_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_1_0_bits_loadStore <= 1'h0;
      shifterReg_1_0_bits_issueInst <= 1'h0;
      shifterReg_1_0_bits_store <= 1'h0;
      shifterReg_1_0_bits_special <= 1'h0;
      shifterReg_1_0_bits_lsWholeReg <= 1'h0;
      shifterReg_1_0_bits_vs1 <= 5'h0;
      shifterReg_1_0_bits_vs2 <= 5'h0;
      shifterReg_1_0_bits_vd <= 5'h0;
      shifterReg_1_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_1_0_bits_mask <= 1'h0;
      shifterReg_1_0_bits_segment <= 3'h0;
      shifterReg_1_0_bits_readFromScalar <= 32'h0;
      shifterReg_1_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_1_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_1_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_1_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_1_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_1_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_1_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_2 <= 1'h0;
      tokenCheck_counter_2 <= 3'h0;
      shifterReg_2_0_valid <= 1'h0;
      shifterReg_2_0_bits_instructionIndex <= 3'h0;
      shifterReg_2_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_2_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_2_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_2_0_bits_decodeResult_float <= 1'h0;
      shifterReg_2_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_2_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_2_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_2_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_2_0_bits_decodeResult_average <= 1'h0;
      shifterReg_2_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_2_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_2_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_2_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_2_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_2_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_2_0_bits_decodeResult_special <= 1'h0;
      shifterReg_2_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_2_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_2_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_2_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_2_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_2_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_2_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_2_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_2_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_2_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_2_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_2_0_bits_decodeResult_red <= 1'h0;
      shifterReg_2_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_2_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_other <= 1'h0;
      shifterReg_2_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_2_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_2_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_2_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_2_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_2_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_2_0_bits_loadStore <= 1'h0;
      shifterReg_2_0_bits_issueInst <= 1'h0;
      shifterReg_2_0_bits_store <= 1'h0;
      shifterReg_2_0_bits_special <= 1'h0;
      shifterReg_2_0_bits_lsWholeReg <= 1'h0;
      shifterReg_2_0_bits_vs1 <= 5'h0;
      shifterReg_2_0_bits_vs2 <= 5'h0;
      shifterReg_2_0_bits_vd <= 5'h0;
      shifterReg_2_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_2_0_bits_mask <= 1'h0;
      shifterReg_2_0_bits_segment <= 3'h0;
      shifterReg_2_0_bits_readFromScalar <= 32'h0;
      shifterReg_2_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_2_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_2_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_2_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_2_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_2_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_2_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_3 <= 1'h0;
      tokenCheck_counter_3 <= 3'h0;
      shifterReg_3_0_valid <= 1'h0;
      shifterReg_3_0_bits_instructionIndex <= 3'h0;
      shifterReg_3_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_3_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_3_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_3_0_bits_decodeResult_float <= 1'h0;
      shifterReg_3_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_3_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_3_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_3_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_3_0_bits_decodeResult_average <= 1'h0;
      shifterReg_3_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_3_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_3_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_3_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_3_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_3_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_3_0_bits_decodeResult_special <= 1'h0;
      shifterReg_3_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_3_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_3_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_3_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_3_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_3_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_3_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_3_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_3_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_3_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_3_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_3_0_bits_decodeResult_red <= 1'h0;
      shifterReg_3_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_3_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_other <= 1'h0;
      shifterReg_3_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_3_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_3_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_3_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_3_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_3_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_3_0_bits_loadStore <= 1'h0;
      shifterReg_3_0_bits_issueInst <= 1'h0;
      shifterReg_3_0_bits_store <= 1'h0;
      shifterReg_3_0_bits_special <= 1'h0;
      shifterReg_3_0_bits_lsWholeReg <= 1'h0;
      shifterReg_3_0_bits_vs1 <= 5'h0;
      shifterReg_3_0_bits_vs2 <= 5'h0;
      shifterReg_3_0_bits_vd <= 5'h0;
      shifterReg_3_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_3_0_bits_mask <= 1'h0;
      shifterReg_3_0_bits_segment <= 3'h0;
      shifterReg_3_0_bits_readFromScalar <= 32'h0;
      shifterReg_3_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_3_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_3_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_3_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_3_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_3_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_3_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_4 <= 1'h0;
      tokenCheck_counter_4 <= 3'h0;
      shifterReg_4_0_valid <= 1'h0;
      shifterReg_4_0_bits_instructionIndex <= 3'h0;
      shifterReg_4_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_4_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_4_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_4_0_bits_decodeResult_float <= 1'h0;
      shifterReg_4_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_4_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_4_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_4_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_4_0_bits_decodeResult_average <= 1'h0;
      shifterReg_4_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_4_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_4_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_4_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_4_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_4_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_4_0_bits_decodeResult_special <= 1'h0;
      shifterReg_4_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_4_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_4_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_4_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_4_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_4_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_4_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_4_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_4_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_4_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_4_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_4_0_bits_decodeResult_red <= 1'h0;
      shifterReg_4_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_4_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_other <= 1'h0;
      shifterReg_4_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_4_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_4_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_4_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_4_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_4_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_4_0_bits_loadStore <= 1'h0;
      shifterReg_4_0_bits_issueInst <= 1'h0;
      shifterReg_4_0_bits_store <= 1'h0;
      shifterReg_4_0_bits_special <= 1'h0;
      shifterReg_4_0_bits_lsWholeReg <= 1'h0;
      shifterReg_4_0_bits_vs1 <= 5'h0;
      shifterReg_4_0_bits_vs2 <= 5'h0;
      shifterReg_4_0_bits_vd <= 5'h0;
      shifterReg_4_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_4_0_bits_mask <= 1'h0;
      shifterReg_4_0_bits_segment <= 3'h0;
      shifterReg_4_0_bits_readFromScalar <= 32'h0;
      shifterReg_4_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_4_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_4_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_4_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_4_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_4_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_4_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_5 <= 1'h0;
      tokenCheck_counter_5 <= 3'h0;
      shifterReg_5_0_valid <= 1'h0;
      shifterReg_5_0_bits_instructionIndex <= 3'h0;
      shifterReg_5_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_5_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_5_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_5_0_bits_decodeResult_float <= 1'h0;
      shifterReg_5_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_5_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_5_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_5_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_5_0_bits_decodeResult_average <= 1'h0;
      shifterReg_5_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_5_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_5_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_5_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_5_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_5_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_5_0_bits_decodeResult_special <= 1'h0;
      shifterReg_5_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_5_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_5_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_5_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_5_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_5_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_5_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_5_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_5_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_5_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_5_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_5_0_bits_decodeResult_red <= 1'h0;
      shifterReg_5_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_5_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_other <= 1'h0;
      shifterReg_5_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_5_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_5_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_5_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_5_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_5_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_5_0_bits_loadStore <= 1'h0;
      shifterReg_5_0_bits_issueInst <= 1'h0;
      shifterReg_5_0_bits_store <= 1'h0;
      shifterReg_5_0_bits_special <= 1'h0;
      shifterReg_5_0_bits_lsWholeReg <= 1'h0;
      shifterReg_5_0_bits_vs1 <= 5'h0;
      shifterReg_5_0_bits_vs2 <= 5'h0;
      shifterReg_5_0_bits_vd <= 5'h0;
      shifterReg_5_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_5_0_bits_mask <= 1'h0;
      shifterReg_5_0_bits_segment <= 3'h0;
      shifterReg_5_0_bits_readFromScalar <= 32'h0;
      shifterReg_5_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_5_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_5_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_5_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_5_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_5_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_5_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_6 <= 1'h0;
      tokenCheck_counter_6 <= 3'h0;
      shifterReg_6_0_valid <= 1'h0;
      shifterReg_6_0_bits_instructionIndex <= 3'h0;
      shifterReg_6_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_6_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_6_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_6_0_bits_decodeResult_float <= 1'h0;
      shifterReg_6_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_6_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_6_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_6_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_6_0_bits_decodeResult_average <= 1'h0;
      shifterReg_6_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_6_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_6_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_6_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_6_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_6_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_6_0_bits_decodeResult_special <= 1'h0;
      shifterReg_6_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_6_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_6_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_6_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_6_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_6_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_6_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_6_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_6_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_6_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_6_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_6_0_bits_decodeResult_red <= 1'h0;
      shifterReg_6_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_6_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_other <= 1'h0;
      shifterReg_6_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_6_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_6_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_6_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_6_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_6_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_6_0_bits_loadStore <= 1'h0;
      shifterReg_6_0_bits_issueInst <= 1'h0;
      shifterReg_6_0_bits_store <= 1'h0;
      shifterReg_6_0_bits_special <= 1'h0;
      shifterReg_6_0_bits_lsWholeReg <= 1'h0;
      shifterReg_6_0_bits_vs1 <= 5'h0;
      shifterReg_6_0_bits_vs2 <= 5'h0;
      shifterReg_6_0_bits_vd <= 5'h0;
      shifterReg_6_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_6_0_bits_mask <= 1'h0;
      shifterReg_6_0_bits_segment <= 3'h0;
      shifterReg_6_0_bits_readFromScalar <= 32'h0;
      shifterReg_6_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_6_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_6_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_6_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_6_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_6_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_6_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_7 <= 1'h0;
      tokenCheck_counter_7 <= 3'h0;
      shifterReg_7_0_valid <= 1'h0;
      shifterReg_7_0_bits_instructionIndex <= 3'h0;
      shifterReg_7_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_7_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_7_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_7_0_bits_decodeResult_float <= 1'h0;
      shifterReg_7_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_7_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_7_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_7_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_7_0_bits_decodeResult_average <= 1'h0;
      shifterReg_7_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_7_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_7_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_7_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_7_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_7_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_7_0_bits_decodeResult_special <= 1'h0;
      shifterReg_7_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_7_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_7_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_7_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_7_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_7_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_7_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_7_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_7_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_7_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_7_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_7_0_bits_decodeResult_red <= 1'h0;
      shifterReg_7_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_7_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_other <= 1'h0;
      shifterReg_7_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_7_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_7_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_7_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_7_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_7_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_7_0_bits_loadStore <= 1'h0;
      shifterReg_7_0_bits_issueInst <= 1'h0;
      shifterReg_7_0_bits_store <= 1'h0;
      shifterReg_7_0_bits_special <= 1'h0;
      shifterReg_7_0_bits_lsWholeReg <= 1'h0;
      shifterReg_7_0_bits_vs1 <= 5'h0;
      shifterReg_7_0_bits_vs2 <= 5'h0;
      shifterReg_7_0_bits_vd <= 5'h0;
      shifterReg_7_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_7_0_bits_mask <= 1'h0;
      shifterReg_7_0_bits_segment <= 3'h0;
      shifterReg_7_0_bits_readFromScalar <= 32'h0;
      shifterReg_7_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_7_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_7_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_7_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_7_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_7_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_7_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_8 <= 1'h0;
      tokenCheck_counter_8 <= 3'h0;
      shifterReg_8_0_valid <= 1'h0;
      shifterReg_8_0_bits_instructionIndex <= 3'h0;
      shifterReg_8_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_8_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_8_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_8_0_bits_decodeResult_float <= 1'h0;
      shifterReg_8_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_8_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_8_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_8_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_8_0_bits_decodeResult_average <= 1'h0;
      shifterReg_8_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_8_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_8_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_8_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_8_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_8_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_8_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_8_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_8_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_8_0_bits_decodeResult_special <= 1'h0;
      shifterReg_8_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_8_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_8_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_8_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_8_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_8_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_8_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_8_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_8_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_8_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_8_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_8_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_8_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_8_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_8_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_8_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_8_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_8_0_bits_decodeResult_red <= 1'h0;
      shifterReg_8_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_8_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_8_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_8_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_8_0_bits_decodeResult_other <= 1'h0;
      shifterReg_8_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_8_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_8_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_8_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_8_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_8_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_8_0_bits_loadStore <= 1'h0;
      shifterReg_8_0_bits_issueInst <= 1'h0;
      shifterReg_8_0_bits_store <= 1'h0;
      shifterReg_8_0_bits_special <= 1'h0;
      shifterReg_8_0_bits_lsWholeReg <= 1'h0;
      shifterReg_8_0_bits_vs1 <= 5'h0;
      shifterReg_8_0_bits_vs2 <= 5'h0;
      shifterReg_8_0_bits_vd <= 5'h0;
      shifterReg_8_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_8_0_bits_mask <= 1'h0;
      shifterReg_8_0_bits_segment <= 3'h0;
      shifterReg_8_0_bits_readFromScalar <= 32'h0;
      shifterReg_8_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_8_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_8_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_8_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_8_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_8_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_8_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_9 <= 1'h0;
      tokenCheck_counter_9 <= 3'h0;
      shifterReg_9_0_valid <= 1'h0;
      shifterReg_9_0_bits_instructionIndex <= 3'h0;
      shifterReg_9_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_9_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_9_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_9_0_bits_decodeResult_float <= 1'h0;
      shifterReg_9_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_9_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_9_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_9_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_9_0_bits_decodeResult_average <= 1'h0;
      shifterReg_9_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_9_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_9_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_9_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_9_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_9_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_9_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_9_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_9_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_9_0_bits_decodeResult_special <= 1'h0;
      shifterReg_9_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_9_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_9_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_9_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_9_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_9_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_9_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_9_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_9_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_9_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_9_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_9_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_9_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_9_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_9_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_9_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_9_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_9_0_bits_decodeResult_red <= 1'h0;
      shifterReg_9_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_9_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_9_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_9_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_9_0_bits_decodeResult_other <= 1'h0;
      shifterReg_9_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_9_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_9_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_9_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_9_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_9_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_9_0_bits_loadStore <= 1'h0;
      shifterReg_9_0_bits_issueInst <= 1'h0;
      shifterReg_9_0_bits_store <= 1'h0;
      shifterReg_9_0_bits_special <= 1'h0;
      shifterReg_9_0_bits_lsWholeReg <= 1'h0;
      shifterReg_9_0_bits_vs1 <= 5'h0;
      shifterReg_9_0_bits_vs2 <= 5'h0;
      shifterReg_9_0_bits_vd <= 5'h0;
      shifterReg_9_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_9_0_bits_mask <= 1'h0;
      shifterReg_9_0_bits_segment <= 3'h0;
      shifterReg_9_0_bits_readFromScalar <= 32'h0;
      shifterReg_9_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_9_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_9_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_9_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_9_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_9_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_9_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_10 <= 1'h0;
      tokenCheck_counter_10 <= 3'h0;
      shifterReg_10_0_valid <= 1'h0;
      shifterReg_10_0_bits_instructionIndex <= 3'h0;
      shifterReg_10_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_10_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_10_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_10_0_bits_decodeResult_float <= 1'h0;
      shifterReg_10_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_10_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_10_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_10_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_10_0_bits_decodeResult_average <= 1'h0;
      shifterReg_10_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_10_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_10_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_10_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_10_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_10_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_10_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_10_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_10_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_10_0_bits_decodeResult_special <= 1'h0;
      shifterReg_10_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_10_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_10_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_10_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_10_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_10_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_10_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_10_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_10_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_10_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_10_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_10_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_10_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_10_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_10_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_10_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_10_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_10_0_bits_decodeResult_red <= 1'h0;
      shifterReg_10_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_10_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_10_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_10_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_10_0_bits_decodeResult_other <= 1'h0;
      shifterReg_10_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_10_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_10_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_10_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_10_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_10_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_10_0_bits_loadStore <= 1'h0;
      shifterReg_10_0_bits_issueInst <= 1'h0;
      shifterReg_10_0_bits_store <= 1'h0;
      shifterReg_10_0_bits_special <= 1'h0;
      shifterReg_10_0_bits_lsWholeReg <= 1'h0;
      shifterReg_10_0_bits_vs1 <= 5'h0;
      shifterReg_10_0_bits_vs2 <= 5'h0;
      shifterReg_10_0_bits_vd <= 5'h0;
      shifterReg_10_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_10_0_bits_mask <= 1'h0;
      shifterReg_10_0_bits_segment <= 3'h0;
      shifterReg_10_0_bits_readFromScalar <= 32'h0;
      shifterReg_10_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_10_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_10_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_10_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_10_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_10_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_10_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_11 <= 1'h0;
      tokenCheck_counter_11 <= 3'h0;
      shifterReg_11_0_valid <= 1'h0;
      shifterReg_11_0_bits_instructionIndex <= 3'h0;
      shifterReg_11_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_11_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_11_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_11_0_bits_decodeResult_float <= 1'h0;
      shifterReg_11_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_11_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_11_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_11_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_11_0_bits_decodeResult_average <= 1'h0;
      shifterReg_11_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_11_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_11_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_11_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_11_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_11_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_11_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_11_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_11_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_11_0_bits_decodeResult_special <= 1'h0;
      shifterReg_11_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_11_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_11_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_11_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_11_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_11_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_11_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_11_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_11_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_11_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_11_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_11_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_11_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_11_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_11_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_11_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_11_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_11_0_bits_decodeResult_red <= 1'h0;
      shifterReg_11_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_11_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_11_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_11_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_11_0_bits_decodeResult_other <= 1'h0;
      shifterReg_11_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_11_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_11_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_11_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_11_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_11_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_11_0_bits_loadStore <= 1'h0;
      shifterReg_11_0_bits_issueInst <= 1'h0;
      shifterReg_11_0_bits_store <= 1'h0;
      shifterReg_11_0_bits_special <= 1'h0;
      shifterReg_11_0_bits_lsWholeReg <= 1'h0;
      shifterReg_11_0_bits_vs1 <= 5'h0;
      shifterReg_11_0_bits_vs2 <= 5'h0;
      shifterReg_11_0_bits_vd <= 5'h0;
      shifterReg_11_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_11_0_bits_mask <= 1'h0;
      shifterReg_11_0_bits_segment <= 3'h0;
      shifterReg_11_0_bits_readFromScalar <= 32'h0;
      shifterReg_11_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_11_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_11_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_11_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_11_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_11_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_11_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_12 <= 1'h0;
      tokenCheck_counter_12 <= 3'h0;
      shifterReg_12_0_valid <= 1'h0;
      shifterReg_12_0_bits_instructionIndex <= 3'h0;
      shifterReg_12_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_12_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_12_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_12_0_bits_decodeResult_float <= 1'h0;
      shifterReg_12_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_12_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_12_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_12_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_12_0_bits_decodeResult_average <= 1'h0;
      shifterReg_12_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_12_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_12_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_12_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_12_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_12_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_12_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_12_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_12_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_12_0_bits_decodeResult_special <= 1'h0;
      shifterReg_12_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_12_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_12_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_12_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_12_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_12_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_12_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_12_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_12_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_12_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_12_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_12_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_12_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_12_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_12_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_12_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_12_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_12_0_bits_decodeResult_red <= 1'h0;
      shifterReg_12_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_12_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_12_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_12_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_12_0_bits_decodeResult_other <= 1'h0;
      shifterReg_12_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_12_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_12_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_12_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_12_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_12_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_12_0_bits_loadStore <= 1'h0;
      shifterReg_12_0_bits_issueInst <= 1'h0;
      shifterReg_12_0_bits_store <= 1'h0;
      shifterReg_12_0_bits_special <= 1'h0;
      shifterReg_12_0_bits_lsWholeReg <= 1'h0;
      shifterReg_12_0_bits_vs1 <= 5'h0;
      shifterReg_12_0_bits_vs2 <= 5'h0;
      shifterReg_12_0_bits_vd <= 5'h0;
      shifterReg_12_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_12_0_bits_mask <= 1'h0;
      shifterReg_12_0_bits_segment <= 3'h0;
      shifterReg_12_0_bits_readFromScalar <= 32'h0;
      shifterReg_12_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_12_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_12_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_12_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_12_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_12_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_12_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_13 <= 1'h0;
      tokenCheck_counter_13 <= 3'h0;
      shifterReg_13_0_valid <= 1'h0;
      shifterReg_13_0_bits_instructionIndex <= 3'h0;
      shifterReg_13_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_13_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_13_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_13_0_bits_decodeResult_float <= 1'h0;
      shifterReg_13_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_13_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_13_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_13_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_13_0_bits_decodeResult_average <= 1'h0;
      shifterReg_13_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_13_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_13_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_13_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_13_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_13_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_13_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_13_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_13_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_13_0_bits_decodeResult_special <= 1'h0;
      shifterReg_13_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_13_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_13_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_13_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_13_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_13_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_13_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_13_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_13_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_13_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_13_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_13_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_13_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_13_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_13_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_13_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_13_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_13_0_bits_decodeResult_red <= 1'h0;
      shifterReg_13_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_13_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_13_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_13_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_13_0_bits_decodeResult_other <= 1'h0;
      shifterReg_13_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_13_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_13_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_13_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_13_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_13_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_13_0_bits_loadStore <= 1'h0;
      shifterReg_13_0_bits_issueInst <= 1'h0;
      shifterReg_13_0_bits_store <= 1'h0;
      shifterReg_13_0_bits_special <= 1'h0;
      shifterReg_13_0_bits_lsWholeReg <= 1'h0;
      shifterReg_13_0_bits_vs1 <= 5'h0;
      shifterReg_13_0_bits_vs2 <= 5'h0;
      shifterReg_13_0_bits_vd <= 5'h0;
      shifterReg_13_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_13_0_bits_mask <= 1'h0;
      shifterReg_13_0_bits_segment <= 3'h0;
      shifterReg_13_0_bits_readFromScalar <= 32'h0;
      shifterReg_13_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_13_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_13_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_13_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_13_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_13_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_13_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_14 <= 1'h0;
      tokenCheck_counter_14 <= 3'h0;
      shifterReg_14_0_valid <= 1'h0;
      shifterReg_14_0_bits_instructionIndex <= 3'h0;
      shifterReg_14_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_14_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_14_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_14_0_bits_decodeResult_float <= 1'h0;
      shifterReg_14_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_14_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_14_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_14_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_14_0_bits_decodeResult_average <= 1'h0;
      shifterReg_14_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_14_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_14_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_14_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_14_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_14_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_14_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_14_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_14_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_14_0_bits_decodeResult_special <= 1'h0;
      shifterReg_14_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_14_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_14_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_14_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_14_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_14_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_14_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_14_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_14_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_14_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_14_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_14_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_14_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_14_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_14_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_14_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_14_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_14_0_bits_decodeResult_red <= 1'h0;
      shifterReg_14_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_14_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_14_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_14_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_14_0_bits_decodeResult_other <= 1'h0;
      shifterReg_14_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_14_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_14_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_14_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_14_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_14_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_14_0_bits_loadStore <= 1'h0;
      shifterReg_14_0_bits_issueInst <= 1'h0;
      shifterReg_14_0_bits_store <= 1'h0;
      shifterReg_14_0_bits_special <= 1'h0;
      shifterReg_14_0_bits_lsWholeReg <= 1'h0;
      shifterReg_14_0_bits_vs1 <= 5'h0;
      shifterReg_14_0_bits_vs2 <= 5'h0;
      shifterReg_14_0_bits_vd <= 5'h0;
      shifterReg_14_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_14_0_bits_mask <= 1'h0;
      shifterReg_14_0_bits_segment <= 3'h0;
      shifterReg_14_0_bits_readFromScalar <= 32'h0;
      shifterReg_14_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_14_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_14_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_14_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_14_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_14_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_14_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_15 <= 1'h0;
      tokenCheck_counter_15 <= 3'h0;
      shifterReg_15_0_valid <= 1'h0;
      shifterReg_15_0_bits_instructionIndex <= 3'h0;
      shifterReg_15_0_bits_decodeResult_orderReduce <= 1'h0;
      shifterReg_15_0_bits_decodeResult_floatMul <= 1'h0;
      shifterReg_15_0_bits_decodeResult_fpExecutionType <= 2'h0;
      shifterReg_15_0_bits_decodeResult_float <= 1'h0;
      shifterReg_15_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_15_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_15_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_15_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_15_0_bits_decodeResult_average <= 1'h0;
      shifterReg_15_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_15_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_15_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_15_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_15_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_15_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_15_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_15_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_15_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_15_0_bits_decodeResult_special <= 1'h0;
      shifterReg_15_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_15_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_15_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_15_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_15_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_15_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_15_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_15_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_15_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_15_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_15_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_15_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_15_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_15_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_15_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_15_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_15_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_15_0_bits_decodeResult_red <= 1'h0;
      shifterReg_15_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_15_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_15_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_15_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_15_0_bits_decodeResult_other <= 1'h0;
      shifterReg_15_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_15_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_15_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_15_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_15_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_15_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_15_0_bits_loadStore <= 1'h0;
      shifterReg_15_0_bits_issueInst <= 1'h0;
      shifterReg_15_0_bits_store <= 1'h0;
      shifterReg_15_0_bits_special <= 1'h0;
      shifterReg_15_0_bits_lsWholeReg <= 1'h0;
      shifterReg_15_0_bits_vs1 <= 5'h0;
      shifterReg_15_0_bits_vs2 <= 5'h0;
      shifterReg_15_0_bits_vd <= 5'h0;
      shifterReg_15_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_15_0_bits_mask <= 1'h0;
      shifterReg_15_0_bits_segment <= 3'h0;
      shifterReg_15_0_bits_readFromScalar <= 32'h0;
      shifterReg_15_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_15_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_15_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_15_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_15_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_15_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_15_0_bits_csrInterface_vma <= 1'h0;
      sinkVec_releasePipe_pipe_v <= 1'h0;
      sinkVec_tokenCheck_counter <= 3'h0;
      sinkVec_shifterReg_0_valid <= 1'h0;
      sinkVec_shifterReg_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_1 <= 1'h0;
      sinkVec_tokenCheck_counter_1 <= 3'h0;
      sinkVec_shifterReg_1_0_valid <= 1'h0;
      sinkVec_shifterReg_1_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_1_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_1_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_1_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst <= 1'h0;
      accessDataValid_pipe_v <= 1'h0;
      accessDataValid_pipe_pipe_v <= 1'h0;
      shifterReg_16_0_valid <= 1'h0;
      shifterReg_16_0_bits <= 32'h0;
      accessDataValid_pipe_v_1 <= 1'h0;
      accessDataValid_pipe_pipe_v_1 <= 1'h0;
      shifterReg_17_0_valid <= 1'h0;
      shifterReg_17_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_2 <= 1'h0;
      sinkVec_tokenCheck_counter_2 <= 3'h0;
      sinkVec_shifterReg_2_0_valid <= 1'h0;
      sinkVec_shifterReg_2_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_2_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_2_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_2_0_bits_data <= 32'h0;
      sinkVec_shifterReg_2_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_3 <= 1'h0;
      sinkVec_tokenCheck_counter_3 <= 3'h0;
      sinkVec_shifterReg_3_0_valid <= 1'h0;
      sinkVec_shifterReg_3_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_3_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_3_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_3_0_bits_data <= 32'h0;
      sinkVec_shifterReg_3_0_bits_last <= 1'h0;
      sinkVec_shifterReg_3_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_1 <= 1'h0;
      view__writeRelease_0_pipe_v <= 1'h0;
      pipe_v <= 1'h0;
      instructionFinishedPipe_pipe_v <= 1'h0;
      pipe_v_1 <= 1'h0;
      pipe_pipe_v <= 1'h0;
      view__laneMaskSelect_0_pipe_v <= 1'h0;
      view__laneMaskSelect_0_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_0_pipe_v <= 1'h0;
      view__laneMaskSewSelect_0_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v <= 1'h0;
      maskLastPipe_pipe_v <= 1'h0;
      pipe_v_2 <= 1'h0;
      sinkVec_releasePipe_pipe_v_4 <= 1'h0;
      sinkVec_tokenCheck_counter_4 <= 3'h0;
      sinkVec_shifterReg_4_0_valid <= 1'h0;
      sinkVec_shifterReg_4_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_4_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_4_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_4_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_5 <= 1'h0;
      sinkVec_tokenCheck_counter_5 <= 3'h0;
      sinkVec_shifterReg_5_0_valid <= 1'h0;
      sinkVec_shifterReg_5_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_5_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_5_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_5_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_2 <= 1'h0;
      accessDataValid_pipe_v_2 <= 1'h0;
      accessDataValid_pipe_pipe_v_2 <= 1'h0;
      shifterReg_18_0_valid <= 1'h0;
      shifterReg_18_0_bits <= 32'h0;
      accessDataValid_pipe_v_3 <= 1'h0;
      accessDataValid_pipe_pipe_v_3 <= 1'h0;
      shifterReg_19_0_valid <= 1'h0;
      shifterReg_19_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_6 <= 1'h0;
      sinkVec_tokenCheck_counter_6 <= 3'h0;
      sinkVec_shifterReg_6_0_valid <= 1'h0;
      sinkVec_shifterReg_6_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_6_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_6_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_6_0_bits_data <= 32'h0;
      sinkVec_shifterReg_6_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_7 <= 1'h0;
      sinkVec_tokenCheck_counter_7 <= 3'h0;
      sinkVec_shifterReg_7_0_valid <= 1'h0;
      sinkVec_shifterReg_7_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_7_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_7_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_7_0_bits_data <= 32'h0;
      sinkVec_shifterReg_7_0_bits_last <= 1'h0;
      sinkVec_shifterReg_7_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_3 <= 1'h0;
      view__writeRelease_1_pipe_v <= 1'h0;
      pipe_v_3 <= 1'h0;
      instructionFinishedPipe_pipe_v_1 <= 1'h0;
      pipe_v_4 <= 1'h0;
      pipe_pipe_v_1 <= 1'h0;
      view__laneMaskSelect_1_pipe_v <= 1'h0;
      view__laneMaskSelect_1_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_1_pipe_v <= 1'h0;
      view__laneMaskSewSelect_1_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_1 <= 1'h0;
      maskLastPipe_pipe_v_1 <= 1'h0;
      pipe_v_5 <= 1'h0;
      sinkVec_releasePipe_pipe_v_8 <= 1'h0;
      sinkVec_tokenCheck_counter_8 <= 3'h0;
      sinkVec_shifterReg_8_0_valid <= 1'h0;
      sinkVec_shifterReg_8_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_8_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_8_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_8_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_9 <= 1'h0;
      sinkVec_tokenCheck_counter_9 <= 3'h0;
      sinkVec_shifterReg_9_0_valid <= 1'h0;
      sinkVec_shifterReg_9_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_9_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_9_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_9_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_4 <= 1'h0;
      accessDataValid_pipe_v_4 <= 1'h0;
      accessDataValid_pipe_pipe_v_4 <= 1'h0;
      shifterReg_20_0_valid <= 1'h0;
      shifterReg_20_0_bits <= 32'h0;
      accessDataValid_pipe_v_5 <= 1'h0;
      accessDataValid_pipe_pipe_v_5 <= 1'h0;
      shifterReg_21_0_valid <= 1'h0;
      shifterReg_21_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_10 <= 1'h0;
      sinkVec_tokenCheck_counter_10 <= 3'h0;
      sinkVec_shifterReg_10_0_valid <= 1'h0;
      sinkVec_shifterReg_10_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_10_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_10_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_10_0_bits_data <= 32'h0;
      sinkVec_shifterReg_10_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_11 <= 1'h0;
      sinkVec_tokenCheck_counter_11 <= 3'h0;
      sinkVec_shifterReg_11_0_valid <= 1'h0;
      sinkVec_shifterReg_11_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_11_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_11_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_11_0_bits_data <= 32'h0;
      sinkVec_shifterReg_11_0_bits_last <= 1'h0;
      sinkVec_shifterReg_11_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_5 <= 1'h0;
      view__writeRelease_2_pipe_v <= 1'h0;
      pipe_v_6 <= 1'h0;
      instructionFinishedPipe_pipe_v_2 <= 1'h0;
      pipe_v_7 <= 1'h0;
      pipe_pipe_v_2 <= 1'h0;
      view__laneMaskSelect_2_pipe_v <= 1'h0;
      view__laneMaskSelect_2_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_2_pipe_v <= 1'h0;
      view__laneMaskSewSelect_2_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_2 <= 1'h0;
      maskLastPipe_pipe_v_2 <= 1'h0;
      pipe_v_8 <= 1'h0;
      sinkVec_releasePipe_pipe_v_12 <= 1'h0;
      sinkVec_tokenCheck_counter_12 <= 3'h0;
      sinkVec_shifterReg_12_0_valid <= 1'h0;
      sinkVec_shifterReg_12_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_12_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_12_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_12_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_13 <= 1'h0;
      sinkVec_tokenCheck_counter_13 <= 3'h0;
      sinkVec_shifterReg_13_0_valid <= 1'h0;
      sinkVec_shifterReg_13_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_13_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_13_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_13_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_6 <= 1'h0;
      accessDataValid_pipe_v_6 <= 1'h0;
      accessDataValid_pipe_pipe_v_6 <= 1'h0;
      shifterReg_22_0_valid <= 1'h0;
      shifterReg_22_0_bits <= 32'h0;
      accessDataValid_pipe_v_7 <= 1'h0;
      accessDataValid_pipe_pipe_v_7 <= 1'h0;
      shifterReg_23_0_valid <= 1'h0;
      shifterReg_23_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_14 <= 1'h0;
      sinkVec_tokenCheck_counter_14 <= 3'h0;
      sinkVec_shifterReg_14_0_valid <= 1'h0;
      sinkVec_shifterReg_14_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_14_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_14_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_14_0_bits_data <= 32'h0;
      sinkVec_shifterReg_14_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_15 <= 1'h0;
      sinkVec_tokenCheck_counter_15 <= 3'h0;
      sinkVec_shifterReg_15_0_valid <= 1'h0;
      sinkVec_shifterReg_15_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_15_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_15_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_15_0_bits_data <= 32'h0;
      sinkVec_shifterReg_15_0_bits_last <= 1'h0;
      sinkVec_shifterReg_15_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_7 <= 1'h0;
      view__writeRelease_3_pipe_v <= 1'h0;
      pipe_v_9 <= 1'h0;
      instructionFinishedPipe_pipe_v_3 <= 1'h0;
      pipe_v_10 <= 1'h0;
      pipe_pipe_v_3 <= 1'h0;
      view__laneMaskSelect_3_pipe_v <= 1'h0;
      view__laneMaskSelect_3_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_3_pipe_v <= 1'h0;
      view__laneMaskSewSelect_3_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_3 <= 1'h0;
      maskLastPipe_pipe_v_3 <= 1'h0;
      pipe_v_11 <= 1'h0;
      sinkVec_releasePipe_pipe_v_16 <= 1'h0;
      sinkVec_tokenCheck_counter_16 <= 3'h0;
      sinkVec_shifterReg_16_0_valid <= 1'h0;
      sinkVec_shifterReg_16_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_16_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_16_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_16_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_17 <= 1'h0;
      sinkVec_tokenCheck_counter_17 <= 3'h0;
      sinkVec_shifterReg_17_0_valid <= 1'h0;
      sinkVec_shifterReg_17_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_17_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_17_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_17_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_8 <= 1'h0;
      accessDataValid_pipe_v_8 <= 1'h0;
      accessDataValid_pipe_pipe_v_8 <= 1'h0;
      shifterReg_24_0_valid <= 1'h0;
      shifterReg_24_0_bits <= 32'h0;
      accessDataValid_pipe_v_9 <= 1'h0;
      accessDataValid_pipe_pipe_v_9 <= 1'h0;
      shifterReg_25_0_valid <= 1'h0;
      shifterReg_25_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_18 <= 1'h0;
      sinkVec_tokenCheck_counter_18 <= 3'h0;
      sinkVec_shifterReg_18_0_valid <= 1'h0;
      sinkVec_shifterReg_18_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_18_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_18_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_18_0_bits_data <= 32'h0;
      sinkVec_shifterReg_18_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_19 <= 1'h0;
      sinkVec_tokenCheck_counter_19 <= 3'h0;
      sinkVec_shifterReg_19_0_valid <= 1'h0;
      sinkVec_shifterReg_19_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_19_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_19_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_19_0_bits_data <= 32'h0;
      sinkVec_shifterReg_19_0_bits_last <= 1'h0;
      sinkVec_shifterReg_19_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_9 <= 1'h0;
      view__writeRelease_4_pipe_v <= 1'h0;
      pipe_v_12 <= 1'h0;
      instructionFinishedPipe_pipe_v_4 <= 1'h0;
      pipe_v_13 <= 1'h0;
      pipe_pipe_v_4 <= 1'h0;
      view__laneMaskSelect_4_pipe_v <= 1'h0;
      view__laneMaskSelect_4_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_4_pipe_v <= 1'h0;
      view__laneMaskSewSelect_4_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_4 <= 1'h0;
      maskLastPipe_pipe_v_4 <= 1'h0;
      pipe_v_14 <= 1'h0;
      sinkVec_releasePipe_pipe_v_20 <= 1'h0;
      sinkVec_tokenCheck_counter_20 <= 3'h0;
      sinkVec_shifterReg_20_0_valid <= 1'h0;
      sinkVec_shifterReg_20_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_20_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_20_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_20_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_21 <= 1'h0;
      sinkVec_tokenCheck_counter_21 <= 3'h0;
      sinkVec_shifterReg_21_0_valid <= 1'h0;
      sinkVec_shifterReg_21_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_21_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_21_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_21_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_10 <= 1'h0;
      accessDataValid_pipe_v_10 <= 1'h0;
      accessDataValid_pipe_pipe_v_10 <= 1'h0;
      shifterReg_26_0_valid <= 1'h0;
      shifterReg_26_0_bits <= 32'h0;
      accessDataValid_pipe_v_11 <= 1'h0;
      accessDataValid_pipe_pipe_v_11 <= 1'h0;
      shifterReg_27_0_valid <= 1'h0;
      shifterReg_27_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_22 <= 1'h0;
      sinkVec_tokenCheck_counter_22 <= 3'h0;
      sinkVec_shifterReg_22_0_valid <= 1'h0;
      sinkVec_shifterReg_22_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_22_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_22_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_22_0_bits_data <= 32'h0;
      sinkVec_shifterReg_22_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_23 <= 1'h0;
      sinkVec_tokenCheck_counter_23 <= 3'h0;
      sinkVec_shifterReg_23_0_valid <= 1'h0;
      sinkVec_shifterReg_23_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_23_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_23_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_23_0_bits_data <= 32'h0;
      sinkVec_shifterReg_23_0_bits_last <= 1'h0;
      sinkVec_shifterReg_23_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_11 <= 1'h0;
      view__writeRelease_5_pipe_v <= 1'h0;
      pipe_v_15 <= 1'h0;
      instructionFinishedPipe_pipe_v_5 <= 1'h0;
      pipe_v_16 <= 1'h0;
      pipe_pipe_v_5 <= 1'h0;
      view__laneMaskSelect_5_pipe_v <= 1'h0;
      view__laneMaskSelect_5_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_5_pipe_v <= 1'h0;
      view__laneMaskSewSelect_5_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_5 <= 1'h0;
      maskLastPipe_pipe_v_5 <= 1'h0;
      pipe_v_17 <= 1'h0;
      sinkVec_releasePipe_pipe_v_24 <= 1'h0;
      sinkVec_tokenCheck_counter_24 <= 3'h0;
      sinkVec_shifterReg_24_0_valid <= 1'h0;
      sinkVec_shifterReg_24_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_24_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_24_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_24_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_25 <= 1'h0;
      sinkVec_tokenCheck_counter_25 <= 3'h0;
      sinkVec_shifterReg_25_0_valid <= 1'h0;
      sinkVec_shifterReg_25_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_25_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_25_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_25_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_12 <= 1'h0;
      accessDataValid_pipe_v_12 <= 1'h0;
      accessDataValid_pipe_pipe_v_12 <= 1'h0;
      shifterReg_28_0_valid <= 1'h0;
      shifterReg_28_0_bits <= 32'h0;
      accessDataValid_pipe_v_13 <= 1'h0;
      accessDataValid_pipe_pipe_v_13 <= 1'h0;
      shifterReg_29_0_valid <= 1'h0;
      shifterReg_29_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_26 <= 1'h0;
      sinkVec_tokenCheck_counter_26 <= 3'h0;
      sinkVec_shifterReg_26_0_valid <= 1'h0;
      sinkVec_shifterReg_26_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_26_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_26_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_26_0_bits_data <= 32'h0;
      sinkVec_shifterReg_26_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_27 <= 1'h0;
      sinkVec_tokenCheck_counter_27 <= 3'h0;
      sinkVec_shifterReg_27_0_valid <= 1'h0;
      sinkVec_shifterReg_27_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_27_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_27_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_27_0_bits_data <= 32'h0;
      sinkVec_shifterReg_27_0_bits_last <= 1'h0;
      sinkVec_shifterReg_27_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_13 <= 1'h0;
      view__writeRelease_6_pipe_v <= 1'h0;
      pipe_v_18 <= 1'h0;
      instructionFinishedPipe_pipe_v_6 <= 1'h0;
      pipe_v_19 <= 1'h0;
      pipe_pipe_v_6 <= 1'h0;
      view__laneMaskSelect_6_pipe_v <= 1'h0;
      view__laneMaskSelect_6_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_6_pipe_v <= 1'h0;
      view__laneMaskSewSelect_6_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_6 <= 1'h0;
      maskLastPipe_pipe_v_6 <= 1'h0;
      pipe_v_20 <= 1'h0;
      sinkVec_releasePipe_pipe_v_28 <= 1'h0;
      sinkVec_tokenCheck_counter_28 <= 3'h0;
      sinkVec_shifterReg_28_0_valid <= 1'h0;
      sinkVec_shifterReg_28_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_28_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_28_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_28_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_29 <= 1'h0;
      sinkVec_tokenCheck_counter_29 <= 3'h0;
      sinkVec_shifterReg_29_0_valid <= 1'h0;
      sinkVec_shifterReg_29_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_29_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_29_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_29_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_14 <= 1'h0;
      accessDataValid_pipe_v_14 <= 1'h0;
      accessDataValid_pipe_pipe_v_14 <= 1'h0;
      shifterReg_30_0_valid <= 1'h0;
      shifterReg_30_0_bits <= 32'h0;
      accessDataValid_pipe_v_15 <= 1'h0;
      accessDataValid_pipe_pipe_v_15 <= 1'h0;
      shifterReg_31_0_valid <= 1'h0;
      shifterReg_31_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_30 <= 1'h0;
      sinkVec_tokenCheck_counter_30 <= 3'h0;
      sinkVec_shifterReg_30_0_valid <= 1'h0;
      sinkVec_shifterReg_30_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_30_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_30_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_30_0_bits_data <= 32'h0;
      sinkVec_shifterReg_30_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_31 <= 1'h0;
      sinkVec_tokenCheck_counter_31 <= 3'h0;
      sinkVec_shifterReg_31_0_valid <= 1'h0;
      sinkVec_shifterReg_31_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_31_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_31_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_31_0_bits_data <= 32'h0;
      sinkVec_shifterReg_31_0_bits_last <= 1'h0;
      sinkVec_shifterReg_31_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_15 <= 1'h0;
      view__writeRelease_7_pipe_v <= 1'h0;
      pipe_v_21 <= 1'h0;
      instructionFinishedPipe_pipe_v_7 <= 1'h0;
      pipe_v_22 <= 1'h0;
      pipe_pipe_v_7 <= 1'h0;
      view__laneMaskSelect_7_pipe_v <= 1'h0;
      view__laneMaskSelect_7_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_7_pipe_v <= 1'h0;
      view__laneMaskSewSelect_7_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_7 <= 1'h0;
      maskLastPipe_pipe_v_7 <= 1'h0;
      pipe_v_23 <= 1'h0;
      sinkVec_releasePipe_pipe_v_32 <= 1'h0;
      sinkVec_tokenCheck_counter_32 <= 3'h0;
      sinkVec_shifterReg_32_0_valid <= 1'h0;
      sinkVec_shifterReg_32_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_32_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_32_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_32_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_33 <= 1'h0;
      sinkVec_tokenCheck_counter_33 <= 3'h0;
      sinkVec_shifterReg_33_0_valid <= 1'h0;
      sinkVec_shifterReg_33_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_33_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_33_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_33_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_16 <= 1'h0;
      accessDataValid_pipe_v_16 <= 1'h0;
      accessDataValid_pipe_pipe_v_16 <= 1'h0;
      shifterReg_32_0_valid <= 1'h0;
      shifterReg_32_0_bits <= 32'h0;
      accessDataValid_pipe_v_17 <= 1'h0;
      accessDataValid_pipe_pipe_v_17 <= 1'h0;
      shifterReg_33_0_valid <= 1'h0;
      shifterReg_33_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_34 <= 1'h0;
      sinkVec_tokenCheck_counter_34 <= 3'h0;
      sinkVec_shifterReg_34_0_valid <= 1'h0;
      sinkVec_shifterReg_34_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_34_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_34_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_34_0_bits_data <= 32'h0;
      sinkVec_shifterReg_34_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_35 <= 1'h0;
      sinkVec_tokenCheck_counter_35 <= 3'h0;
      sinkVec_shifterReg_35_0_valid <= 1'h0;
      sinkVec_shifterReg_35_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_35_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_35_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_35_0_bits_data <= 32'h0;
      sinkVec_shifterReg_35_0_bits_last <= 1'h0;
      sinkVec_shifterReg_35_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_17 <= 1'h0;
      view__writeRelease_8_pipe_v <= 1'h0;
      pipe_v_24 <= 1'h0;
      instructionFinishedPipe_pipe_v_8 <= 1'h0;
      pipe_v_25 <= 1'h0;
      pipe_pipe_v_8 <= 1'h0;
      view__laneMaskSelect_8_pipe_v <= 1'h0;
      view__laneMaskSelect_8_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_8_pipe_v <= 1'h0;
      view__laneMaskSewSelect_8_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_8 <= 1'h0;
      maskLastPipe_pipe_v_8 <= 1'h0;
      pipe_v_26 <= 1'h0;
      sinkVec_releasePipe_pipe_v_36 <= 1'h0;
      sinkVec_tokenCheck_counter_36 <= 3'h0;
      sinkVec_shifterReg_36_0_valid <= 1'h0;
      sinkVec_shifterReg_36_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_36_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_36_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_36_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_37 <= 1'h0;
      sinkVec_tokenCheck_counter_37 <= 3'h0;
      sinkVec_shifterReg_37_0_valid <= 1'h0;
      sinkVec_shifterReg_37_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_37_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_37_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_37_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_18 <= 1'h0;
      accessDataValid_pipe_v_18 <= 1'h0;
      accessDataValid_pipe_pipe_v_18 <= 1'h0;
      shifterReg_34_0_valid <= 1'h0;
      shifterReg_34_0_bits <= 32'h0;
      accessDataValid_pipe_v_19 <= 1'h0;
      accessDataValid_pipe_pipe_v_19 <= 1'h0;
      shifterReg_35_0_valid <= 1'h0;
      shifterReg_35_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_38 <= 1'h0;
      sinkVec_tokenCheck_counter_38 <= 3'h0;
      sinkVec_shifterReg_38_0_valid <= 1'h0;
      sinkVec_shifterReg_38_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_38_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_38_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_38_0_bits_data <= 32'h0;
      sinkVec_shifterReg_38_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_39 <= 1'h0;
      sinkVec_tokenCheck_counter_39 <= 3'h0;
      sinkVec_shifterReg_39_0_valid <= 1'h0;
      sinkVec_shifterReg_39_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_39_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_39_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_39_0_bits_data <= 32'h0;
      sinkVec_shifterReg_39_0_bits_last <= 1'h0;
      sinkVec_shifterReg_39_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_19 <= 1'h0;
      view__writeRelease_9_pipe_v <= 1'h0;
      pipe_v_27 <= 1'h0;
      instructionFinishedPipe_pipe_v_9 <= 1'h0;
      pipe_v_28 <= 1'h0;
      pipe_pipe_v_9 <= 1'h0;
      view__laneMaskSelect_9_pipe_v <= 1'h0;
      view__laneMaskSelect_9_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_9_pipe_v <= 1'h0;
      view__laneMaskSewSelect_9_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_9 <= 1'h0;
      maskLastPipe_pipe_v_9 <= 1'h0;
      pipe_v_29 <= 1'h0;
      sinkVec_releasePipe_pipe_v_40 <= 1'h0;
      sinkVec_tokenCheck_counter_40 <= 3'h0;
      sinkVec_shifterReg_40_0_valid <= 1'h0;
      sinkVec_shifterReg_40_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_40_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_40_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_40_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_41 <= 1'h0;
      sinkVec_tokenCheck_counter_41 <= 3'h0;
      sinkVec_shifterReg_41_0_valid <= 1'h0;
      sinkVec_shifterReg_41_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_41_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_41_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_41_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_20 <= 1'h0;
      accessDataValid_pipe_v_20 <= 1'h0;
      accessDataValid_pipe_pipe_v_20 <= 1'h0;
      shifterReg_36_0_valid <= 1'h0;
      shifterReg_36_0_bits <= 32'h0;
      accessDataValid_pipe_v_21 <= 1'h0;
      accessDataValid_pipe_pipe_v_21 <= 1'h0;
      shifterReg_37_0_valid <= 1'h0;
      shifterReg_37_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_42 <= 1'h0;
      sinkVec_tokenCheck_counter_42 <= 3'h0;
      sinkVec_shifterReg_42_0_valid <= 1'h0;
      sinkVec_shifterReg_42_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_42_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_42_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_42_0_bits_data <= 32'h0;
      sinkVec_shifterReg_42_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_43 <= 1'h0;
      sinkVec_tokenCheck_counter_43 <= 3'h0;
      sinkVec_shifterReg_43_0_valid <= 1'h0;
      sinkVec_shifterReg_43_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_43_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_43_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_43_0_bits_data <= 32'h0;
      sinkVec_shifterReg_43_0_bits_last <= 1'h0;
      sinkVec_shifterReg_43_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_21 <= 1'h0;
      view__writeRelease_10_pipe_v <= 1'h0;
      pipe_v_30 <= 1'h0;
      instructionFinishedPipe_pipe_v_10 <= 1'h0;
      pipe_v_31 <= 1'h0;
      pipe_pipe_v_10 <= 1'h0;
      view__laneMaskSelect_10_pipe_v <= 1'h0;
      view__laneMaskSelect_10_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_10_pipe_v <= 1'h0;
      view__laneMaskSewSelect_10_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_10 <= 1'h0;
      maskLastPipe_pipe_v_10 <= 1'h0;
      pipe_v_32 <= 1'h0;
      sinkVec_releasePipe_pipe_v_44 <= 1'h0;
      sinkVec_tokenCheck_counter_44 <= 3'h0;
      sinkVec_shifterReg_44_0_valid <= 1'h0;
      sinkVec_shifterReg_44_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_44_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_44_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_44_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_45 <= 1'h0;
      sinkVec_tokenCheck_counter_45 <= 3'h0;
      sinkVec_shifterReg_45_0_valid <= 1'h0;
      sinkVec_shifterReg_45_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_45_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_45_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_45_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_22 <= 1'h0;
      accessDataValid_pipe_v_22 <= 1'h0;
      accessDataValid_pipe_pipe_v_22 <= 1'h0;
      shifterReg_38_0_valid <= 1'h0;
      shifterReg_38_0_bits <= 32'h0;
      accessDataValid_pipe_v_23 <= 1'h0;
      accessDataValid_pipe_pipe_v_23 <= 1'h0;
      shifterReg_39_0_valid <= 1'h0;
      shifterReg_39_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_46 <= 1'h0;
      sinkVec_tokenCheck_counter_46 <= 3'h0;
      sinkVec_shifterReg_46_0_valid <= 1'h0;
      sinkVec_shifterReg_46_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_46_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_46_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_46_0_bits_data <= 32'h0;
      sinkVec_shifterReg_46_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_47 <= 1'h0;
      sinkVec_tokenCheck_counter_47 <= 3'h0;
      sinkVec_shifterReg_47_0_valid <= 1'h0;
      sinkVec_shifterReg_47_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_47_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_47_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_47_0_bits_data <= 32'h0;
      sinkVec_shifterReg_47_0_bits_last <= 1'h0;
      sinkVec_shifterReg_47_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_23 <= 1'h0;
      view__writeRelease_11_pipe_v <= 1'h0;
      pipe_v_33 <= 1'h0;
      instructionFinishedPipe_pipe_v_11 <= 1'h0;
      pipe_v_34 <= 1'h0;
      pipe_pipe_v_11 <= 1'h0;
      view__laneMaskSelect_11_pipe_v <= 1'h0;
      view__laneMaskSelect_11_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_11_pipe_v <= 1'h0;
      view__laneMaskSewSelect_11_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_11 <= 1'h0;
      maskLastPipe_pipe_v_11 <= 1'h0;
      pipe_v_35 <= 1'h0;
      sinkVec_releasePipe_pipe_v_48 <= 1'h0;
      sinkVec_tokenCheck_counter_48 <= 3'h0;
      sinkVec_shifterReg_48_0_valid <= 1'h0;
      sinkVec_shifterReg_48_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_48_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_48_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_48_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_49 <= 1'h0;
      sinkVec_tokenCheck_counter_49 <= 3'h0;
      sinkVec_shifterReg_49_0_valid <= 1'h0;
      sinkVec_shifterReg_49_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_49_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_49_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_49_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_24 <= 1'h0;
      accessDataValid_pipe_v_24 <= 1'h0;
      accessDataValid_pipe_pipe_v_24 <= 1'h0;
      shifterReg_40_0_valid <= 1'h0;
      shifterReg_40_0_bits <= 32'h0;
      accessDataValid_pipe_v_25 <= 1'h0;
      accessDataValid_pipe_pipe_v_25 <= 1'h0;
      shifterReg_41_0_valid <= 1'h0;
      shifterReg_41_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_50 <= 1'h0;
      sinkVec_tokenCheck_counter_50 <= 3'h0;
      sinkVec_shifterReg_50_0_valid <= 1'h0;
      sinkVec_shifterReg_50_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_50_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_50_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_50_0_bits_data <= 32'h0;
      sinkVec_shifterReg_50_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_51 <= 1'h0;
      sinkVec_tokenCheck_counter_51 <= 3'h0;
      sinkVec_shifterReg_51_0_valid <= 1'h0;
      sinkVec_shifterReg_51_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_51_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_51_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_51_0_bits_data <= 32'h0;
      sinkVec_shifterReg_51_0_bits_last <= 1'h0;
      sinkVec_shifterReg_51_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_25 <= 1'h0;
      view__writeRelease_12_pipe_v <= 1'h0;
      pipe_v_36 <= 1'h0;
      instructionFinishedPipe_pipe_v_12 <= 1'h0;
      pipe_v_37 <= 1'h0;
      pipe_pipe_v_12 <= 1'h0;
      view__laneMaskSelect_12_pipe_v <= 1'h0;
      view__laneMaskSelect_12_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_12_pipe_v <= 1'h0;
      view__laneMaskSewSelect_12_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_12 <= 1'h0;
      maskLastPipe_pipe_v_12 <= 1'h0;
      pipe_v_38 <= 1'h0;
      sinkVec_releasePipe_pipe_v_52 <= 1'h0;
      sinkVec_tokenCheck_counter_52 <= 3'h0;
      sinkVec_shifterReg_52_0_valid <= 1'h0;
      sinkVec_shifterReg_52_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_52_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_52_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_52_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_53 <= 1'h0;
      sinkVec_tokenCheck_counter_53 <= 3'h0;
      sinkVec_shifterReg_53_0_valid <= 1'h0;
      sinkVec_shifterReg_53_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_53_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_53_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_53_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_26 <= 1'h0;
      accessDataValid_pipe_v_26 <= 1'h0;
      accessDataValid_pipe_pipe_v_26 <= 1'h0;
      shifterReg_42_0_valid <= 1'h0;
      shifterReg_42_0_bits <= 32'h0;
      accessDataValid_pipe_v_27 <= 1'h0;
      accessDataValid_pipe_pipe_v_27 <= 1'h0;
      shifterReg_43_0_valid <= 1'h0;
      shifterReg_43_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_54 <= 1'h0;
      sinkVec_tokenCheck_counter_54 <= 3'h0;
      sinkVec_shifterReg_54_0_valid <= 1'h0;
      sinkVec_shifterReg_54_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_54_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_54_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_54_0_bits_data <= 32'h0;
      sinkVec_shifterReg_54_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_55 <= 1'h0;
      sinkVec_tokenCheck_counter_55 <= 3'h0;
      sinkVec_shifterReg_55_0_valid <= 1'h0;
      sinkVec_shifterReg_55_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_55_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_55_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_55_0_bits_data <= 32'h0;
      sinkVec_shifterReg_55_0_bits_last <= 1'h0;
      sinkVec_shifterReg_55_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_27 <= 1'h0;
      view__writeRelease_13_pipe_v <= 1'h0;
      pipe_v_39 <= 1'h0;
      instructionFinishedPipe_pipe_v_13 <= 1'h0;
      pipe_v_40 <= 1'h0;
      pipe_pipe_v_13 <= 1'h0;
      view__laneMaskSelect_13_pipe_v <= 1'h0;
      view__laneMaskSelect_13_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_13_pipe_v <= 1'h0;
      view__laneMaskSewSelect_13_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_13 <= 1'h0;
      maskLastPipe_pipe_v_13 <= 1'h0;
      pipe_v_41 <= 1'h0;
      sinkVec_releasePipe_pipe_v_56 <= 1'h0;
      sinkVec_tokenCheck_counter_56 <= 3'h0;
      sinkVec_shifterReg_56_0_valid <= 1'h0;
      sinkVec_shifterReg_56_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_56_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_56_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_56_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_57 <= 1'h0;
      sinkVec_tokenCheck_counter_57 <= 3'h0;
      sinkVec_shifterReg_57_0_valid <= 1'h0;
      sinkVec_shifterReg_57_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_57_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_57_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_57_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_28 <= 1'h0;
      accessDataValid_pipe_v_28 <= 1'h0;
      accessDataValid_pipe_pipe_v_28 <= 1'h0;
      shifterReg_44_0_valid <= 1'h0;
      shifterReg_44_0_bits <= 32'h0;
      accessDataValid_pipe_v_29 <= 1'h0;
      accessDataValid_pipe_pipe_v_29 <= 1'h0;
      shifterReg_45_0_valid <= 1'h0;
      shifterReg_45_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_58 <= 1'h0;
      sinkVec_tokenCheck_counter_58 <= 3'h0;
      sinkVec_shifterReg_58_0_valid <= 1'h0;
      sinkVec_shifterReg_58_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_58_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_58_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_58_0_bits_data <= 32'h0;
      sinkVec_shifterReg_58_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_59 <= 1'h0;
      sinkVec_tokenCheck_counter_59 <= 3'h0;
      sinkVec_shifterReg_59_0_valid <= 1'h0;
      sinkVec_shifterReg_59_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_59_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_59_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_59_0_bits_data <= 32'h0;
      sinkVec_shifterReg_59_0_bits_last <= 1'h0;
      sinkVec_shifterReg_59_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_29 <= 1'h0;
      view__writeRelease_14_pipe_v <= 1'h0;
      pipe_v_42 <= 1'h0;
      instructionFinishedPipe_pipe_v_14 <= 1'h0;
      pipe_v_43 <= 1'h0;
      pipe_pipe_v_14 <= 1'h0;
      view__laneMaskSelect_14_pipe_v <= 1'h0;
      view__laneMaskSelect_14_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_14_pipe_v <= 1'h0;
      view__laneMaskSewSelect_14_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_14 <= 1'h0;
      maskLastPipe_pipe_v_14 <= 1'h0;
      pipe_v_44 <= 1'h0;
      sinkVec_releasePipe_pipe_v_60 <= 1'h0;
      sinkVec_tokenCheck_counter_60 <= 3'h0;
      sinkVec_shifterReg_60_0_valid <= 1'h0;
      sinkVec_shifterReg_60_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_60_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_60_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_60_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_61 <= 1'h0;
      sinkVec_tokenCheck_counter_61 <= 3'h0;
      sinkVec_shifterReg_61_0_valid <= 1'h0;
      sinkVec_shifterReg_61_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_61_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_61_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_61_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_30 <= 1'h0;
      accessDataValid_pipe_v_30 <= 1'h0;
      accessDataValid_pipe_pipe_v_30 <= 1'h0;
      shifterReg_46_0_valid <= 1'h0;
      shifterReg_46_0_bits <= 32'h0;
      accessDataValid_pipe_v_31 <= 1'h0;
      accessDataValid_pipe_pipe_v_31 <= 1'h0;
      shifterReg_47_0_valid <= 1'h0;
      shifterReg_47_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_62 <= 1'h0;
      sinkVec_tokenCheck_counter_62 <= 3'h0;
      sinkVec_shifterReg_62_0_valid <= 1'h0;
      sinkVec_shifterReg_62_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_62_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_62_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_62_0_bits_data <= 32'h0;
      sinkVec_shifterReg_62_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_63 <= 1'h0;
      sinkVec_tokenCheck_counter_63 <= 3'h0;
      sinkVec_shifterReg_63_0_valid <= 1'h0;
      sinkVec_shifterReg_63_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_63_0_bits_offset <= 2'h0;
      sinkVec_shifterReg_63_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_63_0_bits_data <= 32'h0;
      sinkVec_shifterReg_63_0_bits_last <= 1'h0;
      sinkVec_shifterReg_63_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_31 <= 1'h0;
      view__writeRelease_15_pipe_v <= 1'h0;
      pipe_v_45 <= 1'h0;
      instructionFinishedPipe_pipe_v_15 <= 1'h0;
      pipe_v_46 <= 1'h0;
      pipe_pipe_v_15 <= 1'h0;
      view__laneMaskSelect_15_pipe_v <= 1'h0;
      view__laneMaskSelect_15_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_15_pipe_v <= 1'h0;
      view__laneMaskSewSelect_15_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_15 <= 1'h0;
      maskLastPipe_pipe_v_15 <= 1'h0;
      pipe_v_47 <= 1'h0;
      pipe_v_48 <= 1'h0;
      shifterReg_48_0_valid <= 1'h0;
      shifterReg_48_0_bits_data <= 32'h0;
      pipe_v_49 <= 1'h0;
      shifterReg_49_0_valid <= 1'h0;
      shifterReg_49_0_bits_data <= 32'h0;
      shifterReg_49_0_bits_mask <= 2'h0;
      shifterReg_49_0_bits_instructionIndex <= 3'h0;
      shifterReg_49_0_bits_counter <= 6'h0;
      pipe_v_50 <= 1'h0;
      shifterReg_50_0_valid <= 1'h0;
      shifterReg_50_0_bits_data <= 32'h0;
      pipe_v_51 <= 1'h0;
      shifterReg_51_0_valid <= 1'h0;
      shifterReg_51_0_bits_data <= 32'h0;
      shifterReg_51_0_bits_mask <= 2'h0;
      shifterReg_51_0_bits_instructionIndex <= 3'h0;
      shifterReg_51_0_bits_counter <= 6'h0;
      pipe_v_52 <= 1'h0;
      shifterReg_52_0_valid <= 1'h0;
      shifterReg_52_0_bits_data <= 32'h0;
      pipe_v_53 <= 1'h0;
      shifterReg_53_0_valid <= 1'h0;
      shifterReg_53_0_bits_data <= 32'h0;
      shifterReg_53_0_bits_mask <= 2'h0;
      shifterReg_53_0_bits_instructionIndex <= 3'h0;
      shifterReg_53_0_bits_counter <= 6'h0;
      pipe_v_54 <= 1'h0;
      shifterReg_54_0_valid <= 1'h0;
      shifterReg_54_0_bits_data <= 32'h0;
      pipe_v_55 <= 1'h0;
      shifterReg_55_0_valid <= 1'h0;
      shifterReg_55_0_bits_data <= 32'h0;
      shifterReg_55_0_bits_mask <= 2'h0;
      shifterReg_55_0_bits_instructionIndex <= 3'h0;
      shifterReg_55_0_bits_counter <= 6'h0;
      pipe_v_56 <= 1'h0;
      shifterReg_56_0_valid <= 1'h0;
      shifterReg_56_0_bits_data <= 32'h0;
      pipe_v_57 <= 1'h0;
      shifterReg_57_0_valid <= 1'h0;
      shifterReg_57_0_bits_data <= 32'h0;
      shifterReg_57_0_bits_mask <= 2'h0;
      shifterReg_57_0_bits_instructionIndex <= 3'h0;
      shifterReg_57_0_bits_counter <= 6'h0;
      pipe_v_58 <= 1'h0;
      shifterReg_58_0_valid <= 1'h0;
      shifterReg_58_0_bits_data <= 32'h0;
      pipe_v_59 <= 1'h0;
      shifterReg_59_0_valid <= 1'h0;
      shifterReg_59_0_bits_data <= 32'h0;
      shifterReg_59_0_bits_mask <= 2'h0;
      shifterReg_59_0_bits_instructionIndex <= 3'h0;
      shifterReg_59_0_bits_counter <= 6'h0;
      pipe_v_60 <= 1'h0;
      shifterReg_60_0_valid <= 1'h0;
      shifterReg_60_0_bits_data <= 32'h0;
      pipe_v_61 <= 1'h0;
      shifterReg_61_0_valid <= 1'h0;
      shifterReg_61_0_bits_data <= 32'h0;
      shifterReg_61_0_bits_mask <= 2'h0;
      shifterReg_61_0_bits_instructionIndex <= 3'h0;
      shifterReg_61_0_bits_counter <= 6'h0;
      pipe_v_62 <= 1'h0;
      shifterReg_62_0_valid <= 1'h0;
      shifterReg_62_0_bits_data <= 32'h0;
      pipe_v_63 <= 1'h0;
      shifterReg_63_0_valid <= 1'h0;
      shifterReg_63_0_bits_data <= 32'h0;
      shifterReg_63_0_bits_mask <= 2'h0;
      shifterReg_63_0_bits_instructionIndex <= 3'h0;
      shifterReg_63_0_bits_counter <= 6'h0;
      pipe_v_64 <= 1'h0;
      shifterReg_64_0_valid <= 1'h0;
      shifterReg_64_0_bits_data <= 32'h0;
      pipe_v_65 <= 1'h0;
      shifterReg_65_0_valid <= 1'h0;
      shifterReg_65_0_bits_data <= 32'h0;
      shifterReg_65_0_bits_mask <= 2'h0;
      shifterReg_65_0_bits_instructionIndex <= 3'h0;
      shifterReg_65_0_bits_counter <= 6'h0;
      pipe_v_66 <= 1'h0;
      shifterReg_66_0_valid <= 1'h0;
      shifterReg_66_0_bits_data <= 32'h0;
      pipe_v_67 <= 1'h0;
      shifterReg_67_0_valid <= 1'h0;
      shifterReg_67_0_bits_data <= 32'h0;
      shifterReg_67_0_bits_mask <= 2'h0;
      shifterReg_67_0_bits_instructionIndex <= 3'h0;
      shifterReg_67_0_bits_counter <= 6'h0;
      pipe_v_68 <= 1'h0;
      shifterReg_68_0_valid <= 1'h0;
      shifterReg_68_0_bits_data <= 32'h0;
      pipe_v_69 <= 1'h0;
      shifterReg_69_0_valid <= 1'h0;
      shifterReg_69_0_bits_data <= 32'h0;
      shifterReg_69_0_bits_mask <= 2'h0;
      shifterReg_69_0_bits_instructionIndex <= 3'h0;
      shifterReg_69_0_bits_counter <= 6'h0;
      pipe_v_70 <= 1'h0;
      shifterReg_70_0_valid <= 1'h0;
      shifterReg_70_0_bits_data <= 32'h0;
      pipe_v_71 <= 1'h0;
      shifterReg_71_0_valid <= 1'h0;
      shifterReg_71_0_bits_data <= 32'h0;
      shifterReg_71_0_bits_mask <= 2'h0;
      shifterReg_71_0_bits_instructionIndex <= 3'h0;
      shifterReg_71_0_bits_counter <= 6'h0;
      pipe_v_72 <= 1'h0;
      shifterReg_72_0_valid <= 1'h0;
      shifterReg_72_0_bits_data <= 32'h0;
      pipe_v_73 <= 1'h0;
      shifterReg_73_0_valid <= 1'h0;
      shifterReg_73_0_bits_data <= 32'h0;
      shifterReg_73_0_bits_mask <= 2'h0;
      shifterReg_73_0_bits_instructionIndex <= 3'h0;
      shifterReg_73_0_bits_counter <= 6'h0;
      pipe_v_74 <= 1'h0;
      shifterReg_74_0_valid <= 1'h0;
      shifterReg_74_0_bits_data <= 32'h0;
      pipe_v_75 <= 1'h0;
      shifterReg_75_0_valid <= 1'h0;
      shifterReg_75_0_bits_data <= 32'h0;
      shifterReg_75_0_bits_mask <= 2'h0;
      shifterReg_75_0_bits_instructionIndex <= 3'h0;
      shifterReg_75_0_bits_counter <= 6'h0;
      pipe_v_76 <= 1'h0;
      shifterReg_76_0_valid <= 1'h0;
      shifterReg_76_0_bits_data <= 32'h0;
      pipe_v_77 <= 1'h0;
      shifterReg_77_0_valid <= 1'h0;
      shifterReg_77_0_bits_data <= 32'h0;
      shifterReg_77_0_bits_mask <= 2'h0;
      shifterReg_77_0_bits_instructionIndex <= 3'h0;
      shifterReg_77_0_bits_counter <= 6'h0;
      pipe_v_78 <= 1'h0;
      shifterReg_78_0_valid <= 1'h0;
      shifterReg_78_0_bits_data <= 32'h0;
      pipe_v_79 <= 1'h0;
      shifterReg_79_0_valid <= 1'h0;
      shifterReg_79_0_bits_data <= 32'h0;
      shifterReg_79_0_bits_mask <= 2'h0;
      shifterReg_79_0_bits_instructionIndex <= 3'h0;
      shifterReg_79_0_bits_counter <= 6'h0;
      pipe_v_80 <= 1'h0;
      shifterReg_80_0_valid <= 1'h0;
      shifterReg_80_0_bits_data <= 32'h0;
      pipe_v_81 <= 1'h0;
      shifterReg_81_0_valid <= 1'h0;
      shifterReg_81_0_bits_data <= 32'h0;
      shifterReg_81_0_bits_mask <= 2'h0;
      shifterReg_81_0_bits_instructionIndex <= 3'h0;
      shifterReg_81_0_bits_counter <= 6'h0;
      pipe_v_82 <= 1'h0;
      shifterReg_82_0_valid <= 1'h0;
      shifterReg_82_0_bits_data <= 32'h0;
      pipe_v_83 <= 1'h0;
      shifterReg_83_0_valid <= 1'h0;
      shifterReg_83_0_bits_data <= 32'h0;
      shifterReg_83_0_bits_mask <= 2'h0;
      shifterReg_83_0_bits_instructionIndex <= 3'h0;
      shifterReg_83_0_bits_counter <= 6'h0;
      pipe_v_84 <= 1'h0;
      shifterReg_84_0_valid <= 1'h0;
      shifterReg_84_0_bits_data <= 32'h0;
      pipe_v_85 <= 1'h0;
      shifterReg_85_0_valid <= 1'h0;
      shifterReg_85_0_bits_data <= 32'h0;
      shifterReg_85_0_bits_mask <= 2'h0;
      shifterReg_85_0_bits_instructionIndex <= 3'h0;
      shifterReg_85_0_bits_counter <= 6'h0;
      pipe_v_86 <= 1'h0;
      shifterReg_86_0_valid <= 1'h0;
      shifterReg_86_0_bits_data <= 32'h0;
      pipe_v_87 <= 1'h0;
      shifterReg_87_0_valid <= 1'h0;
      shifterReg_87_0_bits_data <= 32'h0;
      shifterReg_87_0_bits_mask <= 2'h0;
      shifterReg_87_0_bits_instructionIndex <= 3'h0;
      shifterReg_87_0_bits_counter <= 6'h0;
      pipe_v_88 <= 1'h0;
      shifterReg_88_0_valid <= 1'h0;
      shifterReg_88_0_bits_data <= 32'h0;
      pipe_v_89 <= 1'h0;
      shifterReg_89_0_valid <= 1'h0;
      shifterReg_89_0_bits_data <= 32'h0;
      shifterReg_89_0_bits_mask <= 2'h0;
      shifterReg_89_0_bits_instructionIndex <= 3'h0;
      shifterReg_89_0_bits_counter <= 6'h0;
      pipe_v_90 <= 1'h0;
      shifterReg_90_0_valid <= 1'h0;
      shifterReg_90_0_bits_data <= 32'h0;
      pipe_v_91 <= 1'h0;
      shifterReg_91_0_valid <= 1'h0;
      shifterReg_91_0_bits_data <= 32'h0;
      shifterReg_91_0_bits_mask <= 2'h0;
      shifterReg_91_0_bits_instructionIndex <= 3'h0;
      shifterReg_91_0_bits_counter <= 6'h0;
      pipe_v_92 <= 1'h0;
      shifterReg_92_0_valid <= 1'h0;
      shifterReg_92_0_bits_data <= 32'h0;
      pipe_v_93 <= 1'h0;
      shifterReg_93_0_valid <= 1'h0;
      shifterReg_93_0_bits_data <= 32'h0;
      shifterReg_93_0_bits_mask <= 2'h0;
      shifterReg_93_0_bits_instructionIndex <= 3'h0;
      shifterReg_93_0_bits_counter <= 6'h0;
      pipe_v_94 <= 1'h0;
      shifterReg_94_0_valid <= 1'h0;
      shifterReg_94_0_bits_data <= 32'h0;
      pipe_v_95 <= 1'h0;
      shifterReg_95_0_valid <= 1'h0;
      shifterReg_95_0_bits_data <= 32'h0;
      shifterReg_95_0_bits_mask <= 2'h0;
      shifterReg_95_0_bits_instructionIndex <= 3'h0;
      shifterReg_95_0_bits_counter <= 6'h0;
      pipe_v_96 <= 1'h0;
      shifterReg_96_0_valid <= 1'h0;
      shifterReg_96_0_bits_data <= 32'h0;
      pipe_v_97 <= 1'h0;
      shifterReg_97_0_valid <= 1'h0;
      shifterReg_97_0_bits_data <= 32'h0;
      shifterReg_97_0_bits_mask <= 2'h0;
      shifterReg_97_0_bits_instructionIndex <= 3'h0;
      shifterReg_97_0_bits_counter <= 6'h0;
      pipe_v_98 <= 1'h0;
      shifterReg_98_0_valid <= 1'h0;
      shifterReg_98_0_bits_data <= 32'h0;
      pipe_v_99 <= 1'h0;
      shifterReg_99_0_valid <= 1'h0;
      shifterReg_99_0_bits_data <= 32'h0;
      shifterReg_99_0_bits_mask <= 2'h0;
      shifterReg_99_0_bits_instructionIndex <= 3'h0;
      shifterReg_99_0_bits_counter <= 6'h0;
      pipe_v_100 <= 1'h0;
      shifterReg_100_0_valid <= 1'h0;
      shifterReg_100_0_bits_data <= 32'h0;
      pipe_v_101 <= 1'h0;
      shifterReg_101_0_valid <= 1'h0;
      shifterReg_101_0_bits_data <= 32'h0;
      shifterReg_101_0_bits_mask <= 2'h0;
      shifterReg_101_0_bits_instructionIndex <= 3'h0;
      shifterReg_101_0_bits_counter <= 6'h0;
      pipe_v_102 <= 1'h0;
      shifterReg_102_0_valid <= 1'h0;
      shifterReg_102_0_bits_data <= 32'h0;
      pipe_v_103 <= 1'h0;
      shifterReg_103_0_valid <= 1'h0;
      shifterReg_103_0_bits_data <= 32'h0;
      shifterReg_103_0_bits_mask <= 2'h0;
      shifterReg_103_0_bits_instructionIndex <= 3'h0;
      shifterReg_103_0_bits_counter <= 6'h0;
      pipe_v_104 <= 1'h0;
      shifterReg_104_0_valid <= 1'h0;
      shifterReg_104_0_bits_data <= 32'h0;
      pipe_v_105 <= 1'h0;
      shifterReg_105_0_valid <= 1'h0;
      shifterReg_105_0_bits_data <= 32'h0;
      shifterReg_105_0_bits_mask <= 2'h0;
      shifterReg_105_0_bits_instructionIndex <= 3'h0;
      shifterReg_105_0_bits_counter <= 6'h0;
      pipe_v_106 <= 1'h0;
      shifterReg_106_0_valid <= 1'h0;
      shifterReg_106_0_bits_data <= 32'h0;
      pipe_v_107 <= 1'h0;
      shifterReg_107_0_valid <= 1'h0;
      shifterReg_107_0_bits_data <= 32'h0;
      shifterReg_107_0_bits_mask <= 2'h0;
      shifterReg_107_0_bits_instructionIndex <= 3'h0;
      shifterReg_107_0_bits_counter <= 6'h0;
      pipe_v_108 <= 1'h0;
      shifterReg_108_0_valid <= 1'h0;
      shifterReg_108_0_bits_data <= 32'h0;
      pipe_v_109 <= 1'h0;
      shifterReg_109_0_valid <= 1'h0;
      shifterReg_109_0_bits_data <= 32'h0;
      shifterReg_109_0_bits_mask <= 2'h0;
      shifterReg_109_0_bits_instructionIndex <= 3'h0;
      shifterReg_109_0_bits_counter <= 6'h0;
      pipe_v_110 <= 1'h0;
      shifterReg_110_0_valid <= 1'h0;
      shifterReg_110_0_bits_data <= 32'h0;
      pipe_v_111 <= 1'h0;
      shifterReg_111_0_valid <= 1'h0;
      shifterReg_111_0_bits_data <= 32'h0;
      shifterReg_111_0_bits_mask <= 2'h0;
      shifterReg_111_0_bits_instructionIndex <= 3'h0;
      shifterReg_111_0_bits_counter <= 6'h0;
    end
    else begin
      if (_probeWire_issue_valid_T) begin
        automatic logic [38:0] _requestReg_bits_writeByte_T_8 = {7'h0, issue_bits_vl_0} << issue_bits_vtype_0[5:3] + {2'h0, _decode_decodeResult_crossWrite};
        instructionCounter <= nextInstructionCounter;
        requestReg_bits_issue_instruction <= issue_bits_instruction_0;
        requestReg_bits_issue_rs1Data <= issue_bits_rs1Data_0;
        requestReg_bits_issue_rs2Data <= issue_bits_rs2Data_0;
        requestReg_bits_issue_vtype <= issue_bits_vtype_0;
        requestReg_bits_issue_vl <= issue_bits_vl_0;
        requestReg_bits_issue_vstart <= issue_bits_vstart_0;
        requestReg_bits_issue_vcsr <= issue_bits_vcsr_0;
        requestReg_bits_decodeResult_orderReduce <= _decode_decodeResult_orderReduce;
        requestReg_bits_decodeResult_floatMul <= _decode_decodeResult_floatMul;
        requestReg_bits_decodeResult_fpExecutionType <= _decode_decodeResult_fpExecutionType;
        requestReg_bits_decodeResult_float <= _decode_decodeResult_float;
        requestReg_bits_decodeResult_specialSlot <= _decode_decodeResult_specialSlot;
        requestReg_bits_decodeResult_topUop <= _decode_decodeResult_topUop;
        requestReg_bits_decodeResult_popCount <= _decode_decodeResult_popCount;
        requestReg_bits_decodeResult_ffo <= _decode_decodeResult_ffo;
        requestReg_bits_decodeResult_average <= _decode_decodeResult_average;
        requestReg_bits_decodeResult_reverse <= _decode_decodeResult_reverse;
        requestReg_bits_decodeResult_dontNeedExecuteInLane <= _decode_decodeResult_dontNeedExecuteInLane;
        requestReg_bits_decodeResult_scheduler <= _decode_decodeResult_scheduler;
        requestReg_bits_decodeResult_sReadVD <= _decode_decodeResult_sReadVD;
        requestReg_bits_decodeResult_vtype <= _decode_decodeResult_vtype;
        requestReg_bits_decodeResult_sWrite <= _decode_decodeResult_sWrite;
        requestReg_bits_decodeResult_crossRead <= _decode_decodeResult_crossRead;
        requestReg_bits_decodeResult_crossWrite <= _decode_decodeResult_crossWrite;
        requestReg_bits_decodeResult_maskUnit <= _decode_decodeResult_maskUnit;
        requestReg_bits_decodeResult_special <= _decode_decodeResult_special;
        requestReg_bits_decodeResult_saturate <= _decode_decodeResult_saturate;
        requestReg_bits_decodeResult_vwmacc <= _decode_decodeResult_vwmacc;
        requestReg_bits_decodeResult_readOnly <= _decode_decodeResult_readOnly;
        requestReg_bits_decodeResult_maskSource <= _decode_decodeResult_maskSource;
        requestReg_bits_decodeResult_maskDestination <= _decode_decodeResult_maskDestination;
        requestReg_bits_decodeResult_maskLogic <= _decode_decodeResult_maskLogic;
        requestReg_bits_decodeResult_uop <= _decode_decodeResult_uop;
        requestReg_bits_decodeResult_iota <= _decode_decodeResult_iota;
        requestReg_bits_decodeResult_mv <= _decode_decodeResult_mv;
        requestReg_bits_decodeResult_extend <= _decode_decodeResult_extend;
        requestReg_bits_decodeResult_unOrderWrite <= _decode_decodeResult_unOrderWrite;
        requestReg_bits_decodeResult_compress <= _decode_decodeResult_compress;
        requestReg_bits_decodeResult_gather16 <= _decode_decodeResult_gather16;
        requestReg_bits_decodeResult_gather <= _decode_decodeResult_gather;
        requestReg_bits_decodeResult_slid <= _decode_decodeResult_slid;
        requestReg_bits_decodeResult_targetRd <= _decode_decodeResult_targetRd;
        requestReg_bits_decodeResult_widenReduce <= _decode_decodeResult_widenReduce;
        requestReg_bits_decodeResult_red <= _decode_decodeResult_red;
        requestReg_bits_decodeResult_nr <= _decode_decodeResult_nr;
        requestReg_bits_decodeResult_itype <= _decode_decodeResult_itype;
        requestReg_bits_decodeResult_unsigned1 <= _decode_decodeResult_unsigned1;
        requestReg_bits_decodeResult_unsigned0 <= _decode_decodeResult_unsigned0;
        requestReg_bits_decodeResult_other <= _decode_decodeResult_other;
        requestReg_bits_decodeResult_multiCycle <= _decode_decodeResult_multiCycle;
        requestReg_bits_decodeResult_divider <= _decode_decodeResult_divider;
        requestReg_bits_decodeResult_multiplier <= _decode_decodeResult_multiplier;
        requestReg_bits_decodeResult_shift <= _decode_decodeResult_shift;
        requestReg_bits_decodeResult_adder <= _decode_decodeResult_adder;
        requestReg_bits_decodeResult_logic <= _decode_decodeResult_logic;
        requestReg_bits_instructionIndex <= instructionCounter;
        requestReg_bits_vdIsV0 <= issue_bits_instruction_0[11:7] == 5'h0 & (issue_bits_instruction_0[6] | ~(issue_bits_instruction_0[5]));
        requestReg_bits_writeByte <= _decode_decodeResult_red ? 12'h1 : _decode_decodeResult_maskDestination ? issue_bits_vl_0[14:3] + {11'h0, |(issue_bits_vl_0[2:0])} : _requestReg_bits_writeByte_T_8[11:0];
      end
      if (retire_1)
        responseCounter <= nextResponseCounter;
      if (_probeWire_issue_valid_T ^ maskUnit_gatherData_ready)
        requestReg_valid <= _probeWire_issue_valid_T;
      if (instructionToSlotOH[0]) begin
        slots_0_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_0_record_isLoadStore <= isLoadStoreType;
        slots_0_record_maskType <= maskType;
      end
      slots_0_state_wLast <= ~(instructionToSlotOH[0]) & (slots_laneAndLSUFinish & slots_v0WriteFinish | slots_0_state_wLast);
      slots_0_state_idle <= ~(instructionToSlotOH[0]) & (slots_0_state_sCommit & slots_0_state_wVRFWrite & slots_0_state_wMaskUnitLast | slots_0_state_idle);
      slots_0_state_wMaskUnitLast <= instructionToSlotOH[0] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_0_state_wMaskUnitLast;
      slots_0_state_wVRFWrite <= instructionToSlotOH[0] ? ~requestReg_bits_decodeResult_maskUnit : slots_0_state_wLast & slots_0_state_wMaskUnitLast & ~slots_dataInWritePipeCheck | slots_0_state_wVRFWrite;
      slots_0_state_sCommit <= ~(instructionToSlotOH[0]) & (responseCounter == slots_0_record_instructionIndex & retire_1 | slots_0_state_sCommit);
      slots_0_endTag_0 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_0 | instructionFinished_0_0;
      slots_0_endTag_1 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_1 | instructionFinished_1_0;
      slots_0_endTag_2 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_2 | instructionFinished_2_0;
      slots_0_endTag_3 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_3 | instructionFinished_3_0;
      slots_0_endTag_4 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_4 | instructionFinished_4_0;
      slots_0_endTag_5 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_5 | instructionFinished_5_0;
      slots_0_endTag_6 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_6 | instructionFinished_6_0;
      slots_0_endTag_7 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_7 | instructionFinished_7_0;
      slots_0_endTag_8 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_8 | instructionFinished_8_0;
      slots_0_endTag_9 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_9 | instructionFinished_9_0;
      slots_0_endTag_10 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_10 | instructionFinished_10_0;
      slots_0_endTag_11 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_11 | instructionFinished_11_0;
      slots_0_endTag_12 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_12 | instructionFinished_12_0;
      slots_0_endTag_13 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_13 | instructionFinished_13_0;
      slots_0_endTag_14 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_14 | instructionFinished_14_0;
      slots_0_endTag_15 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_15 | instructionFinished_15_0;
      slots_0_endTag_16 <= instructionToSlotOH[0] ? ~isLoadStoreType : slots_0_endTag_16 | slots_lsuFinished;
      slots_0_vxsat <= ~(instructionToSlotOH[0]) & (slots_vxsatUpdate | slots_0_vxsat);
      if (instructionToSlotOH[1]) begin
        slots_1_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_1_record_isLoadStore <= isLoadStoreType;
        slots_1_record_maskType <= maskType;
      end
      slots_1_state_wLast <= ~(instructionToSlotOH[1]) & (slots_laneAndLSUFinish_1 & slots_v0WriteFinish_1 | slots_1_state_wLast);
      slots_1_state_idle <= ~(instructionToSlotOH[1]) & (slots_1_state_sCommit & slots_1_state_wVRFWrite & slots_1_state_wMaskUnitLast | slots_1_state_idle);
      slots_1_state_wMaskUnitLast <= instructionToSlotOH[1] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_1_state_wMaskUnitLast;
      slots_1_state_wVRFWrite <= instructionToSlotOH[1] ? ~requestReg_bits_decodeResult_maskUnit : slots_1_state_wLast & slots_1_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_1 | slots_1_state_wVRFWrite;
      slots_1_state_sCommit <= ~(instructionToSlotOH[1]) & (responseCounter == slots_1_record_instructionIndex & retire_1 | slots_1_state_sCommit);
      slots_1_endTag_0 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_0 | instructionFinished_0_1;
      slots_1_endTag_1 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_1 | instructionFinished_1_1;
      slots_1_endTag_2 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_2 | instructionFinished_2_1;
      slots_1_endTag_3 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_3 | instructionFinished_3_1;
      slots_1_endTag_4 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_4 | instructionFinished_4_1;
      slots_1_endTag_5 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_5 | instructionFinished_5_1;
      slots_1_endTag_6 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_6 | instructionFinished_6_1;
      slots_1_endTag_7 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_7 | instructionFinished_7_1;
      slots_1_endTag_8 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_8 | instructionFinished_8_1;
      slots_1_endTag_9 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_9 | instructionFinished_9_1;
      slots_1_endTag_10 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_10 | instructionFinished_10_1;
      slots_1_endTag_11 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_11 | instructionFinished_11_1;
      slots_1_endTag_12 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_12 | instructionFinished_12_1;
      slots_1_endTag_13 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_13 | instructionFinished_13_1;
      slots_1_endTag_14 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_14 | instructionFinished_14_1;
      slots_1_endTag_15 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_15 | instructionFinished_15_1;
      slots_1_endTag_16 <= instructionToSlotOH[1] ? ~isLoadStoreType : slots_1_endTag_16 | slots_lsuFinished_1;
      slots_1_vxsat <= ~(instructionToSlotOH[1]) & (slots_vxsatUpdate_1 | slots_1_vxsat);
      if (instructionToSlotOH[2]) begin
        slots_2_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_2_record_isLoadStore <= isLoadStoreType;
        slots_2_record_maskType <= maskType;
      end
      slots_2_state_wLast <= ~(instructionToSlotOH[2]) & (slots_laneAndLSUFinish_2 & slots_v0WriteFinish_2 | slots_2_state_wLast);
      slots_2_state_idle <= ~(instructionToSlotOH[2]) & (slots_2_state_sCommit & slots_2_state_wVRFWrite & slots_2_state_wMaskUnitLast | slots_2_state_idle);
      slots_2_state_wMaskUnitLast <= instructionToSlotOH[2] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_2_state_wMaskUnitLast;
      slots_2_state_wVRFWrite <= instructionToSlotOH[2] ? ~requestReg_bits_decodeResult_maskUnit : slots_2_state_wLast & slots_2_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_2 | slots_2_state_wVRFWrite;
      slots_2_state_sCommit <= ~(instructionToSlotOH[2]) & (responseCounter == slots_2_record_instructionIndex & retire_1 | slots_2_state_sCommit);
      slots_2_endTag_0 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_0 | instructionFinished_0_2;
      slots_2_endTag_1 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_1 | instructionFinished_1_2;
      slots_2_endTag_2 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_2 | instructionFinished_2_2;
      slots_2_endTag_3 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_3 | instructionFinished_3_2;
      slots_2_endTag_4 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_4 | instructionFinished_4_2;
      slots_2_endTag_5 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_5 | instructionFinished_5_2;
      slots_2_endTag_6 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_6 | instructionFinished_6_2;
      slots_2_endTag_7 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_7 | instructionFinished_7_2;
      slots_2_endTag_8 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_8 | instructionFinished_8_2;
      slots_2_endTag_9 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_9 | instructionFinished_9_2;
      slots_2_endTag_10 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_10 | instructionFinished_10_2;
      slots_2_endTag_11 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_11 | instructionFinished_11_2;
      slots_2_endTag_12 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_12 | instructionFinished_12_2;
      slots_2_endTag_13 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_13 | instructionFinished_13_2;
      slots_2_endTag_14 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_14 | instructionFinished_14_2;
      slots_2_endTag_15 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_15 | instructionFinished_15_2;
      slots_2_endTag_16 <= instructionToSlotOH[2] ? ~isLoadStoreType : slots_2_endTag_16 | slots_lsuFinished_2;
      slots_2_vxsat <= ~(instructionToSlotOH[2]) & (slots_vxsatUpdate_2 | slots_2_vxsat);
      if (instructionToSlotOH[3]) begin
        slots_3_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_3_record_isLoadStore <= isLoadStoreType;
        slots_3_record_maskType <= maskType;
        slots_writeRD <= requestReg_bits_decodeResult_targetRd;
        slots_float <= requestReg_bits_decodeResult_float;
        slots_vd <= requestRegDequeue_bits_instruction[11:7];
      end
      slots_3_state_wLast <= ~(instructionToSlotOH[3]) & (slots_laneAndLSUFinish_3 & slots_v0WriteFinish_3 | slots_3_state_wLast);
      slots_3_state_idle <= ~(instructionToSlotOH[3]) & (slots_3_state_sCommit & slots_3_state_wVRFWrite & slots_3_state_wMaskUnitLast | slots_3_state_idle);
      slots_3_state_wMaskUnitLast <= instructionToSlotOH[3] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_3_state_wMaskUnitLast;
      slots_3_state_wVRFWrite <= instructionToSlotOH[3] ? ~requestReg_bits_decodeResult_maskUnit : slots_3_state_wLast & slots_3_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_3 | slots_3_state_wVRFWrite;
      slots_3_state_sCommit <= ~(instructionToSlotOH[3]) & (responseCounter == slots_3_record_instructionIndex & retire_1 | slots_3_state_sCommit);
      slots_3_endTag_0 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_0 | instructionFinished_0_3;
      slots_3_endTag_1 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_1 | instructionFinished_1_3;
      slots_3_endTag_2 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_2 | instructionFinished_2_3;
      slots_3_endTag_3 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_3 | instructionFinished_3_3;
      slots_3_endTag_4 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_4 | instructionFinished_4_3;
      slots_3_endTag_5 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_5 | instructionFinished_5_3;
      slots_3_endTag_6 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_6 | instructionFinished_6_3;
      slots_3_endTag_7 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_7 | instructionFinished_7_3;
      slots_3_endTag_8 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_8 | instructionFinished_8_3;
      slots_3_endTag_9 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_9 | instructionFinished_9_3;
      slots_3_endTag_10 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_10 | instructionFinished_10_3;
      slots_3_endTag_11 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_11 | instructionFinished_11_3;
      slots_3_endTag_12 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_12 | instructionFinished_12_3;
      slots_3_endTag_13 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_13 | instructionFinished_13_3;
      slots_3_endTag_14 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_14 | instructionFinished_14_3;
      slots_3_endTag_15 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_15 | instructionFinished_15_3;
      slots_3_endTag_16 <= instructionToSlotOH[3] ? ~isLoadStoreType : slots_3_endTag_16 | slots_lsuFinished_3;
      slots_3_vxsat <= ~(instructionToSlotOH[3]) & (slots_vxsatUpdate_3 | slots_3_vxsat);
      releasePipe_pipe_v <= laneVec_0_laneRequest_bits_issueInst;
      if (validSource_valid ^ releasePipe_pipe_out_valid)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (shifterValid) begin
        shifterReg_0_valid <= validSource_valid;
        shifterReg_0_bits_instructionIndex <= validSource_bits_instructionIndex;
        shifterReg_0_bits_decodeResult_orderReduce <= validSource_bits_decodeResult_orderReduce;
        shifterReg_0_bits_decodeResult_floatMul <= validSource_bits_decodeResult_floatMul;
        shifterReg_0_bits_decodeResult_fpExecutionType <= validSource_bits_decodeResult_fpExecutionType;
        shifterReg_0_bits_decodeResult_float <= validSource_bits_decodeResult_float;
        shifterReg_0_bits_decodeResult_specialSlot <= validSource_bits_decodeResult_specialSlot;
        shifterReg_0_bits_decodeResult_topUop <= validSource_bits_decodeResult_topUop;
        shifterReg_0_bits_decodeResult_popCount <= validSource_bits_decodeResult_popCount;
        shifterReg_0_bits_decodeResult_ffo <= validSource_bits_decodeResult_ffo;
        shifterReg_0_bits_decodeResult_average <= validSource_bits_decodeResult_average;
        shifterReg_0_bits_decodeResult_reverse <= validSource_bits_decodeResult_reverse;
        shifterReg_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_0_bits_decodeResult_scheduler <= validSource_bits_decodeResult_scheduler;
        shifterReg_0_bits_decodeResult_sReadVD <= validSource_bits_decodeResult_sReadVD;
        shifterReg_0_bits_decodeResult_vtype <= validSource_bits_decodeResult_vtype;
        shifterReg_0_bits_decodeResult_sWrite <= validSource_bits_decodeResult_sWrite;
        shifterReg_0_bits_decodeResult_crossRead <= validSource_bits_decodeResult_crossRead;
        shifterReg_0_bits_decodeResult_crossWrite <= validSource_bits_decodeResult_crossWrite;
        shifterReg_0_bits_decodeResult_maskUnit <= validSource_bits_decodeResult_maskUnit;
        shifterReg_0_bits_decodeResult_special <= validSource_bits_decodeResult_special;
        shifterReg_0_bits_decodeResult_saturate <= validSource_bits_decodeResult_saturate;
        shifterReg_0_bits_decodeResult_vwmacc <= validSource_bits_decodeResult_vwmacc;
        shifterReg_0_bits_decodeResult_readOnly <= validSource_bits_decodeResult_readOnly;
        shifterReg_0_bits_decodeResult_maskSource <= validSource_bits_decodeResult_maskSource;
        shifterReg_0_bits_decodeResult_maskDestination <= validSource_bits_decodeResult_maskDestination;
        shifterReg_0_bits_decodeResult_maskLogic <= validSource_bits_decodeResult_maskLogic;
        shifterReg_0_bits_decodeResult_uop <= validSource_bits_decodeResult_uop;
        shifterReg_0_bits_decodeResult_iota <= validSource_bits_decodeResult_iota;
        shifterReg_0_bits_decodeResult_mv <= validSource_bits_decodeResult_mv;
        shifterReg_0_bits_decodeResult_extend <= validSource_bits_decodeResult_extend;
        shifterReg_0_bits_decodeResult_unOrderWrite <= validSource_bits_decodeResult_unOrderWrite;
        shifterReg_0_bits_decodeResult_compress <= validSource_bits_decodeResult_compress;
        shifterReg_0_bits_decodeResult_gather16 <= validSource_bits_decodeResult_gather16;
        shifterReg_0_bits_decodeResult_gather <= validSource_bits_decodeResult_gather;
        shifterReg_0_bits_decodeResult_slid <= validSource_bits_decodeResult_slid;
        shifterReg_0_bits_decodeResult_targetRd <= validSource_bits_decodeResult_targetRd;
        shifterReg_0_bits_decodeResult_widenReduce <= validSource_bits_decodeResult_widenReduce;
        shifterReg_0_bits_decodeResult_red <= validSource_bits_decodeResult_red;
        shifterReg_0_bits_decodeResult_nr <= validSource_bits_decodeResult_nr;
        shifterReg_0_bits_decodeResult_itype <= validSource_bits_decodeResult_itype;
        shifterReg_0_bits_decodeResult_unsigned1 <= validSource_bits_decodeResult_unsigned1;
        shifterReg_0_bits_decodeResult_unsigned0 <= validSource_bits_decodeResult_unsigned0;
        shifterReg_0_bits_decodeResult_other <= validSource_bits_decodeResult_other;
        shifterReg_0_bits_decodeResult_multiCycle <= validSource_bits_decodeResult_multiCycle;
        shifterReg_0_bits_decodeResult_divider <= validSource_bits_decodeResult_divider;
        shifterReg_0_bits_decodeResult_multiplier <= validSource_bits_decodeResult_multiplier;
        shifterReg_0_bits_decodeResult_shift <= validSource_bits_decodeResult_shift;
        shifterReg_0_bits_decodeResult_adder <= validSource_bits_decodeResult_adder;
        shifterReg_0_bits_decodeResult_logic <= validSource_bits_decodeResult_logic;
        shifterReg_0_bits_loadStore <= validSource_bits_loadStore;
        shifterReg_0_bits_issueInst <= validSource_bits_issueInst;
        shifterReg_0_bits_store <= validSource_bits_store;
        shifterReg_0_bits_special <= validSource_bits_special;
        shifterReg_0_bits_lsWholeReg <= validSource_bits_lsWholeReg;
        shifterReg_0_bits_vs1 <= validSource_bits_vs1;
        shifterReg_0_bits_vs2 <= validSource_bits_vs2;
        shifterReg_0_bits_vd <= validSource_bits_vd;
        shifterReg_0_bits_loadStoreEEW <= validSource_bits_loadStoreEEW;
        shifterReg_0_bits_mask <= validSource_bits_mask;
        shifterReg_0_bits_segment <= validSource_bits_segment;
        shifterReg_0_bits_readFromScalar <= validSource_bits_readFromScalar;
        shifterReg_0_bits_csrInterface_vl <= validSource_bits_csrInterface_vl;
        shifterReg_0_bits_csrInterface_vStart <= validSource_bits_csrInterface_vStart;
        shifterReg_0_bits_csrInterface_vlmul <= validSource_bits_csrInterface_vlmul;
        shifterReg_0_bits_csrInterface_vSew <= validSource_bits_csrInterface_vSew;
        shifterReg_0_bits_csrInterface_vxrm <= validSource_bits_csrInterface_vxrm;
        shifterReg_0_bits_csrInterface_vta <= validSource_bits_csrInterface_vta;
        shifterReg_0_bits_csrInterface_vma <= validSource_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_1 <= laneVec_1_laneRequest_bits_issueInst;
      if (validSource_1_valid ^ releasePipe_pipe_out_1_valid)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (shifterValid_1) begin
        shifterReg_1_0_valid <= validSource_1_valid;
        shifterReg_1_0_bits_instructionIndex <= validSource_1_bits_instructionIndex;
        shifterReg_1_0_bits_decodeResult_orderReduce <= validSource_1_bits_decodeResult_orderReduce;
        shifterReg_1_0_bits_decodeResult_floatMul <= validSource_1_bits_decodeResult_floatMul;
        shifterReg_1_0_bits_decodeResult_fpExecutionType <= validSource_1_bits_decodeResult_fpExecutionType;
        shifterReg_1_0_bits_decodeResult_float <= validSource_1_bits_decodeResult_float;
        shifterReg_1_0_bits_decodeResult_specialSlot <= validSource_1_bits_decodeResult_specialSlot;
        shifterReg_1_0_bits_decodeResult_topUop <= validSource_1_bits_decodeResult_topUop;
        shifterReg_1_0_bits_decodeResult_popCount <= validSource_1_bits_decodeResult_popCount;
        shifterReg_1_0_bits_decodeResult_ffo <= validSource_1_bits_decodeResult_ffo;
        shifterReg_1_0_bits_decodeResult_average <= validSource_1_bits_decodeResult_average;
        shifterReg_1_0_bits_decodeResult_reverse <= validSource_1_bits_decodeResult_reverse;
        shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_1_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_1_0_bits_decodeResult_scheduler <= validSource_1_bits_decodeResult_scheduler;
        shifterReg_1_0_bits_decodeResult_sReadVD <= validSource_1_bits_decodeResult_sReadVD;
        shifterReg_1_0_bits_decodeResult_vtype <= validSource_1_bits_decodeResult_vtype;
        shifterReg_1_0_bits_decodeResult_sWrite <= validSource_1_bits_decodeResult_sWrite;
        shifterReg_1_0_bits_decodeResult_crossRead <= validSource_1_bits_decodeResult_crossRead;
        shifterReg_1_0_bits_decodeResult_crossWrite <= validSource_1_bits_decodeResult_crossWrite;
        shifterReg_1_0_bits_decodeResult_maskUnit <= validSource_1_bits_decodeResult_maskUnit;
        shifterReg_1_0_bits_decodeResult_special <= validSource_1_bits_decodeResult_special;
        shifterReg_1_0_bits_decodeResult_saturate <= validSource_1_bits_decodeResult_saturate;
        shifterReg_1_0_bits_decodeResult_vwmacc <= validSource_1_bits_decodeResult_vwmacc;
        shifterReg_1_0_bits_decodeResult_readOnly <= validSource_1_bits_decodeResult_readOnly;
        shifterReg_1_0_bits_decodeResult_maskSource <= validSource_1_bits_decodeResult_maskSource;
        shifterReg_1_0_bits_decodeResult_maskDestination <= validSource_1_bits_decodeResult_maskDestination;
        shifterReg_1_0_bits_decodeResult_maskLogic <= validSource_1_bits_decodeResult_maskLogic;
        shifterReg_1_0_bits_decodeResult_uop <= validSource_1_bits_decodeResult_uop;
        shifterReg_1_0_bits_decodeResult_iota <= validSource_1_bits_decodeResult_iota;
        shifterReg_1_0_bits_decodeResult_mv <= validSource_1_bits_decodeResult_mv;
        shifterReg_1_0_bits_decodeResult_extend <= validSource_1_bits_decodeResult_extend;
        shifterReg_1_0_bits_decodeResult_unOrderWrite <= validSource_1_bits_decodeResult_unOrderWrite;
        shifterReg_1_0_bits_decodeResult_compress <= validSource_1_bits_decodeResult_compress;
        shifterReg_1_0_bits_decodeResult_gather16 <= validSource_1_bits_decodeResult_gather16;
        shifterReg_1_0_bits_decodeResult_gather <= validSource_1_bits_decodeResult_gather;
        shifterReg_1_0_bits_decodeResult_slid <= validSource_1_bits_decodeResult_slid;
        shifterReg_1_0_bits_decodeResult_targetRd <= validSource_1_bits_decodeResult_targetRd;
        shifterReg_1_0_bits_decodeResult_widenReduce <= validSource_1_bits_decodeResult_widenReduce;
        shifterReg_1_0_bits_decodeResult_red <= validSource_1_bits_decodeResult_red;
        shifterReg_1_0_bits_decodeResult_nr <= validSource_1_bits_decodeResult_nr;
        shifterReg_1_0_bits_decodeResult_itype <= validSource_1_bits_decodeResult_itype;
        shifterReg_1_0_bits_decodeResult_unsigned1 <= validSource_1_bits_decodeResult_unsigned1;
        shifterReg_1_0_bits_decodeResult_unsigned0 <= validSource_1_bits_decodeResult_unsigned0;
        shifterReg_1_0_bits_decodeResult_other <= validSource_1_bits_decodeResult_other;
        shifterReg_1_0_bits_decodeResult_multiCycle <= validSource_1_bits_decodeResult_multiCycle;
        shifterReg_1_0_bits_decodeResult_divider <= validSource_1_bits_decodeResult_divider;
        shifterReg_1_0_bits_decodeResult_multiplier <= validSource_1_bits_decodeResult_multiplier;
        shifterReg_1_0_bits_decodeResult_shift <= validSource_1_bits_decodeResult_shift;
        shifterReg_1_0_bits_decodeResult_adder <= validSource_1_bits_decodeResult_adder;
        shifterReg_1_0_bits_decodeResult_logic <= validSource_1_bits_decodeResult_logic;
        shifterReg_1_0_bits_loadStore <= validSource_1_bits_loadStore;
        shifterReg_1_0_bits_issueInst <= validSource_1_bits_issueInst;
        shifterReg_1_0_bits_store <= validSource_1_bits_store;
        shifterReg_1_0_bits_special <= validSource_1_bits_special;
        shifterReg_1_0_bits_lsWholeReg <= validSource_1_bits_lsWholeReg;
        shifterReg_1_0_bits_vs1 <= validSource_1_bits_vs1;
        shifterReg_1_0_bits_vs2 <= validSource_1_bits_vs2;
        shifterReg_1_0_bits_vd <= validSource_1_bits_vd;
        shifterReg_1_0_bits_loadStoreEEW <= validSource_1_bits_loadStoreEEW;
        shifterReg_1_0_bits_mask <= validSource_1_bits_mask;
        shifterReg_1_0_bits_segment <= validSource_1_bits_segment;
        shifterReg_1_0_bits_readFromScalar <= validSource_1_bits_readFromScalar;
        shifterReg_1_0_bits_csrInterface_vl <= validSource_1_bits_csrInterface_vl;
        shifterReg_1_0_bits_csrInterface_vStart <= validSource_1_bits_csrInterface_vStart;
        shifterReg_1_0_bits_csrInterface_vlmul <= validSource_1_bits_csrInterface_vlmul;
        shifterReg_1_0_bits_csrInterface_vSew <= validSource_1_bits_csrInterface_vSew;
        shifterReg_1_0_bits_csrInterface_vxrm <= validSource_1_bits_csrInterface_vxrm;
        shifterReg_1_0_bits_csrInterface_vta <= validSource_1_bits_csrInterface_vta;
        shifterReg_1_0_bits_csrInterface_vma <= validSource_1_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_2 <= laneVec_2_laneRequest_bits_issueInst;
      if (validSource_2_valid ^ releasePipe_pipe_out_2_valid)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (shifterValid_2) begin
        shifterReg_2_0_valid <= validSource_2_valid;
        shifterReg_2_0_bits_instructionIndex <= validSource_2_bits_instructionIndex;
        shifterReg_2_0_bits_decodeResult_orderReduce <= validSource_2_bits_decodeResult_orderReduce;
        shifterReg_2_0_bits_decodeResult_floatMul <= validSource_2_bits_decodeResult_floatMul;
        shifterReg_2_0_bits_decodeResult_fpExecutionType <= validSource_2_bits_decodeResult_fpExecutionType;
        shifterReg_2_0_bits_decodeResult_float <= validSource_2_bits_decodeResult_float;
        shifterReg_2_0_bits_decodeResult_specialSlot <= validSource_2_bits_decodeResult_specialSlot;
        shifterReg_2_0_bits_decodeResult_topUop <= validSource_2_bits_decodeResult_topUop;
        shifterReg_2_0_bits_decodeResult_popCount <= validSource_2_bits_decodeResult_popCount;
        shifterReg_2_0_bits_decodeResult_ffo <= validSource_2_bits_decodeResult_ffo;
        shifterReg_2_0_bits_decodeResult_average <= validSource_2_bits_decodeResult_average;
        shifterReg_2_0_bits_decodeResult_reverse <= validSource_2_bits_decodeResult_reverse;
        shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_2_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_2_0_bits_decodeResult_scheduler <= validSource_2_bits_decodeResult_scheduler;
        shifterReg_2_0_bits_decodeResult_sReadVD <= validSource_2_bits_decodeResult_sReadVD;
        shifterReg_2_0_bits_decodeResult_vtype <= validSource_2_bits_decodeResult_vtype;
        shifterReg_2_0_bits_decodeResult_sWrite <= validSource_2_bits_decodeResult_sWrite;
        shifterReg_2_0_bits_decodeResult_crossRead <= validSource_2_bits_decodeResult_crossRead;
        shifterReg_2_0_bits_decodeResult_crossWrite <= validSource_2_bits_decodeResult_crossWrite;
        shifterReg_2_0_bits_decodeResult_maskUnit <= validSource_2_bits_decodeResult_maskUnit;
        shifterReg_2_0_bits_decodeResult_special <= validSource_2_bits_decodeResult_special;
        shifterReg_2_0_bits_decodeResult_saturate <= validSource_2_bits_decodeResult_saturate;
        shifterReg_2_0_bits_decodeResult_vwmacc <= validSource_2_bits_decodeResult_vwmacc;
        shifterReg_2_0_bits_decodeResult_readOnly <= validSource_2_bits_decodeResult_readOnly;
        shifterReg_2_0_bits_decodeResult_maskSource <= validSource_2_bits_decodeResult_maskSource;
        shifterReg_2_0_bits_decodeResult_maskDestination <= validSource_2_bits_decodeResult_maskDestination;
        shifterReg_2_0_bits_decodeResult_maskLogic <= validSource_2_bits_decodeResult_maskLogic;
        shifterReg_2_0_bits_decodeResult_uop <= validSource_2_bits_decodeResult_uop;
        shifterReg_2_0_bits_decodeResult_iota <= validSource_2_bits_decodeResult_iota;
        shifterReg_2_0_bits_decodeResult_mv <= validSource_2_bits_decodeResult_mv;
        shifterReg_2_0_bits_decodeResult_extend <= validSource_2_bits_decodeResult_extend;
        shifterReg_2_0_bits_decodeResult_unOrderWrite <= validSource_2_bits_decodeResult_unOrderWrite;
        shifterReg_2_0_bits_decodeResult_compress <= validSource_2_bits_decodeResult_compress;
        shifterReg_2_0_bits_decodeResult_gather16 <= validSource_2_bits_decodeResult_gather16;
        shifterReg_2_0_bits_decodeResult_gather <= validSource_2_bits_decodeResult_gather;
        shifterReg_2_0_bits_decodeResult_slid <= validSource_2_bits_decodeResult_slid;
        shifterReg_2_0_bits_decodeResult_targetRd <= validSource_2_bits_decodeResult_targetRd;
        shifterReg_2_0_bits_decodeResult_widenReduce <= validSource_2_bits_decodeResult_widenReduce;
        shifterReg_2_0_bits_decodeResult_red <= validSource_2_bits_decodeResult_red;
        shifterReg_2_0_bits_decodeResult_nr <= validSource_2_bits_decodeResult_nr;
        shifterReg_2_0_bits_decodeResult_itype <= validSource_2_bits_decodeResult_itype;
        shifterReg_2_0_bits_decodeResult_unsigned1 <= validSource_2_bits_decodeResult_unsigned1;
        shifterReg_2_0_bits_decodeResult_unsigned0 <= validSource_2_bits_decodeResult_unsigned0;
        shifterReg_2_0_bits_decodeResult_other <= validSource_2_bits_decodeResult_other;
        shifterReg_2_0_bits_decodeResult_multiCycle <= validSource_2_bits_decodeResult_multiCycle;
        shifterReg_2_0_bits_decodeResult_divider <= validSource_2_bits_decodeResult_divider;
        shifterReg_2_0_bits_decodeResult_multiplier <= validSource_2_bits_decodeResult_multiplier;
        shifterReg_2_0_bits_decodeResult_shift <= validSource_2_bits_decodeResult_shift;
        shifterReg_2_0_bits_decodeResult_adder <= validSource_2_bits_decodeResult_adder;
        shifterReg_2_0_bits_decodeResult_logic <= validSource_2_bits_decodeResult_logic;
        shifterReg_2_0_bits_loadStore <= validSource_2_bits_loadStore;
        shifterReg_2_0_bits_issueInst <= validSource_2_bits_issueInst;
        shifterReg_2_0_bits_store <= validSource_2_bits_store;
        shifterReg_2_0_bits_special <= validSource_2_bits_special;
        shifterReg_2_0_bits_lsWholeReg <= validSource_2_bits_lsWholeReg;
        shifterReg_2_0_bits_vs1 <= validSource_2_bits_vs1;
        shifterReg_2_0_bits_vs2 <= validSource_2_bits_vs2;
        shifterReg_2_0_bits_vd <= validSource_2_bits_vd;
        shifterReg_2_0_bits_loadStoreEEW <= validSource_2_bits_loadStoreEEW;
        shifterReg_2_0_bits_mask <= validSource_2_bits_mask;
        shifterReg_2_0_bits_segment <= validSource_2_bits_segment;
        shifterReg_2_0_bits_readFromScalar <= validSource_2_bits_readFromScalar;
        shifterReg_2_0_bits_csrInterface_vl <= validSource_2_bits_csrInterface_vl;
        shifterReg_2_0_bits_csrInterface_vStart <= validSource_2_bits_csrInterface_vStart;
        shifterReg_2_0_bits_csrInterface_vlmul <= validSource_2_bits_csrInterface_vlmul;
        shifterReg_2_0_bits_csrInterface_vSew <= validSource_2_bits_csrInterface_vSew;
        shifterReg_2_0_bits_csrInterface_vxrm <= validSource_2_bits_csrInterface_vxrm;
        shifterReg_2_0_bits_csrInterface_vta <= validSource_2_bits_csrInterface_vta;
        shifterReg_2_0_bits_csrInterface_vma <= validSource_2_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_3 <= laneVec_3_laneRequest_bits_issueInst;
      if (validSource_3_valid ^ releasePipe_pipe_out_3_valid)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (shifterValid_3) begin
        shifterReg_3_0_valid <= validSource_3_valid;
        shifterReg_3_0_bits_instructionIndex <= validSource_3_bits_instructionIndex;
        shifterReg_3_0_bits_decodeResult_orderReduce <= validSource_3_bits_decodeResult_orderReduce;
        shifterReg_3_0_bits_decodeResult_floatMul <= validSource_3_bits_decodeResult_floatMul;
        shifterReg_3_0_bits_decodeResult_fpExecutionType <= validSource_3_bits_decodeResult_fpExecutionType;
        shifterReg_3_0_bits_decodeResult_float <= validSource_3_bits_decodeResult_float;
        shifterReg_3_0_bits_decodeResult_specialSlot <= validSource_3_bits_decodeResult_specialSlot;
        shifterReg_3_0_bits_decodeResult_topUop <= validSource_3_bits_decodeResult_topUop;
        shifterReg_3_0_bits_decodeResult_popCount <= validSource_3_bits_decodeResult_popCount;
        shifterReg_3_0_bits_decodeResult_ffo <= validSource_3_bits_decodeResult_ffo;
        shifterReg_3_0_bits_decodeResult_average <= validSource_3_bits_decodeResult_average;
        shifterReg_3_0_bits_decodeResult_reverse <= validSource_3_bits_decodeResult_reverse;
        shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_3_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_3_0_bits_decodeResult_scheduler <= validSource_3_bits_decodeResult_scheduler;
        shifterReg_3_0_bits_decodeResult_sReadVD <= validSource_3_bits_decodeResult_sReadVD;
        shifterReg_3_0_bits_decodeResult_vtype <= validSource_3_bits_decodeResult_vtype;
        shifterReg_3_0_bits_decodeResult_sWrite <= validSource_3_bits_decodeResult_sWrite;
        shifterReg_3_0_bits_decodeResult_crossRead <= validSource_3_bits_decodeResult_crossRead;
        shifterReg_3_0_bits_decodeResult_crossWrite <= validSource_3_bits_decodeResult_crossWrite;
        shifterReg_3_0_bits_decodeResult_maskUnit <= validSource_3_bits_decodeResult_maskUnit;
        shifterReg_3_0_bits_decodeResult_special <= validSource_3_bits_decodeResult_special;
        shifterReg_3_0_bits_decodeResult_saturate <= validSource_3_bits_decodeResult_saturate;
        shifterReg_3_0_bits_decodeResult_vwmacc <= validSource_3_bits_decodeResult_vwmacc;
        shifterReg_3_0_bits_decodeResult_readOnly <= validSource_3_bits_decodeResult_readOnly;
        shifterReg_3_0_bits_decodeResult_maskSource <= validSource_3_bits_decodeResult_maskSource;
        shifterReg_3_0_bits_decodeResult_maskDestination <= validSource_3_bits_decodeResult_maskDestination;
        shifterReg_3_0_bits_decodeResult_maskLogic <= validSource_3_bits_decodeResult_maskLogic;
        shifterReg_3_0_bits_decodeResult_uop <= validSource_3_bits_decodeResult_uop;
        shifterReg_3_0_bits_decodeResult_iota <= validSource_3_bits_decodeResult_iota;
        shifterReg_3_0_bits_decodeResult_mv <= validSource_3_bits_decodeResult_mv;
        shifterReg_3_0_bits_decodeResult_extend <= validSource_3_bits_decodeResult_extend;
        shifterReg_3_0_bits_decodeResult_unOrderWrite <= validSource_3_bits_decodeResult_unOrderWrite;
        shifterReg_3_0_bits_decodeResult_compress <= validSource_3_bits_decodeResult_compress;
        shifterReg_3_0_bits_decodeResult_gather16 <= validSource_3_bits_decodeResult_gather16;
        shifterReg_3_0_bits_decodeResult_gather <= validSource_3_bits_decodeResult_gather;
        shifterReg_3_0_bits_decodeResult_slid <= validSource_3_bits_decodeResult_slid;
        shifterReg_3_0_bits_decodeResult_targetRd <= validSource_3_bits_decodeResult_targetRd;
        shifterReg_3_0_bits_decodeResult_widenReduce <= validSource_3_bits_decodeResult_widenReduce;
        shifterReg_3_0_bits_decodeResult_red <= validSource_3_bits_decodeResult_red;
        shifterReg_3_0_bits_decodeResult_nr <= validSource_3_bits_decodeResult_nr;
        shifterReg_3_0_bits_decodeResult_itype <= validSource_3_bits_decodeResult_itype;
        shifterReg_3_0_bits_decodeResult_unsigned1 <= validSource_3_bits_decodeResult_unsigned1;
        shifterReg_3_0_bits_decodeResult_unsigned0 <= validSource_3_bits_decodeResult_unsigned0;
        shifterReg_3_0_bits_decodeResult_other <= validSource_3_bits_decodeResult_other;
        shifterReg_3_0_bits_decodeResult_multiCycle <= validSource_3_bits_decodeResult_multiCycle;
        shifterReg_3_0_bits_decodeResult_divider <= validSource_3_bits_decodeResult_divider;
        shifterReg_3_0_bits_decodeResult_multiplier <= validSource_3_bits_decodeResult_multiplier;
        shifterReg_3_0_bits_decodeResult_shift <= validSource_3_bits_decodeResult_shift;
        shifterReg_3_0_bits_decodeResult_adder <= validSource_3_bits_decodeResult_adder;
        shifterReg_3_0_bits_decodeResult_logic <= validSource_3_bits_decodeResult_logic;
        shifterReg_3_0_bits_loadStore <= validSource_3_bits_loadStore;
        shifterReg_3_0_bits_issueInst <= validSource_3_bits_issueInst;
        shifterReg_3_0_bits_store <= validSource_3_bits_store;
        shifterReg_3_0_bits_special <= validSource_3_bits_special;
        shifterReg_3_0_bits_lsWholeReg <= validSource_3_bits_lsWholeReg;
        shifterReg_3_0_bits_vs1 <= validSource_3_bits_vs1;
        shifterReg_3_0_bits_vs2 <= validSource_3_bits_vs2;
        shifterReg_3_0_bits_vd <= validSource_3_bits_vd;
        shifterReg_3_0_bits_loadStoreEEW <= validSource_3_bits_loadStoreEEW;
        shifterReg_3_0_bits_mask <= validSource_3_bits_mask;
        shifterReg_3_0_bits_segment <= validSource_3_bits_segment;
        shifterReg_3_0_bits_readFromScalar <= validSource_3_bits_readFromScalar;
        shifterReg_3_0_bits_csrInterface_vl <= validSource_3_bits_csrInterface_vl;
        shifterReg_3_0_bits_csrInterface_vStart <= validSource_3_bits_csrInterface_vStart;
        shifterReg_3_0_bits_csrInterface_vlmul <= validSource_3_bits_csrInterface_vlmul;
        shifterReg_3_0_bits_csrInterface_vSew <= validSource_3_bits_csrInterface_vSew;
        shifterReg_3_0_bits_csrInterface_vxrm <= validSource_3_bits_csrInterface_vxrm;
        shifterReg_3_0_bits_csrInterface_vta <= validSource_3_bits_csrInterface_vta;
        shifterReg_3_0_bits_csrInterface_vma <= validSource_3_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_4 <= laneVec_4_laneRequest_bits_issueInst;
      if (validSource_4_valid ^ releasePipe_pipe_out_4_valid)
        tokenCheck_counter_4 <= tokenCheck_counter_4 + tokenCheck_counterChange_4;
      if (shifterValid_4) begin
        shifterReg_4_0_valid <= validSource_4_valid;
        shifterReg_4_0_bits_instructionIndex <= validSource_4_bits_instructionIndex;
        shifterReg_4_0_bits_decodeResult_orderReduce <= validSource_4_bits_decodeResult_orderReduce;
        shifterReg_4_0_bits_decodeResult_floatMul <= validSource_4_bits_decodeResult_floatMul;
        shifterReg_4_0_bits_decodeResult_fpExecutionType <= validSource_4_bits_decodeResult_fpExecutionType;
        shifterReg_4_0_bits_decodeResult_float <= validSource_4_bits_decodeResult_float;
        shifterReg_4_0_bits_decodeResult_specialSlot <= validSource_4_bits_decodeResult_specialSlot;
        shifterReg_4_0_bits_decodeResult_topUop <= validSource_4_bits_decodeResult_topUop;
        shifterReg_4_0_bits_decodeResult_popCount <= validSource_4_bits_decodeResult_popCount;
        shifterReg_4_0_bits_decodeResult_ffo <= validSource_4_bits_decodeResult_ffo;
        shifterReg_4_0_bits_decodeResult_average <= validSource_4_bits_decodeResult_average;
        shifterReg_4_0_bits_decodeResult_reverse <= validSource_4_bits_decodeResult_reverse;
        shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_4_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_4_0_bits_decodeResult_scheduler <= validSource_4_bits_decodeResult_scheduler;
        shifterReg_4_0_bits_decodeResult_sReadVD <= validSource_4_bits_decodeResult_sReadVD;
        shifterReg_4_0_bits_decodeResult_vtype <= validSource_4_bits_decodeResult_vtype;
        shifterReg_4_0_bits_decodeResult_sWrite <= validSource_4_bits_decodeResult_sWrite;
        shifterReg_4_0_bits_decodeResult_crossRead <= validSource_4_bits_decodeResult_crossRead;
        shifterReg_4_0_bits_decodeResult_crossWrite <= validSource_4_bits_decodeResult_crossWrite;
        shifterReg_4_0_bits_decodeResult_maskUnit <= validSource_4_bits_decodeResult_maskUnit;
        shifterReg_4_0_bits_decodeResult_special <= validSource_4_bits_decodeResult_special;
        shifterReg_4_0_bits_decodeResult_saturate <= validSource_4_bits_decodeResult_saturate;
        shifterReg_4_0_bits_decodeResult_vwmacc <= validSource_4_bits_decodeResult_vwmacc;
        shifterReg_4_0_bits_decodeResult_readOnly <= validSource_4_bits_decodeResult_readOnly;
        shifterReg_4_0_bits_decodeResult_maskSource <= validSource_4_bits_decodeResult_maskSource;
        shifterReg_4_0_bits_decodeResult_maskDestination <= validSource_4_bits_decodeResult_maskDestination;
        shifterReg_4_0_bits_decodeResult_maskLogic <= validSource_4_bits_decodeResult_maskLogic;
        shifterReg_4_0_bits_decodeResult_uop <= validSource_4_bits_decodeResult_uop;
        shifterReg_4_0_bits_decodeResult_iota <= validSource_4_bits_decodeResult_iota;
        shifterReg_4_0_bits_decodeResult_mv <= validSource_4_bits_decodeResult_mv;
        shifterReg_4_0_bits_decodeResult_extend <= validSource_4_bits_decodeResult_extend;
        shifterReg_4_0_bits_decodeResult_unOrderWrite <= validSource_4_bits_decodeResult_unOrderWrite;
        shifterReg_4_0_bits_decodeResult_compress <= validSource_4_bits_decodeResult_compress;
        shifterReg_4_0_bits_decodeResult_gather16 <= validSource_4_bits_decodeResult_gather16;
        shifterReg_4_0_bits_decodeResult_gather <= validSource_4_bits_decodeResult_gather;
        shifterReg_4_0_bits_decodeResult_slid <= validSource_4_bits_decodeResult_slid;
        shifterReg_4_0_bits_decodeResult_targetRd <= validSource_4_bits_decodeResult_targetRd;
        shifterReg_4_0_bits_decodeResult_widenReduce <= validSource_4_bits_decodeResult_widenReduce;
        shifterReg_4_0_bits_decodeResult_red <= validSource_4_bits_decodeResult_red;
        shifterReg_4_0_bits_decodeResult_nr <= validSource_4_bits_decodeResult_nr;
        shifterReg_4_0_bits_decodeResult_itype <= validSource_4_bits_decodeResult_itype;
        shifterReg_4_0_bits_decodeResult_unsigned1 <= validSource_4_bits_decodeResult_unsigned1;
        shifterReg_4_0_bits_decodeResult_unsigned0 <= validSource_4_bits_decodeResult_unsigned0;
        shifterReg_4_0_bits_decodeResult_other <= validSource_4_bits_decodeResult_other;
        shifterReg_4_0_bits_decodeResult_multiCycle <= validSource_4_bits_decodeResult_multiCycle;
        shifterReg_4_0_bits_decodeResult_divider <= validSource_4_bits_decodeResult_divider;
        shifterReg_4_0_bits_decodeResult_multiplier <= validSource_4_bits_decodeResult_multiplier;
        shifterReg_4_0_bits_decodeResult_shift <= validSource_4_bits_decodeResult_shift;
        shifterReg_4_0_bits_decodeResult_adder <= validSource_4_bits_decodeResult_adder;
        shifterReg_4_0_bits_decodeResult_logic <= validSource_4_bits_decodeResult_logic;
        shifterReg_4_0_bits_loadStore <= validSource_4_bits_loadStore;
        shifterReg_4_0_bits_issueInst <= validSource_4_bits_issueInst;
        shifterReg_4_0_bits_store <= validSource_4_bits_store;
        shifterReg_4_0_bits_special <= validSource_4_bits_special;
        shifterReg_4_0_bits_lsWholeReg <= validSource_4_bits_lsWholeReg;
        shifterReg_4_0_bits_vs1 <= validSource_4_bits_vs1;
        shifterReg_4_0_bits_vs2 <= validSource_4_bits_vs2;
        shifterReg_4_0_bits_vd <= validSource_4_bits_vd;
        shifterReg_4_0_bits_loadStoreEEW <= validSource_4_bits_loadStoreEEW;
        shifterReg_4_0_bits_mask <= validSource_4_bits_mask;
        shifterReg_4_0_bits_segment <= validSource_4_bits_segment;
        shifterReg_4_0_bits_readFromScalar <= validSource_4_bits_readFromScalar;
        shifterReg_4_0_bits_csrInterface_vl <= validSource_4_bits_csrInterface_vl;
        shifterReg_4_0_bits_csrInterface_vStart <= validSource_4_bits_csrInterface_vStart;
        shifterReg_4_0_bits_csrInterface_vlmul <= validSource_4_bits_csrInterface_vlmul;
        shifterReg_4_0_bits_csrInterface_vSew <= validSource_4_bits_csrInterface_vSew;
        shifterReg_4_0_bits_csrInterface_vxrm <= validSource_4_bits_csrInterface_vxrm;
        shifterReg_4_0_bits_csrInterface_vta <= validSource_4_bits_csrInterface_vta;
        shifterReg_4_0_bits_csrInterface_vma <= validSource_4_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_5 <= laneVec_5_laneRequest_bits_issueInst;
      if (validSource_5_valid ^ releasePipe_pipe_out_5_valid)
        tokenCheck_counter_5 <= tokenCheck_counter_5 + tokenCheck_counterChange_5;
      if (shifterValid_5) begin
        shifterReg_5_0_valid <= validSource_5_valid;
        shifterReg_5_0_bits_instructionIndex <= validSource_5_bits_instructionIndex;
        shifterReg_5_0_bits_decodeResult_orderReduce <= validSource_5_bits_decodeResult_orderReduce;
        shifterReg_5_0_bits_decodeResult_floatMul <= validSource_5_bits_decodeResult_floatMul;
        shifterReg_5_0_bits_decodeResult_fpExecutionType <= validSource_5_bits_decodeResult_fpExecutionType;
        shifterReg_5_0_bits_decodeResult_float <= validSource_5_bits_decodeResult_float;
        shifterReg_5_0_bits_decodeResult_specialSlot <= validSource_5_bits_decodeResult_specialSlot;
        shifterReg_5_0_bits_decodeResult_topUop <= validSource_5_bits_decodeResult_topUop;
        shifterReg_5_0_bits_decodeResult_popCount <= validSource_5_bits_decodeResult_popCount;
        shifterReg_5_0_bits_decodeResult_ffo <= validSource_5_bits_decodeResult_ffo;
        shifterReg_5_0_bits_decodeResult_average <= validSource_5_bits_decodeResult_average;
        shifterReg_5_0_bits_decodeResult_reverse <= validSource_5_bits_decodeResult_reverse;
        shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_5_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_5_0_bits_decodeResult_scheduler <= validSource_5_bits_decodeResult_scheduler;
        shifterReg_5_0_bits_decodeResult_sReadVD <= validSource_5_bits_decodeResult_sReadVD;
        shifterReg_5_0_bits_decodeResult_vtype <= validSource_5_bits_decodeResult_vtype;
        shifterReg_5_0_bits_decodeResult_sWrite <= validSource_5_bits_decodeResult_sWrite;
        shifterReg_5_0_bits_decodeResult_crossRead <= validSource_5_bits_decodeResult_crossRead;
        shifterReg_5_0_bits_decodeResult_crossWrite <= validSource_5_bits_decodeResult_crossWrite;
        shifterReg_5_0_bits_decodeResult_maskUnit <= validSource_5_bits_decodeResult_maskUnit;
        shifterReg_5_0_bits_decodeResult_special <= validSource_5_bits_decodeResult_special;
        shifterReg_5_0_bits_decodeResult_saturate <= validSource_5_bits_decodeResult_saturate;
        shifterReg_5_0_bits_decodeResult_vwmacc <= validSource_5_bits_decodeResult_vwmacc;
        shifterReg_5_0_bits_decodeResult_readOnly <= validSource_5_bits_decodeResult_readOnly;
        shifterReg_5_0_bits_decodeResult_maskSource <= validSource_5_bits_decodeResult_maskSource;
        shifterReg_5_0_bits_decodeResult_maskDestination <= validSource_5_bits_decodeResult_maskDestination;
        shifterReg_5_0_bits_decodeResult_maskLogic <= validSource_5_bits_decodeResult_maskLogic;
        shifterReg_5_0_bits_decodeResult_uop <= validSource_5_bits_decodeResult_uop;
        shifterReg_5_0_bits_decodeResult_iota <= validSource_5_bits_decodeResult_iota;
        shifterReg_5_0_bits_decodeResult_mv <= validSource_5_bits_decodeResult_mv;
        shifterReg_5_0_bits_decodeResult_extend <= validSource_5_bits_decodeResult_extend;
        shifterReg_5_0_bits_decodeResult_unOrderWrite <= validSource_5_bits_decodeResult_unOrderWrite;
        shifterReg_5_0_bits_decodeResult_compress <= validSource_5_bits_decodeResult_compress;
        shifterReg_5_0_bits_decodeResult_gather16 <= validSource_5_bits_decodeResult_gather16;
        shifterReg_5_0_bits_decodeResult_gather <= validSource_5_bits_decodeResult_gather;
        shifterReg_5_0_bits_decodeResult_slid <= validSource_5_bits_decodeResult_slid;
        shifterReg_5_0_bits_decodeResult_targetRd <= validSource_5_bits_decodeResult_targetRd;
        shifterReg_5_0_bits_decodeResult_widenReduce <= validSource_5_bits_decodeResult_widenReduce;
        shifterReg_5_0_bits_decodeResult_red <= validSource_5_bits_decodeResult_red;
        shifterReg_5_0_bits_decodeResult_nr <= validSource_5_bits_decodeResult_nr;
        shifterReg_5_0_bits_decodeResult_itype <= validSource_5_bits_decodeResult_itype;
        shifterReg_5_0_bits_decodeResult_unsigned1 <= validSource_5_bits_decodeResult_unsigned1;
        shifterReg_5_0_bits_decodeResult_unsigned0 <= validSource_5_bits_decodeResult_unsigned0;
        shifterReg_5_0_bits_decodeResult_other <= validSource_5_bits_decodeResult_other;
        shifterReg_5_0_bits_decodeResult_multiCycle <= validSource_5_bits_decodeResult_multiCycle;
        shifterReg_5_0_bits_decodeResult_divider <= validSource_5_bits_decodeResult_divider;
        shifterReg_5_0_bits_decodeResult_multiplier <= validSource_5_bits_decodeResult_multiplier;
        shifterReg_5_0_bits_decodeResult_shift <= validSource_5_bits_decodeResult_shift;
        shifterReg_5_0_bits_decodeResult_adder <= validSource_5_bits_decodeResult_adder;
        shifterReg_5_0_bits_decodeResult_logic <= validSource_5_bits_decodeResult_logic;
        shifterReg_5_0_bits_loadStore <= validSource_5_bits_loadStore;
        shifterReg_5_0_bits_issueInst <= validSource_5_bits_issueInst;
        shifterReg_5_0_bits_store <= validSource_5_bits_store;
        shifterReg_5_0_bits_special <= validSource_5_bits_special;
        shifterReg_5_0_bits_lsWholeReg <= validSource_5_bits_lsWholeReg;
        shifterReg_5_0_bits_vs1 <= validSource_5_bits_vs1;
        shifterReg_5_0_bits_vs2 <= validSource_5_bits_vs2;
        shifterReg_5_0_bits_vd <= validSource_5_bits_vd;
        shifterReg_5_0_bits_loadStoreEEW <= validSource_5_bits_loadStoreEEW;
        shifterReg_5_0_bits_mask <= validSource_5_bits_mask;
        shifterReg_5_0_bits_segment <= validSource_5_bits_segment;
        shifterReg_5_0_bits_readFromScalar <= validSource_5_bits_readFromScalar;
        shifterReg_5_0_bits_csrInterface_vl <= validSource_5_bits_csrInterface_vl;
        shifterReg_5_0_bits_csrInterface_vStart <= validSource_5_bits_csrInterface_vStart;
        shifterReg_5_0_bits_csrInterface_vlmul <= validSource_5_bits_csrInterface_vlmul;
        shifterReg_5_0_bits_csrInterface_vSew <= validSource_5_bits_csrInterface_vSew;
        shifterReg_5_0_bits_csrInterface_vxrm <= validSource_5_bits_csrInterface_vxrm;
        shifterReg_5_0_bits_csrInterface_vta <= validSource_5_bits_csrInterface_vta;
        shifterReg_5_0_bits_csrInterface_vma <= validSource_5_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_6 <= laneVec_6_laneRequest_bits_issueInst;
      if (validSource_6_valid ^ releasePipe_pipe_out_6_valid)
        tokenCheck_counter_6 <= tokenCheck_counter_6 + tokenCheck_counterChange_6;
      if (shifterValid_6) begin
        shifterReg_6_0_valid <= validSource_6_valid;
        shifterReg_6_0_bits_instructionIndex <= validSource_6_bits_instructionIndex;
        shifterReg_6_0_bits_decodeResult_orderReduce <= validSource_6_bits_decodeResult_orderReduce;
        shifterReg_6_0_bits_decodeResult_floatMul <= validSource_6_bits_decodeResult_floatMul;
        shifterReg_6_0_bits_decodeResult_fpExecutionType <= validSource_6_bits_decodeResult_fpExecutionType;
        shifterReg_6_0_bits_decodeResult_float <= validSource_6_bits_decodeResult_float;
        shifterReg_6_0_bits_decodeResult_specialSlot <= validSource_6_bits_decodeResult_specialSlot;
        shifterReg_6_0_bits_decodeResult_topUop <= validSource_6_bits_decodeResult_topUop;
        shifterReg_6_0_bits_decodeResult_popCount <= validSource_6_bits_decodeResult_popCount;
        shifterReg_6_0_bits_decodeResult_ffo <= validSource_6_bits_decodeResult_ffo;
        shifterReg_6_0_bits_decodeResult_average <= validSource_6_bits_decodeResult_average;
        shifterReg_6_0_bits_decodeResult_reverse <= validSource_6_bits_decodeResult_reverse;
        shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_6_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_6_0_bits_decodeResult_scheduler <= validSource_6_bits_decodeResult_scheduler;
        shifterReg_6_0_bits_decodeResult_sReadVD <= validSource_6_bits_decodeResult_sReadVD;
        shifterReg_6_0_bits_decodeResult_vtype <= validSource_6_bits_decodeResult_vtype;
        shifterReg_6_0_bits_decodeResult_sWrite <= validSource_6_bits_decodeResult_sWrite;
        shifterReg_6_0_bits_decodeResult_crossRead <= validSource_6_bits_decodeResult_crossRead;
        shifterReg_6_0_bits_decodeResult_crossWrite <= validSource_6_bits_decodeResult_crossWrite;
        shifterReg_6_0_bits_decodeResult_maskUnit <= validSource_6_bits_decodeResult_maskUnit;
        shifterReg_6_0_bits_decodeResult_special <= validSource_6_bits_decodeResult_special;
        shifterReg_6_0_bits_decodeResult_saturate <= validSource_6_bits_decodeResult_saturate;
        shifterReg_6_0_bits_decodeResult_vwmacc <= validSource_6_bits_decodeResult_vwmacc;
        shifterReg_6_0_bits_decodeResult_readOnly <= validSource_6_bits_decodeResult_readOnly;
        shifterReg_6_0_bits_decodeResult_maskSource <= validSource_6_bits_decodeResult_maskSource;
        shifterReg_6_0_bits_decodeResult_maskDestination <= validSource_6_bits_decodeResult_maskDestination;
        shifterReg_6_0_bits_decodeResult_maskLogic <= validSource_6_bits_decodeResult_maskLogic;
        shifterReg_6_0_bits_decodeResult_uop <= validSource_6_bits_decodeResult_uop;
        shifterReg_6_0_bits_decodeResult_iota <= validSource_6_bits_decodeResult_iota;
        shifterReg_6_0_bits_decodeResult_mv <= validSource_6_bits_decodeResult_mv;
        shifterReg_6_0_bits_decodeResult_extend <= validSource_6_bits_decodeResult_extend;
        shifterReg_6_0_bits_decodeResult_unOrderWrite <= validSource_6_bits_decodeResult_unOrderWrite;
        shifterReg_6_0_bits_decodeResult_compress <= validSource_6_bits_decodeResult_compress;
        shifterReg_6_0_bits_decodeResult_gather16 <= validSource_6_bits_decodeResult_gather16;
        shifterReg_6_0_bits_decodeResult_gather <= validSource_6_bits_decodeResult_gather;
        shifterReg_6_0_bits_decodeResult_slid <= validSource_6_bits_decodeResult_slid;
        shifterReg_6_0_bits_decodeResult_targetRd <= validSource_6_bits_decodeResult_targetRd;
        shifterReg_6_0_bits_decodeResult_widenReduce <= validSource_6_bits_decodeResult_widenReduce;
        shifterReg_6_0_bits_decodeResult_red <= validSource_6_bits_decodeResult_red;
        shifterReg_6_0_bits_decodeResult_nr <= validSource_6_bits_decodeResult_nr;
        shifterReg_6_0_bits_decodeResult_itype <= validSource_6_bits_decodeResult_itype;
        shifterReg_6_0_bits_decodeResult_unsigned1 <= validSource_6_bits_decodeResult_unsigned1;
        shifterReg_6_0_bits_decodeResult_unsigned0 <= validSource_6_bits_decodeResult_unsigned0;
        shifterReg_6_0_bits_decodeResult_other <= validSource_6_bits_decodeResult_other;
        shifterReg_6_0_bits_decodeResult_multiCycle <= validSource_6_bits_decodeResult_multiCycle;
        shifterReg_6_0_bits_decodeResult_divider <= validSource_6_bits_decodeResult_divider;
        shifterReg_6_0_bits_decodeResult_multiplier <= validSource_6_bits_decodeResult_multiplier;
        shifterReg_6_0_bits_decodeResult_shift <= validSource_6_bits_decodeResult_shift;
        shifterReg_6_0_bits_decodeResult_adder <= validSource_6_bits_decodeResult_adder;
        shifterReg_6_0_bits_decodeResult_logic <= validSource_6_bits_decodeResult_logic;
        shifterReg_6_0_bits_loadStore <= validSource_6_bits_loadStore;
        shifterReg_6_0_bits_issueInst <= validSource_6_bits_issueInst;
        shifterReg_6_0_bits_store <= validSource_6_bits_store;
        shifterReg_6_0_bits_special <= validSource_6_bits_special;
        shifterReg_6_0_bits_lsWholeReg <= validSource_6_bits_lsWholeReg;
        shifterReg_6_0_bits_vs1 <= validSource_6_bits_vs1;
        shifterReg_6_0_bits_vs2 <= validSource_6_bits_vs2;
        shifterReg_6_0_bits_vd <= validSource_6_bits_vd;
        shifterReg_6_0_bits_loadStoreEEW <= validSource_6_bits_loadStoreEEW;
        shifterReg_6_0_bits_mask <= validSource_6_bits_mask;
        shifterReg_6_0_bits_segment <= validSource_6_bits_segment;
        shifterReg_6_0_bits_readFromScalar <= validSource_6_bits_readFromScalar;
        shifterReg_6_0_bits_csrInterface_vl <= validSource_6_bits_csrInterface_vl;
        shifterReg_6_0_bits_csrInterface_vStart <= validSource_6_bits_csrInterface_vStart;
        shifterReg_6_0_bits_csrInterface_vlmul <= validSource_6_bits_csrInterface_vlmul;
        shifterReg_6_0_bits_csrInterface_vSew <= validSource_6_bits_csrInterface_vSew;
        shifterReg_6_0_bits_csrInterface_vxrm <= validSource_6_bits_csrInterface_vxrm;
        shifterReg_6_0_bits_csrInterface_vta <= validSource_6_bits_csrInterface_vta;
        shifterReg_6_0_bits_csrInterface_vma <= validSource_6_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_7 <= laneVec_7_laneRequest_bits_issueInst;
      if (validSource_7_valid ^ releasePipe_pipe_out_7_valid)
        tokenCheck_counter_7 <= tokenCheck_counter_7 + tokenCheck_counterChange_7;
      if (shifterValid_7) begin
        shifterReg_7_0_valid <= validSource_7_valid;
        shifterReg_7_0_bits_instructionIndex <= validSource_7_bits_instructionIndex;
        shifterReg_7_0_bits_decodeResult_orderReduce <= validSource_7_bits_decodeResult_orderReduce;
        shifterReg_7_0_bits_decodeResult_floatMul <= validSource_7_bits_decodeResult_floatMul;
        shifterReg_7_0_bits_decodeResult_fpExecutionType <= validSource_7_bits_decodeResult_fpExecutionType;
        shifterReg_7_0_bits_decodeResult_float <= validSource_7_bits_decodeResult_float;
        shifterReg_7_0_bits_decodeResult_specialSlot <= validSource_7_bits_decodeResult_specialSlot;
        shifterReg_7_0_bits_decodeResult_topUop <= validSource_7_bits_decodeResult_topUop;
        shifterReg_7_0_bits_decodeResult_popCount <= validSource_7_bits_decodeResult_popCount;
        shifterReg_7_0_bits_decodeResult_ffo <= validSource_7_bits_decodeResult_ffo;
        shifterReg_7_0_bits_decodeResult_average <= validSource_7_bits_decodeResult_average;
        shifterReg_7_0_bits_decodeResult_reverse <= validSource_7_bits_decodeResult_reverse;
        shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_7_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_7_0_bits_decodeResult_scheduler <= validSource_7_bits_decodeResult_scheduler;
        shifterReg_7_0_bits_decodeResult_sReadVD <= validSource_7_bits_decodeResult_sReadVD;
        shifterReg_7_0_bits_decodeResult_vtype <= validSource_7_bits_decodeResult_vtype;
        shifterReg_7_0_bits_decodeResult_sWrite <= validSource_7_bits_decodeResult_sWrite;
        shifterReg_7_0_bits_decodeResult_crossRead <= validSource_7_bits_decodeResult_crossRead;
        shifterReg_7_0_bits_decodeResult_crossWrite <= validSource_7_bits_decodeResult_crossWrite;
        shifterReg_7_0_bits_decodeResult_maskUnit <= validSource_7_bits_decodeResult_maskUnit;
        shifterReg_7_0_bits_decodeResult_special <= validSource_7_bits_decodeResult_special;
        shifterReg_7_0_bits_decodeResult_saturate <= validSource_7_bits_decodeResult_saturate;
        shifterReg_7_0_bits_decodeResult_vwmacc <= validSource_7_bits_decodeResult_vwmacc;
        shifterReg_7_0_bits_decodeResult_readOnly <= validSource_7_bits_decodeResult_readOnly;
        shifterReg_7_0_bits_decodeResult_maskSource <= validSource_7_bits_decodeResult_maskSource;
        shifterReg_7_0_bits_decodeResult_maskDestination <= validSource_7_bits_decodeResult_maskDestination;
        shifterReg_7_0_bits_decodeResult_maskLogic <= validSource_7_bits_decodeResult_maskLogic;
        shifterReg_7_0_bits_decodeResult_uop <= validSource_7_bits_decodeResult_uop;
        shifterReg_7_0_bits_decodeResult_iota <= validSource_7_bits_decodeResult_iota;
        shifterReg_7_0_bits_decodeResult_mv <= validSource_7_bits_decodeResult_mv;
        shifterReg_7_0_bits_decodeResult_extend <= validSource_7_bits_decodeResult_extend;
        shifterReg_7_0_bits_decodeResult_unOrderWrite <= validSource_7_bits_decodeResult_unOrderWrite;
        shifterReg_7_0_bits_decodeResult_compress <= validSource_7_bits_decodeResult_compress;
        shifterReg_7_0_bits_decodeResult_gather16 <= validSource_7_bits_decodeResult_gather16;
        shifterReg_7_0_bits_decodeResult_gather <= validSource_7_bits_decodeResult_gather;
        shifterReg_7_0_bits_decodeResult_slid <= validSource_7_bits_decodeResult_slid;
        shifterReg_7_0_bits_decodeResult_targetRd <= validSource_7_bits_decodeResult_targetRd;
        shifterReg_7_0_bits_decodeResult_widenReduce <= validSource_7_bits_decodeResult_widenReduce;
        shifterReg_7_0_bits_decodeResult_red <= validSource_7_bits_decodeResult_red;
        shifterReg_7_0_bits_decodeResult_nr <= validSource_7_bits_decodeResult_nr;
        shifterReg_7_0_bits_decodeResult_itype <= validSource_7_bits_decodeResult_itype;
        shifterReg_7_0_bits_decodeResult_unsigned1 <= validSource_7_bits_decodeResult_unsigned1;
        shifterReg_7_0_bits_decodeResult_unsigned0 <= validSource_7_bits_decodeResult_unsigned0;
        shifterReg_7_0_bits_decodeResult_other <= validSource_7_bits_decodeResult_other;
        shifterReg_7_0_bits_decodeResult_multiCycle <= validSource_7_bits_decodeResult_multiCycle;
        shifterReg_7_0_bits_decodeResult_divider <= validSource_7_bits_decodeResult_divider;
        shifterReg_7_0_bits_decodeResult_multiplier <= validSource_7_bits_decodeResult_multiplier;
        shifterReg_7_0_bits_decodeResult_shift <= validSource_7_bits_decodeResult_shift;
        shifterReg_7_0_bits_decodeResult_adder <= validSource_7_bits_decodeResult_adder;
        shifterReg_7_0_bits_decodeResult_logic <= validSource_7_bits_decodeResult_logic;
        shifterReg_7_0_bits_loadStore <= validSource_7_bits_loadStore;
        shifterReg_7_0_bits_issueInst <= validSource_7_bits_issueInst;
        shifterReg_7_0_bits_store <= validSource_7_bits_store;
        shifterReg_7_0_bits_special <= validSource_7_bits_special;
        shifterReg_7_0_bits_lsWholeReg <= validSource_7_bits_lsWholeReg;
        shifterReg_7_0_bits_vs1 <= validSource_7_bits_vs1;
        shifterReg_7_0_bits_vs2 <= validSource_7_bits_vs2;
        shifterReg_7_0_bits_vd <= validSource_7_bits_vd;
        shifterReg_7_0_bits_loadStoreEEW <= validSource_7_bits_loadStoreEEW;
        shifterReg_7_0_bits_mask <= validSource_7_bits_mask;
        shifterReg_7_0_bits_segment <= validSource_7_bits_segment;
        shifterReg_7_0_bits_readFromScalar <= validSource_7_bits_readFromScalar;
        shifterReg_7_0_bits_csrInterface_vl <= validSource_7_bits_csrInterface_vl;
        shifterReg_7_0_bits_csrInterface_vStart <= validSource_7_bits_csrInterface_vStart;
        shifterReg_7_0_bits_csrInterface_vlmul <= validSource_7_bits_csrInterface_vlmul;
        shifterReg_7_0_bits_csrInterface_vSew <= validSource_7_bits_csrInterface_vSew;
        shifterReg_7_0_bits_csrInterface_vxrm <= validSource_7_bits_csrInterface_vxrm;
        shifterReg_7_0_bits_csrInterface_vta <= validSource_7_bits_csrInterface_vta;
        shifterReg_7_0_bits_csrInterface_vma <= validSource_7_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_8 <= laneVec_8_laneRequest_bits_issueInst;
      if (validSource_8_valid ^ releasePipe_pipe_out_8_valid)
        tokenCheck_counter_8 <= tokenCheck_counter_8 + tokenCheck_counterChange_8;
      if (shifterValid_8) begin
        shifterReg_8_0_valid <= validSource_8_valid;
        shifterReg_8_0_bits_instructionIndex <= validSource_8_bits_instructionIndex;
        shifterReg_8_0_bits_decodeResult_orderReduce <= validSource_8_bits_decodeResult_orderReduce;
        shifterReg_8_0_bits_decodeResult_floatMul <= validSource_8_bits_decodeResult_floatMul;
        shifterReg_8_0_bits_decodeResult_fpExecutionType <= validSource_8_bits_decodeResult_fpExecutionType;
        shifterReg_8_0_bits_decodeResult_float <= validSource_8_bits_decodeResult_float;
        shifterReg_8_0_bits_decodeResult_specialSlot <= validSource_8_bits_decodeResult_specialSlot;
        shifterReg_8_0_bits_decodeResult_topUop <= validSource_8_bits_decodeResult_topUop;
        shifterReg_8_0_bits_decodeResult_popCount <= validSource_8_bits_decodeResult_popCount;
        shifterReg_8_0_bits_decodeResult_ffo <= validSource_8_bits_decodeResult_ffo;
        shifterReg_8_0_bits_decodeResult_average <= validSource_8_bits_decodeResult_average;
        shifterReg_8_0_bits_decodeResult_reverse <= validSource_8_bits_decodeResult_reverse;
        shifterReg_8_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_8_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_8_0_bits_decodeResult_scheduler <= validSource_8_bits_decodeResult_scheduler;
        shifterReg_8_0_bits_decodeResult_sReadVD <= validSource_8_bits_decodeResult_sReadVD;
        shifterReg_8_0_bits_decodeResult_vtype <= validSource_8_bits_decodeResult_vtype;
        shifterReg_8_0_bits_decodeResult_sWrite <= validSource_8_bits_decodeResult_sWrite;
        shifterReg_8_0_bits_decodeResult_crossRead <= validSource_8_bits_decodeResult_crossRead;
        shifterReg_8_0_bits_decodeResult_crossWrite <= validSource_8_bits_decodeResult_crossWrite;
        shifterReg_8_0_bits_decodeResult_maskUnit <= validSource_8_bits_decodeResult_maskUnit;
        shifterReg_8_0_bits_decodeResult_special <= validSource_8_bits_decodeResult_special;
        shifterReg_8_0_bits_decodeResult_saturate <= validSource_8_bits_decodeResult_saturate;
        shifterReg_8_0_bits_decodeResult_vwmacc <= validSource_8_bits_decodeResult_vwmacc;
        shifterReg_8_0_bits_decodeResult_readOnly <= validSource_8_bits_decodeResult_readOnly;
        shifterReg_8_0_bits_decodeResult_maskSource <= validSource_8_bits_decodeResult_maskSource;
        shifterReg_8_0_bits_decodeResult_maskDestination <= validSource_8_bits_decodeResult_maskDestination;
        shifterReg_8_0_bits_decodeResult_maskLogic <= validSource_8_bits_decodeResult_maskLogic;
        shifterReg_8_0_bits_decodeResult_uop <= validSource_8_bits_decodeResult_uop;
        shifterReg_8_0_bits_decodeResult_iota <= validSource_8_bits_decodeResult_iota;
        shifterReg_8_0_bits_decodeResult_mv <= validSource_8_bits_decodeResult_mv;
        shifterReg_8_0_bits_decodeResult_extend <= validSource_8_bits_decodeResult_extend;
        shifterReg_8_0_bits_decodeResult_unOrderWrite <= validSource_8_bits_decodeResult_unOrderWrite;
        shifterReg_8_0_bits_decodeResult_compress <= validSource_8_bits_decodeResult_compress;
        shifterReg_8_0_bits_decodeResult_gather16 <= validSource_8_bits_decodeResult_gather16;
        shifterReg_8_0_bits_decodeResult_gather <= validSource_8_bits_decodeResult_gather;
        shifterReg_8_0_bits_decodeResult_slid <= validSource_8_bits_decodeResult_slid;
        shifterReg_8_0_bits_decodeResult_targetRd <= validSource_8_bits_decodeResult_targetRd;
        shifterReg_8_0_bits_decodeResult_widenReduce <= validSource_8_bits_decodeResult_widenReduce;
        shifterReg_8_0_bits_decodeResult_red <= validSource_8_bits_decodeResult_red;
        shifterReg_8_0_bits_decodeResult_nr <= validSource_8_bits_decodeResult_nr;
        shifterReg_8_0_bits_decodeResult_itype <= validSource_8_bits_decodeResult_itype;
        shifterReg_8_0_bits_decodeResult_unsigned1 <= validSource_8_bits_decodeResult_unsigned1;
        shifterReg_8_0_bits_decodeResult_unsigned0 <= validSource_8_bits_decodeResult_unsigned0;
        shifterReg_8_0_bits_decodeResult_other <= validSource_8_bits_decodeResult_other;
        shifterReg_8_0_bits_decodeResult_multiCycle <= validSource_8_bits_decodeResult_multiCycle;
        shifterReg_8_0_bits_decodeResult_divider <= validSource_8_bits_decodeResult_divider;
        shifterReg_8_0_bits_decodeResult_multiplier <= validSource_8_bits_decodeResult_multiplier;
        shifterReg_8_0_bits_decodeResult_shift <= validSource_8_bits_decodeResult_shift;
        shifterReg_8_0_bits_decodeResult_adder <= validSource_8_bits_decodeResult_adder;
        shifterReg_8_0_bits_decodeResult_logic <= validSource_8_bits_decodeResult_logic;
        shifterReg_8_0_bits_loadStore <= validSource_8_bits_loadStore;
        shifterReg_8_0_bits_issueInst <= validSource_8_bits_issueInst;
        shifterReg_8_0_bits_store <= validSource_8_bits_store;
        shifterReg_8_0_bits_special <= validSource_8_bits_special;
        shifterReg_8_0_bits_lsWholeReg <= validSource_8_bits_lsWholeReg;
        shifterReg_8_0_bits_vs1 <= validSource_8_bits_vs1;
        shifterReg_8_0_bits_vs2 <= validSource_8_bits_vs2;
        shifterReg_8_0_bits_vd <= validSource_8_bits_vd;
        shifterReg_8_0_bits_loadStoreEEW <= validSource_8_bits_loadStoreEEW;
        shifterReg_8_0_bits_mask <= validSource_8_bits_mask;
        shifterReg_8_0_bits_segment <= validSource_8_bits_segment;
        shifterReg_8_0_bits_readFromScalar <= validSource_8_bits_readFromScalar;
        shifterReg_8_0_bits_csrInterface_vl <= validSource_8_bits_csrInterface_vl;
        shifterReg_8_0_bits_csrInterface_vStart <= validSource_8_bits_csrInterface_vStart;
        shifterReg_8_0_bits_csrInterface_vlmul <= validSource_8_bits_csrInterface_vlmul;
        shifterReg_8_0_bits_csrInterface_vSew <= validSource_8_bits_csrInterface_vSew;
        shifterReg_8_0_bits_csrInterface_vxrm <= validSource_8_bits_csrInterface_vxrm;
        shifterReg_8_0_bits_csrInterface_vta <= validSource_8_bits_csrInterface_vta;
        shifterReg_8_0_bits_csrInterface_vma <= validSource_8_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_9 <= laneVec_9_laneRequest_bits_issueInst;
      if (validSource_9_valid ^ releasePipe_pipe_out_9_valid)
        tokenCheck_counter_9 <= tokenCheck_counter_9 + tokenCheck_counterChange_9;
      if (shifterValid_9) begin
        shifterReg_9_0_valid <= validSource_9_valid;
        shifterReg_9_0_bits_instructionIndex <= validSource_9_bits_instructionIndex;
        shifterReg_9_0_bits_decodeResult_orderReduce <= validSource_9_bits_decodeResult_orderReduce;
        shifterReg_9_0_bits_decodeResult_floatMul <= validSource_9_bits_decodeResult_floatMul;
        shifterReg_9_0_bits_decodeResult_fpExecutionType <= validSource_9_bits_decodeResult_fpExecutionType;
        shifterReg_9_0_bits_decodeResult_float <= validSource_9_bits_decodeResult_float;
        shifterReg_9_0_bits_decodeResult_specialSlot <= validSource_9_bits_decodeResult_specialSlot;
        shifterReg_9_0_bits_decodeResult_topUop <= validSource_9_bits_decodeResult_topUop;
        shifterReg_9_0_bits_decodeResult_popCount <= validSource_9_bits_decodeResult_popCount;
        shifterReg_9_0_bits_decodeResult_ffo <= validSource_9_bits_decodeResult_ffo;
        shifterReg_9_0_bits_decodeResult_average <= validSource_9_bits_decodeResult_average;
        shifterReg_9_0_bits_decodeResult_reverse <= validSource_9_bits_decodeResult_reverse;
        shifterReg_9_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_9_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_9_0_bits_decodeResult_scheduler <= validSource_9_bits_decodeResult_scheduler;
        shifterReg_9_0_bits_decodeResult_sReadVD <= validSource_9_bits_decodeResult_sReadVD;
        shifterReg_9_0_bits_decodeResult_vtype <= validSource_9_bits_decodeResult_vtype;
        shifterReg_9_0_bits_decodeResult_sWrite <= validSource_9_bits_decodeResult_sWrite;
        shifterReg_9_0_bits_decodeResult_crossRead <= validSource_9_bits_decodeResult_crossRead;
        shifterReg_9_0_bits_decodeResult_crossWrite <= validSource_9_bits_decodeResult_crossWrite;
        shifterReg_9_0_bits_decodeResult_maskUnit <= validSource_9_bits_decodeResult_maskUnit;
        shifterReg_9_0_bits_decodeResult_special <= validSource_9_bits_decodeResult_special;
        shifterReg_9_0_bits_decodeResult_saturate <= validSource_9_bits_decodeResult_saturate;
        shifterReg_9_0_bits_decodeResult_vwmacc <= validSource_9_bits_decodeResult_vwmacc;
        shifterReg_9_0_bits_decodeResult_readOnly <= validSource_9_bits_decodeResult_readOnly;
        shifterReg_9_0_bits_decodeResult_maskSource <= validSource_9_bits_decodeResult_maskSource;
        shifterReg_9_0_bits_decodeResult_maskDestination <= validSource_9_bits_decodeResult_maskDestination;
        shifterReg_9_0_bits_decodeResult_maskLogic <= validSource_9_bits_decodeResult_maskLogic;
        shifterReg_9_0_bits_decodeResult_uop <= validSource_9_bits_decodeResult_uop;
        shifterReg_9_0_bits_decodeResult_iota <= validSource_9_bits_decodeResult_iota;
        shifterReg_9_0_bits_decodeResult_mv <= validSource_9_bits_decodeResult_mv;
        shifterReg_9_0_bits_decodeResult_extend <= validSource_9_bits_decodeResult_extend;
        shifterReg_9_0_bits_decodeResult_unOrderWrite <= validSource_9_bits_decodeResult_unOrderWrite;
        shifterReg_9_0_bits_decodeResult_compress <= validSource_9_bits_decodeResult_compress;
        shifterReg_9_0_bits_decodeResult_gather16 <= validSource_9_bits_decodeResult_gather16;
        shifterReg_9_0_bits_decodeResult_gather <= validSource_9_bits_decodeResult_gather;
        shifterReg_9_0_bits_decodeResult_slid <= validSource_9_bits_decodeResult_slid;
        shifterReg_9_0_bits_decodeResult_targetRd <= validSource_9_bits_decodeResult_targetRd;
        shifterReg_9_0_bits_decodeResult_widenReduce <= validSource_9_bits_decodeResult_widenReduce;
        shifterReg_9_0_bits_decodeResult_red <= validSource_9_bits_decodeResult_red;
        shifterReg_9_0_bits_decodeResult_nr <= validSource_9_bits_decodeResult_nr;
        shifterReg_9_0_bits_decodeResult_itype <= validSource_9_bits_decodeResult_itype;
        shifterReg_9_0_bits_decodeResult_unsigned1 <= validSource_9_bits_decodeResult_unsigned1;
        shifterReg_9_0_bits_decodeResult_unsigned0 <= validSource_9_bits_decodeResult_unsigned0;
        shifterReg_9_0_bits_decodeResult_other <= validSource_9_bits_decodeResult_other;
        shifterReg_9_0_bits_decodeResult_multiCycle <= validSource_9_bits_decodeResult_multiCycle;
        shifterReg_9_0_bits_decodeResult_divider <= validSource_9_bits_decodeResult_divider;
        shifterReg_9_0_bits_decodeResult_multiplier <= validSource_9_bits_decodeResult_multiplier;
        shifterReg_9_0_bits_decodeResult_shift <= validSource_9_bits_decodeResult_shift;
        shifterReg_9_0_bits_decodeResult_adder <= validSource_9_bits_decodeResult_adder;
        shifterReg_9_0_bits_decodeResult_logic <= validSource_9_bits_decodeResult_logic;
        shifterReg_9_0_bits_loadStore <= validSource_9_bits_loadStore;
        shifterReg_9_0_bits_issueInst <= validSource_9_bits_issueInst;
        shifterReg_9_0_bits_store <= validSource_9_bits_store;
        shifterReg_9_0_bits_special <= validSource_9_bits_special;
        shifterReg_9_0_bits_lsWholeReg <= validSource_9_bits_lsWholeReg;
        shifterReg_9_0_bits_vs1 <= validSource_9_bits_vs1;
        shifterReg_9_0_bits_vs2 <= validSource_9_bits_vs2;
        shifterReg_9_0_bits_vd <= validSource_9_bits_vd;
        shifterReg_9_0_bits_loadStoreEEW <= validSource_9_bits_loadStoreEEW;
        shifterReg_9_0_bits_mask <= validSource_9_bits_mask;
        shifterReg_9_0_bits_segment <= validSource_9_bits_segment;
        shifterReg_9_0_bits_readFromScalar <= validSource_9_bits_readFromScalar;
        shifterReg_9_0_bits_csrInterface_vl <= validSource_9_bits_csrInterface_vl;
        shifterReg_9_0_bits_csrInterface_vStart <= validSource_9_bits_csrInterface_vStart;
        shifterReg_9_0_bits_csrInterface_vlmul <= validSource_9_bits_csrInterface_vlmul;
        shifterReg_9_0_bits_csrInterface_vSew <= validSource_9_bits_csrInterface_vSew;
        shifterReg_9_0_bits_csrInterface_vxrm <= validSource_9_bits_csrInterface_vxrm;
        shifterReg_9_0_bits_csrInterface_vta <= validSource_9_bits_csrInterface_vta;
        shifterReg_9_0_bits_csrInterface_vma <= validSource_9_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_10 <= laneVec_10_laneRequest_bits_issueInst;
      if (validSource_10_valid ^ releasePipe_pipe_out_10_valid)
        tokenCheck_counter_10 <= tokenCheck_counter_10 + tokenCheck_counterChange_10;
      if (shifterValid_10) begin
        shifterReg_10_0_valid <= validSource_10_valid;
        shifterReg_10_0_bits_instructionIndex <= validSource_10_bits_instructionIndex;
        shifterReg_10_0_bits_decodeResult_orderReduce <= validSource_10_bits_decodeResult_orderReduce;
        shifterReg_10_0_bits_decodeResult_floatMul <= validSource_10_bits_decodeResult_floatMul;
        shifterReg_10_0_bits_decodeResult_fpExecutionType <= validSource_10_bits_decodeResult_fpExecutionType;
        shifterReg_10_0_bits_decodeResult_float <= validSource_10_bits_decodeResult_float;
        shifterReg_10_0_bits_decodeResult_specialSlot <= validSource_10_bits_decodeResult_specialSlot;
        shifterReg_10_0_bits_decodeResult_topUop <= validSource_10_bits_decodeResult_topUop;
        shifterReg_10_0_bits_decodeResult_popCount <= validSource_10_bits_decodeResult_popCount;
        shifterReg_10_0_bits_decodeResult_ffo <= validSource_10_bits_decodeResult_ffo;
        shifterReg_10_0_bits_decodeResult_average <= validSource_10_bits_decodeResult_average;
        shifterReg_10_0_bits_decodeResult_reverse <= validSource_10_bits_decodeResult_reverse;
        shifterReg_10_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_10_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_10_0_bits_decodeResult_scheduler <= validSource_10_bits_decodeResult_scheduler;
        shifterReg_10_0_bits_decodeResult_sReadVD <= validSource_10_bits_decodeResult_sReadVD;
        shifterReg_10_0_bits_decodeResult_vtype <= validSource_10_bits_decodeResult_vtype;
        shifterReg_10_0_bits_decodeResult_sWrite <= validSource_10_bits_decodeResult_sWrite;
        shifterReg_10_0_bits_decodeResult_crossRead <= validSource_10_bits_decodeResult_crossRead;
        shifterReg_10_0_bits_decodeResult_crossWrite <= validSource_10_bits_decodeResult_crossWrite;
        shifterReg_10_0_bits_decodeResult_maskUnit <= validSource_10_bits_decodeResult_maskUnit;
        shifterReg_10_0_bits_decodeResult_special <= validSource_10_bits_decodeResult_special;
        shifterReg_10_0_bits_decodeResult_saturate <= validSource_10_bits_decodeResult_saturate;
        shifterReg_10_0_bits_decodeResult_vwmacc <= validSource_10_bits_decodeResult_vwmacc;
        shifterReg_10_0_bits_decodeResult_readOnly <= validSource_10_bits_decodeResult_readOnly;
        shifterReg_10_0_bits_decodeResult_maskSource <= validSource_10_bits_decodeResult_maskSource;
        shifterReg_10_0_bits_decodeResult_maskDestination <= validSource_10_bits_decodeResult_maskDestination;
        shifterReg_10_0_bits_decodeResult_maskLogic <= validSource_10_bits_decodeResult_maskLogic;
        shifterReg_10_0_bits_decodeResult_uop <= validSource_10_bits_decodeResult_uop;
        shifterReg_10_0_bits_decodeResult_iota <= validSource_10_bits_decodeResult_iota;
        shifterReg_10_0_bits_decodeResult_mv <= validSource_10_bits_decodeResult_mv;
        shifterReg_10_0_bits_decodeResult_extend <= validSource_10_bits_decodeResult_extend;
        shifterReg_10_0_bits_decodeResult_unOrderWrite <= validSource_10_bits_decodeResult_unOrderWrite;
        shifterReg_10_0_bits_decodeResult_compress <= validSource_10_bits_decodeResult_compress;
        shifterReg_10_0_bits_decodeResult_gather16 <= validSource_10_bits_decodeResult_gather16;
        shifterReg_10_0_bits_decodeResult_gather <= validSource_10_bits_decodeResult_gather;
        shifterReg_10_0_bits_decodeResult_slid <= validSource_10_bits_decodeResult_slid;
        shifterReg_10_0_bits_decodeResult_targetRd <= validSource_10_bits_decodeResult_targetRd;
        shifterReg_10_0_bits_decodeResult_widenReduce <= validSource_10_bits_decodeResult_widenReduce;
        shifterReg_10_0_bits_decodeResult_red <= validSource_10_bits_decodeResult_red;
        shifterReg_10_0_bits_decodeResult_nr <= validSource_10_bits_decodeResult_nr;
        shifterReg_10_0_bits_decodeResult_itype <= validSource_10_bits_decodeResult_itype;
        shifterReg_10_0_bits_decodeResult_unsigned1 <= validSource_10_bits_decodeResult_unsigned1;
        shifterReg_10_0_bits_decodeResult_unsigned0 <= validSource_10_bits_decodeResult_unsigned0;
        shifterReg_10_0_bits_decodeResult_other <= validSource_10_bits_decodeResult_other;
        shifterReg_10_0_bits_decodeResult_multiCycle <= validSource_10_bits_decodeResult_multiCycle;
        shifterReg_10_0_bits_decodeResult_divider <= validSource_10_bits_decodeResult_divider;
        shifterReg_10_0_bits_decodeResult_multiplier <= validSource_10_bits_decodeResult_multiplier;
        shifterReg_10_0_bits_decodeResult_shift <= validSource_10_bits_decodeResult_shift;
        shifterReg_10_0_bits_decodeResult_adder <= validSource_10_bits_decodeResult_adder;
        shifterReg_10_0_bits_decodeResult_logic <= validSource_10_bits_decodeResult_logic;
        shifterReg_10_0_bits_loadStore <= validSource_10_bits_loadStore;
        shifterReg_10_0_bits_issueInst <= validSource_10_bits_issueInst;
        shifterReg_10_0_bits_store <= validSource_10_bits_store;
        shifterReg_10_0_bits_special <= validSource_10_bits_special;
        shifterReg_10_0_bits_lsWholeReg <= validSource_10_bits_lsWholeReg;
        shifterReg_10_0_bits_vs1 <= validSource_10_bits_vs1;
        shifterReg_10_0_bits_vs2 <= validSource_10_bits_vs2;
        shifterReg_10_0_bits_vd <= validSource_10_bits_vd;
        shifterReg_10_0_bits_loadStoreEEW <= validSource_10_bits_loadStoreEEW;
        shifterReg_10_0_bits_mask <= validSource_10_bits_mask;
        shifterReg_10_0_bits_segment <= validSource_10_bits_segment;
        shifterReg_10_0_bits_readFromScalar <= validSource_10_bits_readFromScalar;
        shifterReg_10_0_bits_csrInterface_vl <= validSource_10_bits_csrInterface_vl;
        shifterReg_10_0_bits_csrInterface_vStart <= validSource_10_bits_csrInterface_vStart;
        shifterReg_10_0_bits_csrInterface_vlmul <= validSource_10_bits_csrInterface_vlmul;
        shifterReg_10_0_bits_csrInterface_vSew <= validSource_10_bits_csrInterface_vSew;
        shifterReg_10_0_bits_csrInterface_vxrm <= validSource_10_bits_csrInterface_vxrm;
        shifterReg_10_0_bits_csrInterface_vta <= validSource_10_bits_csrInterface_vta;
        shifterReg_10_0_bits_csrInterface_vma <= validSource_10_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_11 <= laneVec_11_laneRequest_bits_issueInst;
      if (validSource_11_valid ^ releasePipe_pipe_out_11_valid)
        tokenCheck_counter_11 <= tokenCheck_counter_11 + tokenCheck_counterChange_11;
      if (shifterValid_11) begin
        shifterReg_11_0_valid <= validSource_11_valid;
        shifterReg_11_0_bits_instructionIndex <= validSource_11_bits_instructionIndex;
        shifterReg_11_0_bits_decodeResult_orderReduce <= validSource_11_bits_decodeResult_orderReduce;
        shifterReg_11_0_bits_decodeResult_floatMul <= validSource_11_bits_decodeResult_floatMul;
        shifterReg_11_0_bits_decodeResult_fpExecutionType <= validSource_11_bits_decodeResult_fpExecutionType;
        shifterReg_11_0_bits_decodeResult_float <= validSource_11_bits_decodeResult_float;
        shifterReg_11_0_bits_decodeResult_specialSlot <= validSource_11_bits_decodeResult_specialSlot;
        shifterReg_11_0_bits_decodeResult_topUop <= validSource_11_bits_decodeResult_topUop;
        shifterReg_11_0_bits_decodeResult_popCount <= validSource_11_bits_decodeResult_popCount;
        shifterReg_11_0_bits_decodeResult_ffo <= validSource_11_bits_decodeResult_ffo;
        shifterReg_11_0_bits_decodeResult_average <= validSource_11_bits_decodeResult_average;
        shifterReg_11_0_bits_decodeResult_reverse <= validSource_11_bits_decodeResult_reverse;
        shifterReg_11_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_11_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_11_0_bits_decodeResult_scheduler <= validSource_11_bits_decodeResult_scheduler;
        shifterReg_11_0_bits_decodeResult_sReadVD <= validSource_11_bits_decodeResult_sReadVD;
        shifterReg_11_0_bits_decodeResult_vtype <= validSource_11_bits_decodeResult_vtype;
        shifterReg_11_0_bits_decodeResult_sWrite <= validSource_11_bits_decodeResult_sWrite;
        shifterReg_11_0_bits_decodeResult_crossRead <= validSource_11_bits_decodeResult_crossRead;
        shifterReg_11_0_bits_decodeResult_crossWrite <= validSource_11_bits_decodeResult_crossWrite;
        shifterReg_11_0_bits_decodeResult_maskUnit <= validSource_11_bits_decodeResult_maskUnit;
        shifterReg_11_0_bits_decodeResult_special <= validSource_11_bits_decodeResult_special;
        shifterReg_11_0_bits_decodeResult_saturate <= validSource_11_bits_decodeResult_saturate;
        shifterReg_11_0_bits_decodeResult_vwmacc <= validSource_11_bits_decodeResult_vwmacc;
        shifterReg_11_0_bits_decodeResult_readOnly <= validSource_11_bits_decodeResult_readOnly;
        shifterReg_11_0_bits_decodeResult_maskSource <= validSource_11_bits_decodeResult_maskSource;
        shifterReg_11_0_bits_decodeResult_maskDestination <= validSource_11_bits_decodeResult_maskDestination;
        shifterReg_11_0_bits_decodeResult_maskLogic <= validSource_11_bits_decodeResult_maskLogic;
        shifterReg_11_0_bits_decodeResult_uop <= validSource_11_bits_decodeResult_uop;
        shifterReg_11_0_bits_decodeResult_iota <= validSource_11_bits_decodeResult_iota;
        shifterReg_11_0_bits_decodeResult_mv <= validSource_11_bits_decodeResult_mv;
        shifterReg_11_0_bits_decodeResult_extend <= validSource_11_bits_decodeResult_extend;
        shifterReg_11_0_bits_decodeResult_unOrderWrite <= validSource_11_bits_decodeResult_unOrderWrite;
        shifterReg_11_0_bits_decodeResult_compress <= validSource_11_bits_decodeResult_compress;
        shifterReg_11_0_bits_decodeResult_gather16 <= validSource_11_bits_decodeResult_gather16;
        shifterReg_11_0_bits_decodeResult_gather <= validSource_11_bits_decodeResult_gather;
        shifterReg_11_0_bits_decodeResult_slid <= validSource_11_bits_decodeResult_slid;
        shifterReg_11_0_bits_decodeResult_targetRd <= validSource_11_bits_decodeResult_targetRd;
        shifterReg_11_0_bits_decodeResult_widenReduce <= validSource_11_bits_decodeResult_widenReduce;
        shifterReg_11_0_bits_decodeResult_red <= validSource_11_bits_decodeResult_red;
        shifterReg_11_0_bits_decodeResult_nr <= validSource_11_bits_decodeResult_nr;
        shifterReg_11_0_bits_decodeResult_itype <= validSource_11_bits_decodeResult_itype;
        shifterReg_11_0_bits_decodeResult_unsigned1 <= validSource_11_bits_decodeResult_unsigned1;
        shifterReg_11_0_bits_decodeResult_unsigned0 <= validSource_11_bits_decodeResult_unsigned0;
        shifterReg_11_0_bits_decodeResult_other <= validSource_11_bits_decodeResult_other;
        shifterReg_11_0_bits_decodeResult_multiCycle <= validSource_11_bits_decodeResult_multiCycle;
        shifterReg_11_0_bits_decodeResult_divider <= validSource_11_bits_decodeResult_divider;
        shifterReg_11_0_bits_decodeResult_multiplier <= validSource_11_bits_decodeResult_multiplier;
        shifterReg_11_0_bits_decodeResult_shift <= validSource_11_bits_decodeResult_shift;
        shifterReg_11_0_bits_decodeResult_adder <= validSource_11_bits_decodeResult_adder;
        shifterReg_11_0_bits_decodeResult_logic <= validSource_11_bits_decodeResult_logic;
        shifterReg_11_0_bits_loadStore <= validSource_11_bits_loadStore;
        shifterReg_11_0_bits_issueInst <= validSource_11_bits_issueInst;
        shifterReg_11_0_bits_store <= validSource_11_bits_store;
        shifterReg_11_0_bits_special <= validSource_11_bits_special;
        shifterReg_11_0_bits_lsWholeReg <= validSource_11_bits_lsWholeReg;
        shifterReg_11_0_bits_vs1 <= validSource_11_bits_vs1;
        shifterReg_11_0_bits_vs2 <= validSource_11_bits_vs2;
        shifterReg_11_0_bits_vd <= validSource_11_bits_vd;
        shifterReg_11_0_bits_loadStoreEEW <= validSource_11_bits_loadStoreEEW;
        shifterReg_11_0_bits_mask <= validSource_11_bits_mask;
        shifterReg_11_0_bits_segment <= validSource_11_bits_segment;
        shifterReg_11_0_bits_readFromScalar <= validSource_11_bits_readFromScalar;
        shifterReg_11_0_bits_csrInterface_vl <= validSource_11_bits_csrInterface_vl;
        shifterReg_11_0_bits_csrInterface_vStart <= validSource_11_bits_csrInterface_vStart;
        shifterReg_11_0_bits_csrInterface_vlmul <= validSource_11_bits_csrInterface_vlmul;
        shifterReg_11_0_bits_csrInterface_vSew <= validSource_11_bits_csrInterface_vSew;
        shifterReg_11_0_bits_csrInterface_vxrm <= validSource_11_bits_csrInterface_vxrm;
        shifterReg_11_0_bits_csrInterface_vta <= validSource_11_bits_csrInterface_vta;
        shifterReg_11_0_bits_csrInterface_vma <= validSource_11_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_12 <= laneVec_12_laneRequest_bits_issueInst;
      if (validSource_12_valid ^ releasePipe_pipe_out_12_valid)
        tokenCheck_counter_12 <= tokenCheck_counter_12 + tokenCheck_counterChange_12;
      if (shifterValid_12) begin
        shifterReg_12_0_valid <= validSource_12_valid;
        shifterReg_12_0_bits_instructionIndex <= validSource_12_bits_instructionIndex;
        shifterReg_12_0_bits_decodeResult_orderReduce <= validSource_12_bits_decodeResult_orderReduce;
        shifterReg_12_0_bits_decodeResult_floatMul <= validSource_12_bits_decodeResult_floatMul;
        shifterReg_12_0_bits_decodeResult_fpExecutionType <= validSource_12_bits_decodeResult_fpExecutionType;
        shifterReg_12_0_bits_decodeResult_float <= validSource_12_bits_decodeResult_float;
        shifterReg_12_0_bits_decodeResult_specialSlot <= validSource_12_bits_decodeResult_specialSlot;
        shifterReg_12_0_bits_decodeResult_topUop <= validSource_12_bits_decodeResult_topUop;
        shifterReg_12_0_bits_decodeResult_popCount <= validSource_12_bits_decodeResult_popCount;
        shifterReg_12_0_bits_decodeResult_ffo <= validSource_12_bits_decodeResult_ffo;
        shifterReg_12_0_bits_decodeResult_average <= validSource_12_bits_decodeResult_average;
        shifterReg_12_0_bits_decodeResult_reverse <= validSource_12_bits_decodeResult_reverse;
        shifterReg_12_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_12_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_12_0_bits_decodeResult_scheduler <= validSource_12_bits_decodeResult_scheduler;
        shifterReg_12_0_bits_decodeResult_sReadVD <= validSource_12_bits_decodeResult_sReadVD;
        shifterReg_12_0_bits_decodeResult_vtype <= validSource_12_bits_decodeResult_vtype;
        shifterReg_12_0_bits_decodeResult_sWrite <= validSource_12_bits_decodeResult_sWrite;
        shifterReg_12_0_bits_decodeResult_crossRead <= validSource_12_bits_decodeResult_crossRead;
        shifterReg_12_0_bits_decodeResult_crossWrite <= validSource_12_bits_decodeResult_crossWrite;
        shifterReg_12_0_bits_decodeResult_maskUnit <= validSource_12_bits_decodeResult_maskUnit;
        shifterReg_12_0_bits_decodeResult_special <= validSource_12_bits_decodeResult_special;
        shifterReg_12_0_bits_decodeResult_saturate <= validSource_12_bits_decodeResult_saturate;
        shifterReg_12_0_bits_decodeResult_vwmacc <= validSource_12_bits_decodeResult_vwmacc;
        shifterReg_12_0_bits_decodeResult_readOnly <= validSource_12_bits_decodeResult_readOnly;
        shifterReg_12_0_bits_decodeResult_maskSource <= validSource_12_bits_decodeResult_maskSource;
        shifterReg_12_0_bits_decodeResult_maskDestination <= validSource_12_bits_decodeResult_maskDestination;
        shifterReg_12_0_bits_decodeResult_maskLogic <= validSource_12_bits_decodeResult_maskLogic;
        shifterReg_12_0_bits_decodeResult_uop <= validSource_12_bits_decodeResult_uop;
        shifterReg_12_0_bits_decodeResult_iota <= validSource_12_bits_decodeResult_iota;
        shifterReg_12_0_bits_decodeResult_mv <= validSource_12_bits_decodeResult_mv;
        shifterReg_12_0_bits_decodeResult_extend <= validSource_12_bits_decodeResult_extend;
        shifterReg_12_0_bits_decodeResult_unOrderWrite <= validSource_12_bits_decodeResult_unOrderWrite;
        shifterReg_12_0_bits_decodeResult_compress <= validSource_12_bits_decodeResult_compress;
        shifterReg_12_0_bits_decodeResult_gather16 <= validSource_12_bits_decodeResult_gather16;
        shifterReg_12_0_bits_decodeResult_gather <= validSource_12_bits_decodeResult_gather;
        shifterReg_12_0_bits_decodeResult_slid <= validSource_12_bits_decodeResult_slid;
        shifterReg_12_0_bits_decodeResult_targetRd <= validSource_12_bits_decodeResult_targetRd;
        shifterReg_12_0_bits_decodeResult_widenReduce <= validSource_12_bits_decodeResult_widenReduce;
        shifterReg_12_0_bits_decodeResult_red <= validSource_12_bits_decodeResult_red;
        shifterReg_12_0_bits_decodeResult_nr <= validSource_12_bits_decodeResult_nr;
        shifterReg_12_0_bits_decodeResult_itype <= validSource_12_bits_decodeResult_itype;
        shifterReg_12_0_bits_decodeResult_unsigned1 <= validSource_12_bits_decodeResult_unsigned1;
        shifterReg_12_0_bits_decodeResult_unsigned0 <= validSource_12_bits_decodeResult_unsigned0;
        shifterReg_12_0_bits_decodeResult_other <= validSource_12_bits_decodeResult_other;
        shifterReg_12_0_bits_decodeResult_multiCycle <= validSource_12_bits_decodeResult_multiCycle;
        shifterReg_12_0_bits_decodeResult_divider <= validSource_12_bits_decodeResult_divider;
        shifterReg_12_0_bits_decodeResult_multiplier <= validSource_12_bits_decodeResult_multiplier;
        shifterReg_12_0_bits_decodeResult_shift <= validSource_12_bits_decodeResult_shift;
        shifterReg_12_0_bits_decodeResult_adder <= validSource_12_bits_decodeResult_adder;
        shifterReg_12_0_bits_decodeResult_logic <= validSource_12_bits_decodeResult_logic;
        shifterReg_12_0_bits_loadStore <= validSource_12_bits_loadStore;
        shifterReg_12_0_bits_issueInst <= validSource_12_bits_issueInst;
        shifterReg_12_0_bits_store <= validSource_12_bits_store;
        shifterReg_12_0_bits_special <= validSource_12_bits_special;
        shifterReg_12_0_bits_lsWholeReg <= validSource_12_bits_lsWholeReg;
        shifterReg_12_0_bits_vs1 <= validSource_12_bits_vs1;
        shifterReg_12_0_bits_vs2 <= validSource_12_bits_vs2;
        shifterReg_12_0_bits_vd <= validSource_12_bits_vd;
        shifterReg_12_0_bits_loadStoreEEW <= validSource_12_bits_loadStoreEEW;
        shifterReg_12_0_bits_mask <= validSource_12_bits_mask;
        shifterReg_12_0_bits_segment <= validSource_12_bits_segment;
        shifterReg_12_0_bits_readFromScalar <= validSource_12_bits_readFromScalar;
        shifterReg_12_0_bits_csrInterface_vl <= validSource_12_bits_csrInterface_vl;
        shifterReg_12_0_bits_csrInterface_vStart <= validSource_12_bits_csrInterface_vStart;
        shifterReg_12_0_bits_csrInterface_vlmul <= validSource_12_bits_csrInterface_vlmul;
        shifterReg_12_0_bits_csrInterface_vSew <= validSource_12_bits_csrInterface_vSew;
        shifterReg_12_0_bits_csrInterface_vxrm <= validSource_12_bits_csrInterface_vxrm;
        shifterReg_12_0_bits_csrInterface_vta <= validSource_12_bits_csrInterface_vta;
        shifterReg_12_0_bits_csrInterface_vma <= validSource_12_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_13 <= laneVec_13_laneRequest_bits_issueInst;
      if (validSource_13_valid ^ releasePipe_pipe_out_13_valid)
        tokenCheck_counter_13 <= tokenCheck_counter_13 + tokenCheck_counterChange_13;
      if (shifterValid_13) begin
        shifterReg_13_0_valid <= validSource_13_valid;
        shifterReg_13_0_bits_instructionIndex <= validSource_13_bits_instructionIndex;
        shifterReg_13_0_bits_decodeResult_orderReduce <= validSource_13_bits_decodeResult_orderReduce;
        shifterReg_13_0_bits_decodeResult_floatMul <= validSource_13_bits_decodeResult_floatMul;
        shifterReg_13_0_bits_decodeResult_fpExecutionType <= validSource_13_bits_decodeResult_fpExecutionType;
        shifterReg_13_0_bits_decodeResult_float <= validSource_13_bits_decodeResult_float;
        shifterReg_13_0_bits_decodeResult_specialSlot <= validSource_13_bits_decodeResult_specialSlot;
        shifterReg_13_0_bits_decodeResult_topUop <= validSource_13_bits_decodeResult_topUop;
        shifterReg_13_0_bits_decodeResult_popCount <= validSource_13_bits_decodeResult_popCount;
        shifterReg_13_0_bits_decodeResult_ffo <= validSource_13_bits_decodeResult_ffo;
        shifterReg_13_0_bits_decodeResult_average <= validSource_13_bits_decodeResult_average;
        shifterReg_13_0_bits_decodeResult_reverse <= validSource_13_bits_decodeResult_reverse;
        shifterReg_13_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_13_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_13_0_bits_decodeResult_scheduler <= validSource_13_bits_decodeResult_scheduler;
        shifterReg_13_0_bits_decodeResult_sReadVD <= validSource_13_bits_decodeResult_sReadVD;
        shifterReg_13_0_bits_decodeResult_vtype <= validSource_13_bits_decodeResult_vtype;
        shifterReg_13_0_bits_decodeResult_sWrite <= validSource_13_bits_decodeResult_sWrite;
        shifterReg_13_0_bits_decodeResult_crossRead <= validSource_13_bits_decodeResult_crossRead;
        shifterReg_13_0_bits_decodeResult_crossWrite <= validSource_13_bits_decodeResult_crossWrite;
        shifterReg_13_0_bits_decodeResult_maskUnit <= validSource_13_bits_decodeResult_maskUnit;
        shifterReg_13_0_bits_decodeResult_special <= validSource_13_bits_decodeResult_special;
        shifterReg_13_0_bits_decodeResult_saturate <= validSource_13_bits_decodeResult_saturate;
        shifterReg_13_0_bits_decodeResult_vwmacc <= validSource_13_bits_decodeResult_vwmacc;
        shifterReg_13_0_bits_decodeResult_readOnly <= validSource_13_bits_decodeResult_readOnly;
        shifterReg_13_0_bits_decodeResult_maskSource <= validSource_13_bits_decodeResult_maskSource;
        shifterReg_13_0_bits_decodeResult_maskDestination <= validSource_13_bits_decodeResult_maskDestination;
        shifterReg_13_0_bits_decodeResult_maskLogic <= validSource_13_bits_decodeResult_maskLogic;
        shifterReg_13_0_bits_decodeResult_uop <= validSource_13_bits_decodeResult_uop;
        shifterReg_13_0_bits_decodeResult_iota <= validSource_13_bits_decodeResult_iota;
        shifterReg_13_0_bits_decodeResult_mv <= validSource_13_bits_decodeResult_mv;
        shifterReg_13_0_bits_decodeResult_extend <= validSource_13_bits_decodeResult_extend;
        shifterReg_13_0_bits_decodeResult_unOrderWrite <= validSource_13_bits_decodeResult_unOrderWrite;
        shifterReg_13_0_bits_decodeResult_compress <= validSource_13_bits_decodeResult_compress;
        shifterReg_13_0_bits_decodeResult_gather16 <= validSource_13_bits_decodeResult_gather16;
        shifterReg_13_0_bits_decodeResult_gather <= validSource_13_bits_decodeResult_gather;
        shifterReg_13_0_bits_decodeResult_slid <= validSource_13_bits_decodeResult_slid;
        shifterReg_13_0_bits_decodeResult_targetRd <= validSource_13_bits_decodeResult_targetRd;
        shifterReg_13_0_bits_decodeResult_widenReduce <= validSource_13_bits_decodeResult_widenReduce;
        shifterReg_13_0_bits_decodeResult_red <= validSource_13_bits_decodeResult_red;
        shifterReg_13_0_bits_decodeResult_nr <= validSource_13_bits_decodeResult_nr;
        shifterReg_13_0_bits_decodeResult_itype <= validSource_13_bits_decodeResult_itype;
        shifterReg_13_0_bits_decodeResult_unsigned1 <= validSource_13_bits_decodeResult_unsigned1;
        shifterReg_13_0_bits_decodeResult_unsigned0 <= validSource_13_bits_decodeResult_unsigned0;
        shifterReg_13_0_bits_decodeResult_other <= validSource_13_bits_decodeResult_other;
        shifterReg_13_0_bits_decodeResult_multiCycle <= validSource_13_bits_decodeResult_multiCycle;
        shifterReg_13_0_bits_decodeResult_divider <= validSource_13_bits_decodeResult_divider;
        shifterReg_13_0_bits_decodeResult_multiplier <= validSource_13_bits_decodeResult_multiplier;
        shifterReg_13_0_bits_decodeResult_shift <= validSource_13_bits_decodeResult_shift;
        shifterReg_13_0_bits_decodeResult_adder <= validSource_13_bits_decodeResult_adder;
        shifterReg_13_0_bits_decodeResult_logic <= validSource_13_bits_decodeResult_logic;
        shifterReg_13_0_bits_loadStore <= validSource_13_bits_loadStore;
        shifterReg_13_0_bits_issueInst <= validSource_13_bits_issueInst;
        shifterReg_13_0_bits_store <= validSource_13_bits_store;
        shifterReg_13_0_bits_special <= validSource_13_bits_special;
        shifterReg_13_0_bits_lsWholeReg <= validSource_13_bits_lsWholeReg;
        shifterReg_13_0_bits_vs1 <= validSource_13_bits_vs1;
        shifterReg_13_0_bits_vs2 <= validSource_13_bits_vs2;
        shifterReg_13_0_bits_vd <= validSource_13_bits_vd;
        shifterReg_13_0_bits_loadStoreEEW <= validSource_13_bits_loadStoreEEW;
        shifterReg_13_0_bits_mask <= validSource_13_bits_mask;
        shifterReg_13_0_bits_segment <= validSource_13_bits_segment;
        shifterReg_13_0_bits_readFromScalar <= validSource_13_bits_readFromScalar;
        shifterReg_13_0_bits_csrInterface_vl <= validSource_13_bits_csrInterface_vl;
        shifterReg_13_0_bits_csrInterface_vStart <= validSource_13_bits_csrInterface_vStart;
        shifterReg_13_0_bits_csrInterface_vlmul <= validSource_13_bits_csrInterface_vlmul;
        shifterReg_13_0_bits_csrInterface_vSew <= validSource_13_bits_csrInterface_vSew;
        shifterReg_13_0_bits_csrInterface_vxrm <= validSource_13_bits_csrInterface_vxrm;
        shifterReg_13_0_bits_csrInterface_vta <= validSource_13_bits_csrInterface_vta;
        shifterReg_13_0_bits_csrInterface_vma <= validSource_13_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_14 <= laneVec_14_laneRequest_bits_issueInst;
      if (validSource_14_valid ^ releasePipe_pipe_out_14_valid)
        tokenCheck_counter_14 <= tokenCheck_counter_14 + tokenCheck_counterChange_14;
      if (shifterValid_14) begin
        shifterReg_14_0_valid <= validSource_14_valid;
        shifterReg_14_0_bits_instructionIndex <= validSource_14_bits_instructionIndex;
        shifterReg_14_0_bits_decodeResult_orderReduce <= validSource_14_bits_decodeResult_orderReduce;
        shifterReg_14_0_bits_decodeResult_floatMul <= validSource_14_bits_decodeResult_floatMul;
        shifterReg_14_0_bits_decodeResult_fpExecutionType <= validSource_14_bits_decodeResult_fpExecutionType;
        shifterReg_14_0_bits_decodeResult_float <= validSource_14_bits_decodeResult_float;
        shifterReg_14_0_bits_decodeResult_specialSlot <= validSource_14_bits_decodeResult_specialSlot;
        shifterReg_14_0_bits_decodeResult_topUop <= validSource_14_bits_decodeResult_topUop;
        shifterReg_14_0_bits_decodeResult_popCount <= validSource_14_bits_decodeResult_popCount;
        shifterReg_14_0_bits_decodeResult_ffo <= validSource_14_bits_decodeResult_ffo;
        shifterReg_14_0_bits_decodeResult_average <= validSource_14_bits_decodeResult_average;
        shifterReg_14_0_bits_decodeResult_reverse <= validSource_14_bits_decodeResult_reverse;
        shifterReg_14_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_14_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_14_0_bits_decodeResult_scheduler <= validSource_14_bits_decodeResult_scheduler;
        shifterReg_14_0_bits_decodeResult_sReadVD <= validSource_14_bits_decodeResult_sReadVD;
        shifterReg_14_0_bits_decodeResult_vtype <= validSource_14_bits_decodeResult_vtype;
        shifterReg_14_0_bits_decodeResult_sWrite <= validSource_14_bits_decodeResult_sWrite;
        shifterReg_14_0_bits_decodeResult_crossRead <= validSource_14_bits_decodeResult_crossRead;
        shifterReg_14_0_bits_decodeResult_crossWrite <= validSource_14_bits_decodeResult_crossWrite;
        shifterReg_14_0_bits_decodeResult_maskUnit <= validSource_14_bits_decodeResult_maskUnit;
        shifterReg_14_0_bits_decodeResult_special <= validSource_14_bits_decodeResult_special;
        shifterReg_14_0_bits_decodeResult_saturate <= validSource_14_bits_decodeResult_saturate;
        shifterReg_14_0_bits_decodeResult_vwmacc <= validSource_14_bits_decodeResult_vwmacc;
        shifterReg_14_0_bits_decodeResult_readOnly <= validSource_14_bits_decodeResult_readOnly;
        shifterReg_14_0_bits_decodeResult_maskSource <= validSource_14_bits_decodeResult_maskSource;
        shifterReg_14_0_bits_decodeResult_maskDestination <= validSource_14_bits_decodeResult_maskDestination;
        shifterReg_14_0_bits_decodeResult_maskLogic <= validSource_14_bits_decodeResult_maskLogic;
        shifterReg_14_0_bits_decodeResult_uop <= validSource_14_bits_decodeResult_uop;
        shifterReg_14_0_bits_decodeResult_iota <= validSource_14_bits_decodeResult_iota;
        shifterReg_14_0_bits_decodeResult_mv <= validSource_14_bits_decodeResult_mv;
        shifterReg_14_0_bits_decodeResult_extend <= validSource_14_bits_decodeResult_extend;
        shifterReg_14_0_bits_decodeResult_unOrderWrite <= validSource_14_bits_decodeResult_unOrderWrite;
        shifterReg_14_0_bits_decodeResult_compress <= validSource_14_bits_decodeResult_compress;
        shifterReg_14_0_bits_decodeResult_gather16 <= validSource_14_bits_decodeResult_gather16;
        shifterReg_14_0_bits_decodeResult_gather <= validSource_14_bits_decodeResult_gather;
        shifterReg_14_0_bits_decodeResult_slid <= validSource_14_bits_decodeResult_slid;
        shifterReg_14_0_bits_decodeResult_targetRd <= validSource_14_bits_decodeResult_targetRd;
        shifterReg_14_0_bits_decodeResult_widenReduce <= validSource_14_bits_decodeResult_widenReduce;
        shifterReg_14_0_bits_decodeResult_red <= validSource_14_bits_decodeResult_red;
        shifterReg_14_0_bits_decodeResult_nr <= validSource_14_bits_decodeResult_nr;
        shifterReg_14_0_bits_decodeResult_itype <= validSource_14_bits_decodeResult_itype;
        shifterReg_14_0_bits_decodeResult_unsigned1 <= validSource_14_bits_decodeResult_unsigned1;
        shifterReg_14_0_bits_decodeResult_unsigned0 <= validSource_14_bits_decodeResult_unsigned0;
        shifterReg_14_0_bits_decodeResult_other <= validSource_14_bits_decodeResult_other;
        shifterReg_14_0_bits_decodeResult_multiCycle <= validSource_14_bits_decodeResult_multiCycle;
        shifterReg_14_0_bits_decodeResult_divider <= validSource_14_bits_decodeResult_divider;
        shifterReg_14_0_bits_decodeResult_multiplier <= validSource_14_bits_decodeResult_multiplier;
        shifterReg_14_0_bits_decodeResult_shift <= validSource_14_bits_decodeResult_shift;
        shifterReg_14_0_bits_decodeResult_adder <= validSource_14_bits_decodeResult_adder;
        shifterReg_14_0_bits_decodeResult_logic <= validSource_14_bits_decodeResult_logic;
        shifterReg_14_0_bits_loadStore <= validSource_14_bits_loadStore;
        shifterReg_14_0_bits_issueInst <= validSource_14_bits_issueInst;
        shifterReg_14_0_bits_store <= validSource_14_bits_store;
        shifterReg_14_0_bits_special <= validSource_14_bits_special;
        shifterReg_14_0_bits_lsWholeReg <= validSource_14_bits_lsWholeReg;
        shifterReg_14_0_bits_vs1 <= validSource_14_bits_vs1;
        shifterReg_14_0_bits_vs2 <= validSource_14_bits_vs2;
        shifterReg_14_0_bits_vd <= validSource_14_bits_vd;
        shifterReg_14_0_bits_loadStoreEEW <= validSource_14_bits_loadStoreEEW;
        shifterReg_14_0_bits_mask <= validSource_14_bits_mask;
        shifterReg_14_0_bits_segment <= validSource_14_bits_segment;
        shifterReg_14_0_bits_readFromScalar <= validSource_14_bits_readFromScalar;
        shifterReg_14_0_bits_csrInterface_vl <= validSource_14_bits_csrInterface_vl;
        shifterReg_14_0_bits_csrInterface_vStart <= validSource_14_bits_csrInterface_vStart;
        shifterReg_14_0_bits_csrInterface_vlmul <= validSource_14_bits_csrInterface_vlmul;
        shifterReg_14_0_bits_csrInterface_vSew <= validSource_14_bits_csrInterface_vSew;
        shifterReg_14_0_bits_csrInterface_vxrm <= validSource_14_bits_csrInterface_vxrm;
        shifterReg_14_0_bits_csrInterface_vta <= validSource_14_bits_csrInterface_vta;
        shifterReg_14_0_bits_csrInterface_vma <= validSource_14_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_15 <= laneVec_15_laneRequest_bits_issueInst;
      if (validSource_15_valid ^ releasePipe_pipe_out_15_valid)
        tokenCheck_counter_15 <= tokenCheck_counter_15 + tokenCheck_counterChange_15;
      if (shifterValid_15) begin
        shifterReg_15_0_valid <= validSource_15_valid;
        shifterReg_15_0_bits_instructionIndex <= validSource_15_bits_instructionIndex;
        shifterReg_15_0_bits_decodeResult_orderReduce <= validSource_15_bits_decodeResult_orderReduce;
        shifterReg_15_0_bits_decodeResult_floatMul <= validSource_15_bits_decodeResult_floatMul;
        shifterReg_15_0_bits_decodeResult_fpExecutionType <= validSource_15_bits_decodeResult_fpExecutionType;
        shifterReg_15_0_bits_decodeResult_float <= validSource_15_bits_decodeResult_float;
        shifterReg_15_0_bits_decodeResult_specialSlot <= validSource_15_bits_decodeResult_specialSlot;
        shifterReg_15_0_bits_decodeResult_topUop <= validSource_15_bits_decodeResult_topUop;
        shifterReg_15_0_bits_decodeResult_popCount <= validSource_15_bits_decodeResult_popCount;
        shifterReg_15_0_bits_decodeResult_ffo <= validSource_15_bits_decodeResult_ffo;
        shifterReg_15_0_bits_decodeResult_average <= validSource_15_bits_decodeResult_average;
        shifterReg_15_0_bits_decodeResult_reverse <= validSource_15_bits_decodeResult_reverse;
        shifterReg_15_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_15_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_15_0_bits_decodeResult_scheduler <= validSource_15_bits_decodeResult_scheduler;
        shifterReg_15_0_bits_decodeResult_sReadVD <= validSource_15_bits_decodeResult_sReadVD;
        shifterReg_15_0_bits_decodeResult_vtype <= validSource_15_bits_decodeResult_vtype;
        shifterReg_15_0_bits_decodeResult_sWrite <= validSource_15_bits_decodeResult_sWrite;
        shifterReg_15_0_bits_decodeResult_crossRead <= validSource_15_bits_decodeResult_crossRead;
        shifterReg_15_0_bits_decodeResult_crossWrite <= validSource_15_bits_decodeResult_crossWrite;
        shifterReg_15_0_bits_decodeResult_maskUnit <= validSource_15_bits_decodeResult_maskUnit;
        shifterReg_15_0_bits_decodeResult_special <= validSource_15_bits_decodeResult_special;
        shifterReg_15_0_bits_decodeResult_saturate <= validSource_15_bits_decodeResult_saturate;
        shifterReg_15_0_bits_decodeResult_vwmacc <= validSource_15_bits_decodeResult_vwmacc;
        shifterReg_15_0_bits_decodeResult_readOnly <= validSource_15_bits_decodeResult_readOnly;
        shifterReg_15_0_bits_decodeResult_maskSource <= validSource_15_bits_decodeResult_maskSource;
        shifterReg_15_0_bits_decodeResult_maskDestination <= validSource_15_bits_decodeResult_maskDestination;
        shifterReg_15_0_bits_decodeResult_maskLogic <= validSource_15_bits_decodeResult_maskLogic;
        shifterReg_15_0_bits_decodeResult_uop <= validSource_15_bits_decodeResult_uop;
        shifterReg_15_0_bits_decodeResult_iota <= validSource_15_bits_decodeResult_iota;
        shifterReg_15_0_bits_decodeResult_mv <= validSource_15_bits_decodeResult_mv;
        shifterReg_15_0_bits_decodeResult_extend <= validSource_15_bits_decodeResult_extend;
        shifterReg_15_0_bits_decodeResult_unOrderWrite <= validSource_15_bits_decodeResult_unOrderWrite;
        shifterReg_15_0_bits_decodeResult_compress <= validSource_15_bits_decodeResult_compress;
        shifterReg_15_0_bits_decodeResult_gather16 <= validSource_15_bits_decodeResult_gather16;
        shifterReg_15_0_bits_decodeResult_gather <= validSource_15_bits_decodeResult_gather;
        shifterReg_15_0_bits_decodeResult_slid <= validSource_15_bits_decodeResult_slid;
        shifterReg_15_0_bits_decodeResult_targetRd <= validSource_15_bits_decodeResult_targetRd;
        shifterReg_15_0_bits_decodeResult_widenReduce <= validSource_15_bits_decodeResult_widenReduce;
        shifterReg_15_0_bits_decodeResult_red <= validSource_15_bits_decodeResult_red;
        shifterReg_15_0_bits_decodeResult_nr <= validSource_15_bits_decodeResult_nr;
        shifterReg_15_0_bits_decodeResult_itype <= validSource_15_bits_decodeResult_itype;
        shifterReg_15_0_bits_decodeResult_unsigned1 <= validSource_15_bits_decodeResult_unsigned1;
        shifterReg_15_0_bits_decodeResult_unsigned0 <= validSource_15_bits_decodeResult_unsigned0;
        shifterReg_15_0_bits_decodeResult_other <= validSource_15_bits_decodeResult_other;
        shifterReg_15_0_bits_decodeResult_multiCycle <= validSource_15_bits_decodeResult_multiCycle;
        shifterReg_15_0_bits_decodeResult_divider <= validSource_15_bits_decodeResult_divider;
        shifterReg_15_0_bits_decodeResult_multiplier <= validSource_15_bits_decodeResult_multiplier;
        shifterReg_15_0_bits_decodeResult_shift <= validSource_15_bits_decodeResult_shift;
        shifterReg_15_0_bits_decodeResult_adder <= validSource_15_bits_decodeResult_adder;
        shifterReg_15_0_bits_decodeResult_logic <= validSource_15_bits_decodeResult_logic;
        shifterReg_15_0_bits_loadStore <= validSource_15_bits_loadStore;
        shifterReg_15_0_bits_issueInst <= validSource_15_bits_issueInst;
        shifterReg_15_0_bits_store <= validSource_15_bits_store;
        shifterReg_15_0_bits_special <= validSource_15_bits_special;
        shifterReg_15_0_bits_lsWholeReg <= validSource_15_bits_lsWholeReg;
        shifterReg_15_0_bits_vs1 <= validSource_15_bits_vs1;
        shifterReg_15_0_bits_vs2 <= validSource_15_bits_vs2;
        shifterReg_15_0_bits_vd <= validSource_15_bits_vd;
        shifterReg_15_0_bits_loadStoreEEW <= validSource_15_bits_loadStoreEEW;
        shifterReg_15_0_bits_mask <= validSource_15_bits_mask;
        shifterReg_15_0_bits_segment <= validSource_15_bits_segment;
        shifterReg_15_0_bits_readFromScalar <= validSource_15_bits_readFromScalar;
        shifterReg_15_0_bits_csrInterface_vl <= validSource_15_bits_csrInterface_vl;
        shifterReg_15_0_bits_csrInterface_vStart <= validSource_15_bits_csrInterface_vStart;
        shifterReg_15_0_bits_csrInterface_vlmul <= validSource_15_bits_csrInterface_vlmul;
        shifterReg_15_0_bits_csrInterface_vSew <= validSource_15_bits_csrInterface_vSew;
        shifterReg_15_0_bits_csrInterface_vxrm <= validSource_15_bits_csrInterface_vxrm;
        shifterReg_15_0_bits_csrInterface_vta <= validSource_15_bits_csrInterface_vta;
        shifterReg_15_0_bits_csrInterface_vma <= validSource_15_bits_csrInterface_vma;
      end
      sinkVec_releasePipe_pipe_v <= sinkVec_sinkWire_ready & sinkVec_sinkWire_valid;
      if (sinkVec_validSource_valid ^ sinkVec_releasePipe_pipe_out_valid)
        sinkVec_tokenCheck_counter <= sinkVec_tokenCheck_counter + sinkVec_tokenCheck_counterChange;
      if (sinkVec_shifterValid) begin
        sinkVec_shifterReg_0_valid <= sinkVec_validSource_valid;
        sinkVec_shifterReg_0_bits_vs <= sinkVec_validSource_bits_vs;
        sinkVec_shifterReg_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_0_bits_offset <= sinkVec_validSource_bits_offset;
        sinkVec_shifterReg_0_bits_instructionIndex <= sinkVec_validSource_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_1 <= sinkVec_sinkWire_1_ready & sinkVec_sinkWire_1_valid;
      if (sinkVec_validSource_1_valid ^ sinkVec_releasePipe_pipe_out_1_valid)
        sinkVec_tokenCheck_counter_1 <= sinkVec_tokenCheck_counter_1 + sinkVec_tokenCheck_counterChange_1;
      if (sinkVec_shifterValid_1) begin
        sinkVec_shifterReg_1_0_valid <= sinkVec_validSource_1_valid;
        sinkVec_shifterReg_1_0_bits_vs <= sinkVec_validSource_1_bits_vs;
        sinkVec_shifterReg_1_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_1_0_bits_offset <= sinkVec_validSource_1_bits_offset;
        sinkVec_shifterReg_1_0_bits_instructionIndex <= sinkVec_validSource_1_bits_instructionIndex;
      end
      maskUnitFirst <= tryToRead & ~(sinkWire_ready & sinkWire_valid) ^ maskUnitFirst;
      accessDataValid_pipe_v <= sinkVec_0_ready & sinkVec_0_valid;
      accessDataValid_pipe_pipe_v <= accessDataValid_pipe_v;
      if (shifterValid_16) begin
        shifterReg_16_0_valid <= accessDataSource_valid;
        shifterReg_16_0_bits <= accessDataSource_bits;
      end
      accessDataValid_pipe_v_1 <= sinkVec_1_ready & sinkVec_1_valid;
      accessDataValid_pipe_pipe_v_1 <= accessDataValid_pipe_v_1;
      if (shifterValid_17) begin
        shifterReg_17_0_valid <= accessDataSource_1_valid;
        shifterReg_17_0_bits <= accessDataSource_1_bits;
      end
      sinkVec_releasePipe_pipe_v_2 <= sinkVec_sinkWire_2_ready & sinkVec_sinkWire_2_valid;
      if (sinkVec_validSource_2_valid ^ sinkVec_releasePipe_pipe_out_2_valid)
        sinkVec_tokenCheck_counter_2 <= sinkVec_tokenCheck_counter_2 + sinkVec_tokenCheck_counterChange_2;
      if (sinkVec_shifterValid_2) begin
        sinkVec_shifterReg_2_0_valid <= sinkVec_validSource_2_valid;
        sinkVec_shifterReg_2_0_bits_vd <= sinkVec_validSource_2_bits_vd;
        sinkVec_shifterReg_2_0_bits_offset <= sinkVec_validSource_2_bits_offset;
        sinkVec_shifterReg_2_0_bits_mask <= sinkVec_validSource_2_bits_mask;
        sinkVec_shifterReg_2_0_bits_data <= sinkVec_validSource_2_bits_data;
        sinkVec_shifterReg_2_0_bits_instructionIndex <= sinkVec_validSource_2_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_3 <= sinkVec_sinkWire_3_ready & sinkVec_sinkWire_3_valid;
      if (sinkVec_validSource_3_valid ^ sinkVec_releasePipe_pipe_out_3_valid)
        sinkVec_tokenCheck_counter_3 <= sinkVec_tokenCheck_counter_3 + sinkVec_tokenCheck_counterChange_3;
      if (sinkVec_shifterValid_3) begin
        sinkVec_shifterReg_3_0_valid <= sinkVec_validSource_3_valid;
        sinkVec_shifterReg_3_0_bits_vd <= sinkVec_validSource_3_bits_vd;
        sinkVec_shifterReg_3_0_bits_offset <= sinkVec_validSource_3_bits_offset;
        sinkVec_shifterReg_3_0_bits_mask <= sinkVec_validSource_3_bits_mask;
        sinkVec_shifterReg_3_0_bits_data <= sinkVec_validSource_3_bits_data;
        sinkVec_shifterReg_3_0_bits_last <= sinkVec_validSource_3_bits_last;
        sinkVec_shifterReg_3_0_bits_instructionIndex <= sinkVec_validSource_3_bits_instructionIndex;
      end
      maskUnitFirst_1 <= tryToRead_1 & ~(sinkWire_1_ready & sinkWire_1_valid) ^ maskUnitFirst_1;
      view__writeRelease_0_pipe_v <= sinkVec_1_0_ready & sinkVec_1_0_valid;
      pipe_v <= sinkVec_1_1_ready & sinkVec_1_1_valid;
      instructionFinishedPipe_pipe_v <= 1'h1;
      pipe_v_1 <= 1'h1;
      pipe_pipe_v <= pipe_v_1;
      view__laneMaskSelect_0_pipe_v <= 1'h1;
      view__laneMaskSelect_0_pipe_pipe_v <= view__laneMaskSelect_0_pipe_v;
      view__laneMaskSewSelect_0_pipe_v <= 1'h1;
      view__laneMaskSewSelect_0_pipe_pipe_v <= view__laneMaskSewSelect_0_pipe_v;
      lsuLastPipe_pipe_v <= 1'h1;
      maskLastPipe_pipe_v <= 1'h1;
      pipe_v_2 <= 1'h1;
      sinkVec_releasePipe_pipe_v_4 <= sinkVec_sinkWire_4_ready & sinkVec_sinkWire_4_valid;
      if (sinkVec_validSource_4_valid ^ sinkVec_releasePipe_pipe_out_4_valid)
        sinkVec_tokenCheck_counter_4 <= sinkVec_tokenCheck_counter_4 + sinkVec_tokenCheck_counterChange_4;
      if (sinkVec_shifterValid_4) begin
        sinkVec_shifterReg_4_0_valid <= sinkVec_validSource_4_valid;
        sinkVec_shifterReg_4_0_bits_vs <= sinkVec_validSource_4_bits_vs;
        sinkVec_shifterReg_4_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_4_0_bits_offset <= sinkVec_validSource_4_bits_offset;
        sinkVec_shifterReg_4_0_bits_instructionIndex <= sinkVec_validSource_4_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_5 <= sinkVec_sinkWire_5_ready & sinkVec_sinkWire_5_valid;
      if (sinkVec_validSource_5_valid ^ sinkVec_releasePipe_pipe_out_5_valid)
        sinkVec_tokenCheck_counter_5 <= sinkVec_tokenCheck_counter_5 + sinkVec_tokenCheck_counterChange_5;
      if (sinkVec_shifterValid_5) begin
        sinkVec_shifterReg_5_0_valid <= sinkVec_validSource_5_valid;
        sinkVec_shifterReg_5_0_bits_vs <= sinkVec_validSource_5_bits_vs;
        sinkVec_shifterReg_5_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_5_0_bits_offset <= sinkVec_validSource_5_bits_offset;
        sinkVec_shifterReg_5_0_bits_instructionIndex <= sinkVec_validSource_5_bits_instructionIndex;
      end
      maskUnitFirst_2 <= tryToRead_2 & ~(sinkWire_2_ready & sinkWire_2_valid) ^ maskUnitFirst_2;
      accessDataValid_pipe_v_2 <= sinkVec_2_0_ready & sinkVec_2_0_valid;
      accessDataValid_pipe_pipe_v_2 <= accessDataValid_pipe_v_2;
      if (shifterValid_18) begin
        shifterReg_18_0_valid <= accessDataSource_2_valid;
        shifterReg_18_0_bits <= accessDataSource_2_bits;
      end
      accessDataValid_pipe_v_3 <= sinkVec_2_1_ready & sinkVec_2_1_valid;
      accessDataValid_pipe_pipe_v_3 <= accessDataValid_pipe_v_3;
      if (shifterValid_19) begin
        shifterReg_19_0_valid <= accessDataSource_3_valid;
        shifterReg_19_0_bits <= accessDataSource_3_bits;
      end
      sinkVec_releasePipe_pipe_v_6 <= sinkVec_sinkWire_6_ready & sinkVec_sinkWire_6_valid;
      if (sinkVec_validSource_6_valid ^ sinkVec_releasePipe_pipe_out_6_valid)
        sinkVec_tokenCheck_counter_6 <= sinkVec_tokenCheck_counter_6 + sinkVec_tokenCheck_counterChange_6;
      if (sinkVec_shifterValid_6) begin
        sinkVec_shifterReg_6_0_valid <= sinkVec_validSource_6_valid;
        sinkVec_shifterReg_6_0_bits_vd <= sinkVec_validSource_6_bits_vd;
        sinkVec_shifterReg_6_0_bits_offset <= sinkVec_validSource_6_bits_offset;
        sinkVec_shifterReg_6_0_bits_mask <= sinkVec_validSource_6_bits_mask;
        sinkVec_shifterReg_6_0_bits_data <= sinkVec_validSource_6_bits_data;
        sinkVec_shifterReg_6_0_bits_instructionIndex <= sinkVec_validSource_6_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_7 <= sinkVec_sinkWire_7_ready & sinkVec_sinkWire_7_valid;
      if (sinkVec_validSource_7_valid ^ sinkVec_releasePipe_pipe_out_7_valid)
        sinkVec_tokenCheck_counter_7 <= sinkVec_tokenCheck_counter_7 + sinkVec_tokenCheck_counterChange_7;
      if (sinkVec_shifterValid_7) begin
        sinkVec_shifterReg_7_0_valid <= sinkVec_validSource_7_valid;
        sinkVec_shifterReg_7_0_bits_vd <= sinkVec_validSource_7_bits_vd;
        sinkVec_shifterReg_7_0_bits_offset <= sinkVec_validSource_7_bits_offset;
        sinkVec_shifterReg_7_0_bits_mask <= sinkVec_validSource_7_bits_mask;
        sinkVec_shifterReg_7_0_bits_data <= sinkVec_validSource_7_bits_data;
        sinkVec_shifterReg_7_0_bits_last <= sinkVec_validSource_7_bits_last;
        sinkVec_shifterReg_7_0_bits_instructionIndex <= sinkVec_validSource_7_bits_instructionIndex;
      end
      maskUnitFirst_3 <= tryToRead_3 & ~(sinkWire_3_ready & sinkWire_3_valid) ^ maskUnitFirst_3;
      view__writeRelease_1_pipe_v <= sinkVec_3_0_ready & sinkVec_3_0_valid;
      pipe_v_3 <= sinkVec_3_1_ready & sinkVec_3_1_valid;
      instructionFinishedPipe_pipe_v_1 <= 1'h1;
      pipe_v_4 <= 1'h1;
      pipe_pipe_v_1 <= pipe_v_4;
      view__laneMaskSelect_1_pipe_v <= 1'h1;
      view__laneMaskSelect_1_pipe_pipe_v <= view__laneMaskSelect_1_pipe_v;
      view__laneMaskSewSelect_1_pipe_v <= 1'h1;
      view__laneMaskSewSelect_1_pipe_pipe_v <= view__laneMaskSewSelect_1_pipe_v;
      lsuLastPipe_pipe_v_1 <= 1'h1;
      maskLastPipe_pipe_v_1 <= 1'h1;
      pipe_v_5 <= 1'h1;
      sinkVec_releasePipe_pipe_v_8 <= sinkVec_sinkWire_8_ready & sinkVec_sinkWire_8_valid;
      if (sinkVec_validSource_8_valid ^ sinkVec_releasePipe_pipe_out_8_valid)
        sinkVec_tokenCheck_counter_8 <= sinkVec_tokenCheck_counter_8 + sinkVec_tokenCheck_counterChange_8;
      if (sinkVec_shifterValid_8) begin
        sinkVec_shifterReg_8_0_valid <= sinkVec_validSource_8_valid;
        sinkVec_shifterReg_8_0_bits_vs <= sinkVec_validSource_8_bits_vs;
        sinkVec_shifterReg_8_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_8_0_bits_offset <= sinkVec_validSource_8_bits_offset;
        sinkVec_shifterReg_8_0_bits_instructionIndex <= sinkVec_validSource_8_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_9 <= sinkVec_sinkWire_9_ready & sinkVec_sinkWire_9_valid;
      if (sinkVec_validSource_9_valid ^ sinkVec_releasePipe_pipe_out_9_valid)
        sinkVec_tokenCheck_counter_9 <= sinkVec_tokenCheck_counter_9 + sinkVec_tokenCheck_counterChange_9;
      if (sinkVec_shifterValid_9) begin
        sinkVec_shifterReg_9_0_valid <= sinkVec_validSource_9_valid;
        sinkVec_shifterReg_9_0_bits_vs <= sinkVec_validSource_9_bits_vs;
        sinkVec_shifterReg_9_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_9_0_bits_offset <= sinkVec_validSource_9_bits_offset;
        sinkVec_shifterReg_9_0_bits_instructionIndex <= sinkVec_validSource_9_bits_instructionIndex;
      end
      maskUnitFirst_4 <= tryToRead_4 & ~(sinkWire_4_ready & sinkWire_4_valid) ^ maskUnitFirst_4;
      accessDataValid_pipe_v_4 <= sinkVec_4_0_ready & sinkVec_4_0_valid;
      accessDataValid_pipe_pipe_v_4 <= accessDataValid_pipe_v_4;
      if (shifterValid_20) begin
        shifterReg_20_0_valid <= accessDataSource_4_valid;
        shifterReg_20_0_bits <= accessDataSource_4_bits;
      end
      accessDataValid_pipe_v_5 <= sinkVec_4_1_ready & sinkVec_4_1_valid;
      accessDataValid_pipe_pipe_v_5 <= accessDataValid_pipe_v_5;
      if (shifterValid_21) begin
        shifterReg_21_0_valid <= accessDataSource_5_valid;
        shifterReg_21_0_bits <= accessDataSource_5_bits;
      end
      sinkVec_releasePipe_pipe_v_10 <= sinkVec_sinkWire_10_ready & sinkVec_sinkWire_10_valid;
      if (sinkVec_validSource_10_valid ^ sinkVec_releasePipe_pipe_out_10_valid)
        sinkVec_tokenCheck_counter_10 <= sinkVec_tokenCheck_counter_10 + sinkVec_tokenCheck_counterChange_10;
      if (sinkVec_shifterValid_10) begin
        sinkVec_shifterReg_10_0_valid <= sinkVec_validSource_10_valid;
        sinkVec_shifterReg_10_0_bits_vd <= sinkVec_validSource_10_bits_vd;
        sinkVec_shifterReg_10_0_bits_offset <= sinkVec_validSource_10_bits_offset;
        sinkVec_shifterReg_10_0_bits_mask <= sinkVec_validSource_10_bits_mask;
        sinkVec_shifterReg_10_0_bits_data <= sinkVec_validSource_10_bits_data;
        sinkVec_shifterReg_10_0_bits_instructionIndex <= sinkVec_validSource_10_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_11 <= sinkVec_sinkWire_11_ready & sinkVec_sinkWire_11_valid;
      if (sinkVec_validSource_11_valid ^ sinkVec_releasePipe_pipe_out_11_valid)
        sinkVec_tokenCheck_counter_11 <= sinkVec_tokenCheck_counter_11 + sinkVec_tokenCheck_counterChange_11;
      if (sinkVec_shifterValid_11) begin
        sinkVec_shifterReg_11_0_valid <= sinkVec_validSource_11_valid;
        sinkVec_shifterReg_11_0_bits_vd <= sinkVec_validSource_11_bits_vd;
        sinkVec_shifterReg_11_0_bits_offset <= sinkVec_validSource_11_bits_offset;
        sinkVec_shifterReg_11_0_bits_mask <= sinkVec_validSource_11_bits_mask;
        sinkVec_shifterReg_11_0_bits_data <= sinkVec_validSource_11_bits_data;
        sinkVec_shifterReg_11_0_bits_last <= sinkVec_validSource_11_bits_last;
        sinkVec_shifterReg_11_0_bits_instructionIndex <= sinkVec_validSource_11_bits_instructionIndex;
      end
      maskUnitFirst_5 <= tryToRead_5 & ~(sinkWire_5_ready & sinkWire_5_valid) ^ maskUnitFirst_5;
      view__writeRelease_2_pipe_v <= sinkVec_5_0_ready & sinkVec_5_0_valid;
      pipe_v_6 <= sinkVec_5_1_ready & sinkVec_5_1_valid;
      instructionFinishedPipe_pipe_v_2 <= 1'h1;
      pipe_v_7 <= 1'h1;
      pipe_pipe_v_2 <= pipe_v_7;
      view__laneMaskSelect_2_pipe_v <= 1'h1;
      view__laneMaskSelect_2_pipe_pipe_v <= view__laneMaskSelect_2_pipe_v;
      view__laneMaskSewSelect_2_pipe_v <= 1'h1;
      view__laneMaskSewSelect_2_pipe_pipe_v <= view__laneMaskSewSelect_2_pipe_v;
      lsuLastPipe_pipe_v_2 <= 1'h1;
      maskLastPipe_pipe_v_2 <= 1'h1;
      pipe_v_8 <= 1'h1;
      sinkVec_releasePipe_pipe_v_12 <= sinkVec_sinkWire_12_ready & sinkVec_sinkWire_12_valid;
      if (sinkVec_validSource_12_valid ^ sinkVec_releasePipe_pipe_out_12_valid)
        sinkVec_tokenCheck_counter_12 <= sinkVec_tokenCheck_counter_12 + sinkVec_tokenCheck_counterChange_12;
      if (sinkVec_shifterValid_12) begin
        sinkVec_shifterReg_12_0_valid <= sinkVec_validSource_12_valid;
        sinkVec_shifterReg_12_0_bits_vs <= sinkVec_validSource_12_bits_vs;
        sinkVec_shifterReg_12_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_12_0_bits_offset <= sinkVec_validSource_12_bits_offset;
        sinkVec_shifterReg_12_0_bits_instructionIndex <= sinkVec_validSource_12_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_13 <= sinkVec_sinkWire_13_ready & sinkVec_sinkWire_13_valid;
      if (sinkVec_validSource_13_valid ^ sinkVec_releasePipe_pipe_out_13_valid)
        sinkVec_tokenCheck_counter_13 <= sinkVec_tokenCheck_counter_13 + sinkVec_tokenCheck_counterChange_13;
      if (sinkVec_shifterValid_13) begin
        sinkVec_shifterReg_13_0_valid <= sinkVec_validSource_13_valid;
        sinkVec_shifterReg_13_0_bits_vs <= sinkVec_validSource_13_bits_vs;
        sinkVec_shifterReg_13_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_13_0_bits_offset <= sinkVec_validSource_13_bits_offset;
        sinkVec_shifterReg_13_0_bits_instructionIndex <= sinkVec_validSource_13_bits_instructionIndex;
      end
      maskUnitFirst_6 <= tryToRead_6 & ~(sinkWire_6_ready & sinkWire_6_valid) ^ maskUnitFirst_6;
      accessDataValid_pipe_v_6 <= sinkVec_6_0_ready & sinkVec_6_0_valid;
      accessDataValid_pipe_pipe_v_6 <= accessDataValid_pipe_v_6;
      if (shifterValid_22) begin
        shifterReg_22_0_valid <= accessDataSource_6_valid;
        shifterReg_22_0_bits <= accessDataSource_6_bits;
      end
      accessDataValid_pipe_v_7 <= sinkVec_6_1_ready & sinkVec_6_1_valid;
      accessDataValid_pipe_pipe_v_7 <= accessDataValid_pipe_v_7;
      if (shifterValid_23) begin
        shifterReg_23_0_valid <= accessDataSource_7_valid;
        shifterReg_23_0_bits <= accessDataSource_7_bits;
      end
      sinkVec_releasePipe_pipe_v_14 <= sinkVec_sinkWire_14_ready & sinkVec_sinkWire_14_valid;
      if (sinkVec_validSource_14_valid ^ sinkVec_releasePipe_pipe_out_14_valid)
        sinkVec_tokenCheck_counter_14 <= sinkVec_tokenCheck_counter_14 + sinkVec_tokenCheck_counterChange_14;
      if (sinkVec_shifterValid_14) begin
        sinkVec_shifterReg_14_0_valid <= sinkVec_validSource_14_valid;
        sinkVec_shifterReg_14_0_bits_vd <= sinkVec_validSource_14_bits_vd;
        sinkVec_shifterReg_14_0_bits_offset <= sinkVec_validSource_14_bits_offset;
        sinkVec_shifterReg_14_0_bits_mask <= sinkVec_validSource_14_bits_mask;
        sinkVec_shifterReg_14_0_bits_data <= sinkVec_validSource_14_bits_data;
        sinkVec_shifterReg_14_0_bits_instructionIndex <= sinkVec_validSource_14_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_15 <= sinkVec_sinkWire_15_ready & sinkVec_sinkWire_15_valid;
      if (sinkVec_validSource_15_valid ^ sinkVec_releasePipe_pipe_out_15_valid)
        sinkVec_tokenCheck_counter_15 <= sinkVec_tokenCheck_counter_15 + sinkVec_tokenCheck_counterChange_15;
      if (sinkVec_shifterValid_15) begin
        sinkVec_shifterReg_15_0_valid <= sinkVec_validSource_15_valid;
        sinkVec_shifterReg_15_0_bits_vd <= sinkVec_validSource_15_bits_vd;
        sinkVec_shifterReg_15_0_bits_offset <= sinkVec_validSource_15_bits_offset;
        sinkVec_shifterReg_15_0_bits_mask <= sinkVec_validSource_15_bits_mask;
        sinkVec_shifterReg_15_0_bits_data <= sinkVec_validSource_15_bits_data;
        sinkVec_shifterReg_15_0_bits_last <= sinkVec_validSource_15_bits_last;
        sinkVec_shifterReg_15_0_bits_instructionIndex <= sinkVec_validSource_15_bits_instructionIndex;
      end
      maskUnitFirst_7 <= tryToRead_7 & ~(sinkWire_7_ready & sinkWire_7_valid) ^ maskUnitFirst_7;
      view__writeRelease_3_pipe_v <= sinkVec_7_0_ready & sinkVec_7_0_valid;
      pipe_v_9 <= sinkVec_7_1_ready & sinkVec_7_1_valid;
      instructionFinishedPipe_pipe_v_3 <= 1'h1;
      pipe_v_10 <= 1'h1;
      pipe_pipe_v_3 <= pipe_v_10;
      view__laneMaskSelect_3_pipe_v <= 1'h1;
      view__laneMaskSelect_3_pipe_pipe_v <= view__laneMaskSelect_3_pipe_v;
      view__laneMaskSewSelect_3_pipe_v <= 1'h1;
      view__laneMaskSewSelect_3_pipe_pipe_v <= view__laneMaskSewSelect_3_pipe_v;
      lsuLastPipe_pipe_v_3 <= 1'h1;
      maskLastPipe_pipe_v_3 <= 1'h1;
      pipe_v_11 <= 1'h1;
      sinkVec_releasePipe_pipe_v_16 <= sinkVec_sinkWire_16_ready & sinkVec_sinkWire_16_valid;
      if (sinkVec_validSource_16_valid ^ sinkVec_releasePipe_pipe_out_16_valid)
        sinkVec_tokenCheck_counter_16 <= sinkVec_tokenCheck_counter_16 + sinkVec_tokenCheck_counterChange_16;
      if (sinkVec_shifterValid_16) begin
        sinkVec_shifterReg_16_0_valid <= sinkVec_validSource_16_valid;
        sinkVec_shifterReg_16_0_bits_vs <= sinkVec_validSource_16_bits_vs;
        sinkVec_shifterReg_16_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_16_0_bits_offset <= sinkVec_validSource_16_bits_offset;
        sinkVec_shifterReg_16_0_bits_instructionIndex <= sinkVec_validSource_16_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_17 <= sinkVec_sinkWire_17_ready & sinkVec_sinkWire_17_valid;
      if (sinkVec_validSource_17_valid ^ sinkVec_releasePipe_pipe_out_17_valid)
        sinkVec_tokenCheck_counter_17 <= sinkVec_tokenCheck_counter_17 + sinkVec_tokenCheck_counterChange_17;
      if (sinkVec_shifterValid_17) begin
        sinkVec_shifterReg_17_0_valid <= sinkVec_validSource_17_valid;
        sinkVec_shifterReg_17_0_bits_vs <= sinkVec_validSource_17_bits_vs;
        sinkVec_shifterReg_17_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_17_0_bits_offset <= sinkVec_validSource_17_bits_offset;
        sinkVec_shifterReg_17_0_bits_instructionIndex <= sinkVec_validSource_17_bits_instructionIndex;
      end
      maskUnitFirst_8 <= tryToRead_8 & ~(sinkWire_8_ready & sinkWire_8_valid) ^ maskUnitFirst_8;
      accessDataValid_pipe_v_8 <= sinkVec_8_0_ready & sinkVec_8_0_valid;
      accessDataValid_pipe_pipe_v_8 <= accessDataValid_pipe_v_8;
      if (shifterValid_24) begin
        shifterReg_24_0_valid <= accessDataSource_8_valid;
        shifterReg_24_0_bits <= accessDataSource_8_bits;
      end
      accessDataValid_pipe_v_9 <= sinkVec_8_1_ready & sinkVec_8_1_valid;
      accessDataValid_pipe_pipe_v_9 <= accessDataValid_pipe_v_9;
      if (shifterValid_25) begin
        shifterReg_25_0_valid <= accessDataSource_9_valid;
        shifterReg_25_0_bits <= accessDataSource_9_bits;
      end
      sinkVec_releasePipe_pipe_v_18 <= sinkVec_sinkWire_18_ready & sinkVec_sinkWire_18_valid;
      if (sinkVec_validSource_18_valid ^ sinkVec_releasePipe_pipe_out_18_valid)
        sinkVec_tokenCheck_counter_18 <= sinkVec_tokenCheck_counter_18 + sinkVec_tokenCheck_counterChange_18;
      if (sinkVec_shifterValid_18) begin
        sinkVec_shifterReg_18_0_valid <= sinkVec_validSource_18_valid;
        sinkVec_shifterReg_18_0_bits_vd <= sinkVec_validSource_18_bits_vd;
        sinkVec_shifterReg_18_0_bits_offset <= sinkVec_validSource_18_bits_offset;
        sinkVec_shifterReg_18_0_bits_mask <= sinkVec_validSource_18_bits_mask;
        sinkVec_shifterReg_18_0_bits_data <= sinkVec_validSource_18_bits_data;
        sinkVec_shifterReg_18_0_bits_instructionIndex <= sinkVec_validSource_18_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_19 <= sinkVec_sinkWire_19_ready & sinkVec_sinkWire_19_valid;
      if (sinkVec_validSource_19_valid ^ sinkVec_releasePipe_pipe_out_19_valid)
        sinkVec_tokenCheck_counter_19 <= sinkVec_tokenCheck_counter_19 + sinkVec_tokenCheck_counterChange_19;
      if (sinkVec_shifterValid_19) begin
        sinkVec_shifterReg_19_0_valid <= sinkVec_validSource_19_valid;
        sinkVec_shifterReg_19_0_bits_vd <= sinkVec_validSource_19_bits_vd;
        sinkVec_shifterReg_19_0_bits_offset <= sinkVec_validSource_19_bits_offset;
        sinkVec_shifterReg_19_0_bits_mask <= sinkVec_validSource_19_bits_mask;
        sinkVec_shifterReg_19_0_bits_data <= sinkVec_validSource_19_bits_data;
        sinkVec_shifterReg_19_0_bits_last <= sinkVec_validSource_19_bits_last;
        sinkVec_shifterReg_19_0_bits_instructionIndex <= sinkVec_validSource_19_bits_instructionIndex;
      end
      maskUnitFirst_9 <= tryToRead_9 & ~(sinkWire_9_ready & sinkWire_9_valid) ^ maskUnitFirst_9;
      view__writeRelease_4_pipe_v <= sinkVec_9_0_ready & sinkVec_9_0_valid;
      pipe_v_12 <= sinkVec_9_1_ready & sinkVec_9_1_valid;
      instructionFinishedPipe_pipe_v_4 <= 1'h1;
      pipe_v_13 <= 1'h1;
      pipe_pipe_v_4 <= pipe_v_13;
      view__laneMaskSelect_4_pipe_v <= 1'h1;
      view__laneMaskSelect_4_pipe_pipe_v <= view__laneMaskSelect_4_pipe_v;
      view__laneMaskSewSelect_4_pipe_v <= 1'h1;
      view__laneMaskSewSelect_4_pipe_pipe_v <= view__laneMaskSewSelect_4_pipe_v;
      lsuLastPipe_pipe_v_4 <= 1'h1;
      maskLastPipe_pipe_v_4 <= 1'h1;
      pipe_v_14 <= 1'h1;
      sinkVec_releasePipe_pipe_v_20 <= sinkVec_sinkWire_20_ready & sinkVec_sinkWire_20_valid;
      if (sinkVec_validSource_20_valid ^ sinkVec_releasePipe_pipe_out_20_valid)
        sinkVec_tokenCheck_counter_20 <= sinkVec_tokenCheck_counter_20 + sinkVec_tokenCheck_counterChange_20;
      if (sinkVec_shifterValid_20) begin
        sinkVec_shifterReg_20_0_valid <= sinkVec_validSource_20_valid;
        sinkVec_shifterReg_20_0_bits_vs <= sinkVec_validSource_20_bits_vs;
        sinkVec_shifterReg_20_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_20_0_bits_offset <= sinkVec_validSource_20_bits_offset;
        sinkVec_shifterReg_20_0_bits_instructionIndex <= sinkVec_validSource_20_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_21 <= sinkVec_sinkWire_21_ready & sinkVec_sinkWire_21_valid;
      if (sinkVec_validSource_21_valid ^ sinkVec_releasePipe_pipe_out_21_valid)
        sinkVec_tokenCheck_counter_21 <= sinkVec_tokenCheck_counter_21 + sinkVec_tokenCheck_counterChange_21;
      if (sinkVec_shifterValid_21) begin
        sinkVec_shifterReg_21_0_valid <= sinkVec_validSource_21_valid;
        sinkVec_shifterReg_21_0_bits_vs <= sinkVec_validSource_21_bits_vs;
        sinkVec_shifterReg_21_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_21_0_bits_offset <= sinkVec_validSource_21_bits_offset;
        sinkVec_shifterReg_21_0_bits_instructionIndex <= sinkVec_validSource_21_bits_instructionIndex;
      end
      maskUnitFirst_10 <= tryToRead_10 & ~(sinkWire_10_ready & sinkWire_10_valid) ^ maskUnitFirst_10;
      accessDataValid_pipe_v_10 <= sinkVec_10_0_ready & sinkVec_10_0_valid;
      accessDataValid_pipe_pipe_v_10 <= accessDataValid_pipe_v_10;
      if (shifterValid_26) begin
        shifterReg_26_0_valid <= accessDataSource_10_valid;
        shifterReg_26_0_bits <= accessDataSource_10_bits;
      end
      accessDataValid_pipe_v_11 <= sinkVec_10_1_ready & sinkVec_10_1_valid;
      accessDataValid_pipe_pipe_v_11 <= accessDataValid_pipe_v_11;
      if (shifterValid_27) begin
        shifterReg_27_0_valid <= accessDataSource_11_valid;
        shifterReg_27_0_bits <= accessDataSource_11_bits;
      end
      sinkVec_releasePipe_pipe_v_22 <= sinkVec_sinkWire_22_ready & sinkVec_sinkWire_22_valid;
      if (sinkVec_validSource_22_valid ^ sinkVec_releasePipe_pipe_out_22_valid)
        sinkVec_tokenCheck_counter_22 <= sinkVec_tokenCheck_counter_22 + sinkVec_tokenCheck_counterChange_22;
      if (sinkVec_shifterValid_22) begin
        sinkVec_shifterReg_22_0_valid <= sinkVec_validSource_22_valid;
        sinkVec_shifterReg_22_0_bits_vd <= sinkVec_validSource_22_bits_vd;
        sinkVec_shifterReg_22_0_bits_offset <= sinkVec_validSource_22_bits_offset;
        sinkVec_shifterReg_22_0_bits_mask <= sinkVec_validSource_22_bits_mask;
        sinkVec_shifterReg_22_0_bits_data <= sinkVec_validSource_22_bits_data;
        sinkVec_shifterReg_22_0_bits_instructionIndex <= sinkVec_validSource_22_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_23 <= sinkVec_sinkWire_23_ready & sinkVec_sinkWire_23_valid;
      if (sinkVec_validSource_23_valid ^ sinkVec_releasePipe_pipe_out_23_valid)
        sinkVec_tokenCheck_counter_23 <= sinkVec_tokenCheck_counter_23 + sinkVec_tokenCheck_counterChange_23;
      if (sinkVec_shifterValid_23) begin
        sinkVec_shifterReg_23_0_valid <= sinkVec_validSource_23_valid;
        sinkVec_shifterReg_23_0_bits_vd <= sinkVec_validSource_23_bits_vd;
        sinkVec_shifterReg_23_0_bits_offset <= sinkVec_validSource_23_bits_offset;
        sinkVec_shifterReg_23_0_bits_mask <= sinkVec_validSource_23_bits_mask;
        sinkVec_shifterReg_23_0_bits_data <= sinkVec_validSource_23_bits_data;
        sinkVec_shifterReg_23_0_bits_last <= sinkVec_validSource_23_bits_last;
        sinkVec_shifterReg_23_0_bits_instructionIndex <= sinkVec_validSource_23_bits_instructionIndex;
      end
      maskUnitFirst_11 <= tryToRead_11 & ~(sinkWire_11_ready & sinkWire_11_valid) ^ maskUnitFirst_11;
      view__writeRelease_5_pipe_v <= sinkVec_11_0_ready & sinkVec_11_0_valid;
      pipe_v_15 <= sinkVec_11_1_ready & sinkVec_11_1_valid;
      instructionFinishedPipe_pipe_v_5 <= 1'h1;
      pipe_v_16 <= 1'h1;
      pipe_pipe_v_5 <= pipe_v_16;
      view__laneMaskSelect_5_pipe_v <= 1'h1;
      view__laneMaskSelect_5_pipe_pipe_v <= view__laneMaskSelect_5_pipe_v;
      view__laneMaskSewSelect_5_pipe_v <= 1'h1;
      view__laneMaskSewSelect_5_pipe_pipe_v <= view__laneMaskSewSelect_5_pipe_v;
      lsuLastPipe_pipe_v_5 <= 1'h1;
      maskLastPipe_pipe_v_5 <= 1'h1;
      pipe_v_17 <= 1'h1;
      sinkVec_releasePipe_pipe_v_24 <= sinkVec_sinkWire_24_ready & sinkVec_sinkWire_24_valid;
      if (sinkVec_validSource_24_valid ^ sinkVec_releasePipe_pipe_out_24_valid)
        sinkVec_tokenCheck_counter_24 <= sinkVec_tokenCheck_counter_24 + sinkVec_tokenCheck_counterChange_24;
      if (sinkVec_shifterValid_24) begin
        sinkVec_shifterReg_24_0_valid <= sinkVec_validSource_24_valid;
        sinkVec_shifterReg_24_0_bits_vs <= sinkVec_validSource_24_bits_vs;
        sinkVec_shifterReg_24_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_24_0_bits_offset <= sinkVec_validSource_24_bits_offset;
        sinkVec_shifterReg_24_0_bits_instructionIndex <= sinkVec_validSource_24_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_25 <= sinkVec_sinkWire_25_ready & sinkVec_sinkWire_25_valid;
      if (sinkVec_validSource_25_valid ^ sinkVec_releasePipe_pipe_out_25_valid)
        sinkVec_tokenCheck_counter_25 <= sinkVec_tokenCheck_counter_25 + sinkVec_tokenCheck_counterChange_25;
      if (sinkVec_shifterValid_25) begin
        sinkVec_shifterReg_25_0_valid <= sinkVec_validSource_25_valid;
        sinkVec_shifterReg_25_0_bits_vs <= sinkVec_validSource_25_bits_vs;
        sinkVec_shifterReg_25_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_25_0_bits_offset <= sinkVec_validSource_25_bits_offset;
        sinkVec_shifterReg_25_0_bits_instructionIndex <= sinkVec_validSource_25_bits_instructionIndex;
      end
      maskUnitFirst_12 <= tryToRead_12 & ~(sinkWire_12_ready & sinkWire_12_valid) ^ maskUnitFirst_12;
      accessDataValid_pipe_v_12 <= sinkVec_12_0_ready & sinkVec_12_0_valid;
      accessDataValid_pipe_pipe_v_12 <= accessDataValid_pipe_v_12;
      if (shifterValid_28) begin
        shifterReg_28_0_valid <= accessDataSource_12_valid;
        shifterReg_28_0_bits <= accessDataSource_12_bits;
      end
      accessDataValid_pipe_v_13 <= sinkVec_12_1_ready & sinkVec_12_1_valid;
      accessDataValid_pipe_pipe_v_13 <= accessDataValid_pipe_v_13;
      if (shifterValid_29) begin
        shifterReg_29_0_valid <= accessDataSource_13_valid;
        shifterReg_29_0_bits <= accessDataSource_13_bits;
      end
      sinkVec_releasePipe_pipe_v_26 <= sinkVec_sinkWire_26_ready & sinkVec_sinkWire_26_valid;
      if (sinkVec_validSource_26_valid ^ sinkVec_releasePipe_pipe_out_26_valid)
        sinkVec_tokenCheck_counter_26 <= sinkVec_tokenCheck_counter_26 + sinkVec_tokenCheck_counterChange_26;
      if (sinkVec_shifterValid_26) begin
        sinkVec_shifterReg_26_0_valid <= sinkVec_validSource_26_valid;
        sinkVec_shifterReg_26_0_bits_vd <= sinkVec_validSource_26_bits_vd;
        sinkVec_shifterReg_26_0_bits_offset <= sinkVec_validSource_26_bits_offset;
        sinkVec_shifterReg_26_0_bits_mask <= sinkVec_validSource_26_bits_mask;
        sinkVec_shifterReg_26_0_bits_data <= sinkVec_validSource_26_bits_data;
        sinkVec_shifterReg_26_0_bits_instructionIndex <= sinkVec_validSource_26_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_27 <= sinkVec_sinkWire_27_ready & sinkVec_sinkWire_27_valid;
      if (sinkVec_validSource_27_valid ^ sinkVec_releasePipe_pipe_out_27_valid)
        sinkVec_tokenCheck_counter_27 <= sinkVec_tokenCheck_counter_27 + sinkVec_tokenCheck_counterChange_27;
      if (sinkVec_shifterValid_27) begin
        sinkVec_shifterReg_27_0_valid <= sinkVec_validSource_27_valid;
        sinkVec_shifterReg_27_0_bits_vd <= sinkVec_validSource_27_bits_vd;
        sinkVec_shifterReg_27_0_bits_offset <= sinkVec_validSource_27_bits_offset;
        sinkVec_shifterReg_27_0_bits_mask <= sinkVec_validSource_27_bits_mask;
        sinkVec_shifterReg_27_0_bits_data <= sinkVec_validSource_27_bits_data;
        sinkVec_shifterReg_27_0_bits_last <= sinkVec_validSource_27_bits_last;
        sinkVec_shifterReg_27_0_bits_instructionIndex <= sinkVec_validSource_27_bits_instructionIndex;
      end
      maskUnitFirst_13 <= tryToRead_13 & ~(sinkWire_13_ready & sinkWire_13_valid) ^ maskUnitFirst_13;
      view__writeRelease_6_pipe_v <= sinkVec_13_0_ready & sinkVec_13_0_valid;
      pipe_v_18 <= sinkVec_13_1_ready & sinkVec_13_1_valid;
      instructionFinishedPipe_pipe_v_6 <= 1'h1;
      pipe_v_19 <= 1'h1;
      pipe_pipe_v_6 <= pipe_v_19;
      view__laneMaskSelect_6_pipe_v <= 1'h1;
      view__laneMaskSelect_6_pipe_pipe_v <= view__laneMaskSelect_6_pipe_v;
      view__laneMaskSewSelect_6_pipe_v <= 1'h1;
      view__laneMaskSewSelect_6_pipe_pipe_v <= view__laneMaskSewSelect_6_pipe_v;
      lsuLastPipe_pipe_v_6 <= 1'h1;
      maskLastPipe_pipe_v_6 <= 1'h1;
      pipe_v_20 <= 1'h1;
      sinkVec_releasePipe_pipe_v_28 <= sinkVec_sinkWire_28_ready & sinkVec_sinkWire_28_valid;
      if (sinkVec_validSource_28_valid ^ sinkVec_releasePipe_pipe_out_28_valid)
        sinkVec_tokenCheck_counter_28 <= sinkVec_tokenCheck_counter_28 + sinkVec_tokenCheck_counterChange_28;
      if (sinkVec_shifterValid_28) begin
        sinkVec_shifterReg_28_0_valid <= sinkVec_validSource_28_valid;
        sinkVec_shifterReg_28_0_bits_vs <= sinkVec_validSource_28_bits_vs;
        sinkVec_shifterReg_28_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_28_0_bits_offset <= sinkVec_validSource_28_bits_offset;
        sinkVec_shifterReg_28_0_bits_instructionIndex <= sinkVec_validSource_28_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_29 <= sinkVec_sinkWire_29_ready & sinkVec_sinkWire_29_valid;
      if (sinkVec_validSource_29_valid ^ sinkVec_releasePipe_pipe_out_29_valid)
        sinkVec_tokenCheck_counter_29 <= sinkVec_tokenCheck_counter_29 + sinkVec_tokenCheck_counterChange_29;
      if (sinkVec_shifterValid_29) begin
        sinkVec_shifterReg_29_0_valid <= sinkVec_validSource_29_valid;
        sinkVec_shifterReg_29_0_bits_vs <= sinkVec_validSource_29_bits_vs;
        sinkVec_shifterReg_29_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_29_0_bits_offset <= sinkVec_validSource_29_bits_offset;
        sinkVec_shifterReg_29_0_bits_instructionIndex <= sinkVec_validSource_29_bits_instructionIndex;
      end
      maskUnitFirst_14 <= tryToRead_14 & ~(sinkWire_14_ready & sinkWire_14_valid) ^ maskUnitFirst_14;
      accessDataValid_pipe_v_14 <= sinkVec_14_0_ready & sinkVec_14_0_valid;
      accessDataValid_pipe_pipe_v_14 <= accessDataValid_pipe_v_14;
      if (shifterValid_30) begin
        shifterReg_30_0_valid <= accessDataSource_14_valid;
        shifterReg_30_0_bits <= accessDataSource_14_bits;
      end
      accessDataValid_pipe_v_15 <= sinkVec_14_1_ready & sinkVec_14_1_valid;
      accessDataValid_pipe_pipe_v_15 <= accessDataValid_pipe_v_15;
      if (shifterValid_31) begin
        shifterReg_31_0_valid <= accessDataSource_15_valid;
        shifterReg_31_0_bits <= accessDataSource_15_bits;
      end
      sinkVec_releasePipe_pipe_v_30 <= sinkVec_sinkWire_30_ready & sinkVec_sinkWire_30_valid;
      if (sinkVec_validSource_30_valid ^ sinkVec_releasePipe_pipe_out_30_valid)
        sinkVec_tokenCheck_counter_30 <= sinkVec_tokenCheck_counter_30 + sinkVec_tokenCheck_counterChange_30;
      if (sinkVec_shifterValid_30) begin
        sinkVec_shifterReg_30_0_valid <= sinkVec_validSource_30_valid;
        sinkVec_shifterReg_30_0_bits_vd <= sinkVec_validSource_30_bits_vd;
        sinkVec_shifterReg_30_0_bits_offset <= sinkVec_validSource_30_bits_offset;
        sinkVec_shifterReg_30_0_bits_mask <= sinkVec_validSource_30_bits_mask;
        sinkVec_shifterReg_30_0_bits_data <= sinkVec_validSource_30_bits_data;
        sinkVec_shifterReg_30_0_bits_instructionIndex <= sinkVec_validSource_30_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_31 <= sinkVec_sinkWire_31_ready & sinkVec_sinkWire_31_valid;
      if (sinkVec_validSource_31_valid ^ sinkVec_releasePipe_pipe_out_31_valid)
        sinkVec_tokenCheck_counter_31 <= sinkVec_tokenCheck_counter_31 + sinkVec_tokenCheck_counterChange_31;
      if (sinkVec_shifterValid_31) begin
        sinkVec_shifterReg_31_0_valid <= sinkVec_validSource_31_valid;
        sinkVec_shifterReg_31_0_bits_vd <= sinkVec_validSource_31_bits_vd;
        sinkVec_shifterReg_31_0_bits_offset <= sinkVec_validSource_31_bits_offset;
        sinkVec_shifterReg_31_0_bits_mask <= sinkVec_validSource_31_bits_mask;
        sinkVec_shifterReg_31_0_bits_data <= sinkVec_validSource_31_bits_data;
        sinkVec_shifterReg_31_0_bits_last <= sinkVec_validSource_31_bits_last;
        sinkVec_shifterReg_31_0_bits_instructionIndex <= sinkVec_validSource_31_bits_instructionIndex;
      end
      maskUnitFirst_15 <= tryToRead_15 & ~(sinkWire_15_ready & sinkWire_15_valid) ^ maskUnitFirst_15;
      view__writeRelease_7_pipe_v <= sinkVec_15_0_ready & sinkVec_15_0_valid;
      pipe_v_21 <= sinkVec_15_1_ready & sinkVec_15_1_valid;
      instructionFinishedPipe_pipe_v_7 <= 1'h1;
      pipe_v_22 <= 1'h1;
      pipe_pipe_v_7 <= pipe_v_22;
      view__laneMaskSelect_7_pipe_v <= 1'h1;
      view__laneMaskSelect_7_pipe_pipe_v <= view__laneMaskSelect_7_pipe_v;
      view__laneMaskSewSelect_7_pipe_v <= 1'h1;
      view__laneMaskSewSelect_7_pipe_pipe_v <= view__laneMaskSewSelect_7_pipe_v;
      lsuLastPipe_pipe_v_7 <= 1'h1;
      maskLastPipe_pipe_v_7 <= 1'h1;
      pipe_v_23 <= 1'h1;
      sinkVec_releasePipe_pipe_v_32 <= sinkVec_sinkWire_32_ready & sinkVec_sinkWire_32_valid;
      if (sinkVec_validSource_32_valid ^ sinkVec_releasePipe_pipe_out_32_valid)
        sinkVec_tokenCheck_counter_32 <= sinkVec_tokenCheck_counter_32 + sinkVec_tokenCheck_counterChange_32;
      if (sinkVec_shifterValid_32) begin
        sinkVec_shifterReg_32_0_valid <= sinkVec_validSource_32_valid;
        sinkVec_shifterReg_32_0_bits_vs <= sinkVec_validSource_32_bits_vs;
        sinkVec_shifterReg_32_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_32_0_bits_offset <= sinkVec_validSource_32_bits_offset;
        sinkVec_shifterReg_32_0_bits_instructionIndex <= sinkVec_validSource_32_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_33 <= sinkVec_sinkWire_33_ready & sinkVec_sinkWire_33_valid;
      if (sinkVec_validSource_33_valid ^ sinkVec_releasePipe_pipe_out_33_valid)
        sinkVec_tokenCheck_counter_33 <= sinkVec_tokenCheck_counter_33 + sinkVec_tokenCheck_counterChange_33;
      if (sinkVec_shifterValid_33) begin
        sinkVec_shifterReg_33_0_valid <= sinkVec_validSource_33_valid;
        sinkVec_shifterReg_33_0_bits_vs <= sinkVec_validSource_33_bits_vs;
        sinkVec_shifterReg_33_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_33_0_bits_offset <= sinkVec_validSource_33_bits_offset;
        sinkVec_shifterReg_33_0_bits_instructionIndex <= sinkVec_validSource_33_bits_instructionIndex;
      end
      maskUnitFirst_16 <= tryToRead_16 & ~(sinkWire_16_ready & sinkWire_16_valid) ^ maskUnitFirst_16;
      accessDataValid_pipe_v_16 <= sinkVec_16_0_ready & sinkVec_16_0_valid;
      accessDataValid_pipe_pipe_v_16 <= accessDataValid_pipe_v_16;
      if (shifterValid_32) begin
        shifterReg_32_0_valid <= accessDataSource_16_valid;
        shifterReg_32_0_bits <= accessDataSource_16_bits;
      end
      accessDataValid_pipe_v_17 <= sinkVec_16_1_ready & sinkVec_16_1_valid;
      accessDataValid_pipe_pipe_v_17 <= accessDataValid_pipe_v_17;
      if (shifterValid_33) begin
        shifterReg_33_0_valid <= accessDataSource_17_valid;
        shifterReg_33_0_bits <= accessDataSource_17_bits;
      end
      sinkVec_releasePipe_pipe_v_34 <= sinkVec_sinkWire_34_ready & sinkVec_sinkWire_34_valid;
      if (sinkVec_validSource_34_valid ^ sinkVec_releasePipe_pipe_out_34_valid)
        sinkVec_tokenCheck_counter_34 <= sinkVec_tokenCheck_counter_34 + sinkVec_tokenCheck_counterChange_34;
      if (sinkVec_shifterValid_34) begin
        sinkVec_shifterReg_34_0_valid <= sinkVec_validSource_34_valid;
        sinkVec_shifterReg_34_0_bits_vd <= sinkVec_validSource_34_bits_vd;
        sinkVec_shifterReg_34_0_bits_offset <= sinkVec_validSource_34_bits_offset;
        sinkVec_shifterReg_34_0_bits_mask <= sinkVec_validSource_34_bits_mask;
        sinkVec_shifterReg_34_0_bits_data <= sinkVec_validSource_34_bits_data;
        sinkVec_shifterReg_34_0_bits_instructionIndex <= sinkVec_validSource_34_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_35 <= sinkVec_sinkWire_35_ready & sinkVec_sinkWire_35_valid;
      if (sinkVec_validSource_35_valid ^ sinkVec_releasePipe_pipe_out_35_valid)
        sinkVec_tokenCheck_counter_35 <= sinkVec_tokenCheck_counter_35 + sinkVec_tokenCheck_counterChange_35;
      if (sinkVec_shifterValid_35) begin
        sinkVec_shifterReg_35_0_valid <= sinkVec_validSource_35_valid;
        sinkVec_shifterReg_35_0_bits_vd <= sinkVec_validSource_35_bits_vd;
        sinkVec_shifterReg_35_0_bits_offset <= sinkVec_validSource_35_bits_offset;
        sinkVec_shifterReg_35_0_bits_mask <= sinkVec_validSource_35_bits_mask;
        sinkVec_shifterReg_35_0_bits_data <= sinkVec_validSource_35_bits_data;
        sinkVec_shifterReg_35_0_bits_last <= sinkVec_validSource_35_bits_last;
        sinkVec_shifterReg_35_0_bits_instructionIndex <= sinkVec_validSource_35_bits_instructionIndex;
      end
      maskUnitFirst_17 <= tryToRead_17 & ~(sinkWire_17_ready & sinkWire_17_valid) ^ maskUnitFirst_17;
      view__writeRelease_8_pipe_v <= sinkVec_17_0_ready & sinkVec_17_0_valid;
      pipe_v_24 <= sinkVec_17_1_ready & sinkVec_17_1_valid;
      instructionFinishedPipe_pipe_v_8 <= 1'h1;
      pipe_v_25 <= 1'h1;
      pipe_pipe_v_8 <= pipe_v_25;
      view__laneMaskSelect_8_pipe_v <= 1'h1;
      view__laneMaskSelect_8_pipe_pipe_v <= view__laneMaskSelect_8_pipe_v;
      view__laneMaskSewSelect_8_pipe_v <= 1'h1;
      view__laneMaskSewSelect_8_pipe_pipe_v <= view__laneMaskSewSelect_8_pipe_v;
      lsuLastPipe_pipe_v_8 <= 1'h1;
      maskLastPipe_pipe_v_8 <= 1'h1;
      pipe_v_26 <= 1'h1;
      sinkVec_releasePipe_pipe_v_36 <= sinkVec_sinkWire_36_ready & sinkVec_sinkWire_36_valid;
      if (sinkVec_validSource_36_valid ^ sinkVec_releasePipe_pipe_out_36_valid)
        sinkVec_tokenCheck_counter_36 <= sinkVec_tokenCheck_counter_36 + sinkVec_tokenCheck_counterChange_36;
      if (sinkVec_shifterValid_36) begin
        sinkVec_shifterReg_36_0_valid <= sinkVec_validSource_36_valid;
        sinkVec_shifterReg_36_0_bits_vs <= sinkVec_validSource_36_bits_vs;
        sinkVec_shifterReg_36_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_36_0_bits_offset <= sinkVec_validSource_36_bits_offset;
        sinkVec_shifterReg_36_0_bits_instructionIndex <= sinkVec_validSource_36_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_37 <= sinkVec_sinkWire_37_ready & sinkVec_sinkWire_37_valid;
      if (sinkVec_validSource_37_valid ^ sinkVec_releasePipe_pipe_out_37_valid)
        sinkVec_tokenCheck_counter_37 <= sinkVec_tokenCheck_counter_37 + sinkVec_tokenCheck_counterChange_37;
      if (sinkVec_shifterValid_37) begin
        sinkVec_shifterReg_37_0_valid <= sinkVec_validSource_37_valid;
        sinkVec_shifterReg_37_0_bits_vs <= sinkVec_validSource_37_bits_vs;
        sinkVec_shifterReg_37_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_37_0_bits_offset <= sinkVec_validSource_37_bits_offset;
        sinkVec_shifterReg_37_0_bits_instructionIndex <= sinkVec_validSource_37_bits_instructionIndex;
      end
      maskUnitFirst_18 <= tryToRead_18 & ~(sinkWire_18_ready & sinkWire_18_valid) ^ maskUnitFirst_18;
      accessDataValid_pipe_v_18 <= sinkVec_18_0_ready & sinkVec_18_0_valid;
      accessDataValid_pipe_pipe_v_18 <= accessDataValid_pipe_v_18;
      if (shifterValid_34) begin
        shifterReg_34_0_valid <= accessDataSource_18_valid;
        shifterReg_34_0_bits <= accessDataSource_18_bits;
      end
      accessDataValid_pipe_v_19 <= sinkVec_18_1_ready & sinkVec_18_1_valid;
      accessDataValid_pipe_pipe_v_19 <= accessDataValid_pipe_v_19;
      if (shifterValid_35) begin
        shifterReg_35_0_valid <= accessDataSource_19_valid;
        shifterReg_35_0_bits <= accessDataSource_19_bits;
      end
      sinkVec_releasePipe_pipe_v_38 <= sinkVec_sinkWire_38_ready & sinkVec_sinkWire_38_valid;
      if (sinkVec_validSource_38_valid ^ sinkVec_releasePipe_pipe_out_38_valid)
        sinkVec_tokenCheck_counter_38 <= sinkVec_tokenCheck_counter_38 + sinkVec_tokenCheck_counterChange_38;
      if (sinkVec_shifterValid_38) begin
        sinkVec_shifterReg_38_0_valid <= sinkVec_validSource_38_valid;
        sinkVec_shifterReg_38_0_bits_vd <= sinkVec_validSource_38_bits_vd;
        sinkVec_shifterReg_38_0_bits_offset <= sinkVec_validSource_38_bits_offset;
        sinkVec_shifterReg_38_0_bits_mask <= sinkVec_validSource_38_bits_mask;
        sinkVec_shifterReg_38_0_bits_data <= sinkVec_validSource_38_bits_data;
        sinkVec_shifterReg_38_0_bits_instructionIndex <= sinkVec_validSource_38_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_39 <= sinkVec_sinkWire_39_ready & sinkVec_sinkWire_39_valid;
      if (sinkVec_validSource_39_valid ^ sinkVec_releasePipe_pipe_out_39_valid)
        sinkVec_tokenCheck_counter_39 <= sinkVec_tokenCheck_counter_39 + sinkVec_tokenCheck_counterChange_39;
      if (sinkVec_shifterValid_39) begin
        sinkVec_shifterReg_39_0_valid <= sinkVec_validSource_39_valid;
        sinkVec_shifterReg_39_0_bits_vd <= sinkVec_validSource_39_bits_vd;
        sinkVec_shifterReg_39_0_bits_offset <= sinkVec_validSource_39_bits_offset;
        sinkVec_shifterReg_39_0_bits_mask <= sinkVec_validSource_39_bits_mask;
        sinkVec_shifterReg_39_0_bits_data <= sinkVec_validSource_39_bits_data;
        sinkVec_shifterReg_39_0_bits_last <= sinkVec_validSource_39_bits_last;
        sinkVec_shifterReg_39_0_bits_instructionIndex <= sinkVec_validSource_39_bits_instructionIndex;
      end
      maskUnitFirst_19 <= tryToRead_19 & ~(sinkWire_19_ready & sinkWire_19_valid) ^ maskUnitFirst_19;
      view__writeRelease_9_pipe_v <= sinkVec_19_0_ready & sinkVec_19_0_valid;
      pipe_v_27 <= sinkVec_19_1_ready & sinkVec_19_1_valid;
      instructionFinishedPipe_pipe_v_9 <= 1'h1;
      pipe_v_28 <= 1'h1;
      pipe_pipe_v_9 <= pipe_v_28;
      view__laneMaskSelect_9_pipe_v <= 1'h1;
      view__laneMaskSelect_9_pipe_pipe_v <= view__laneMaskSelect_9_pipe_v;
      view__laneMaskSewSelect_9_pipe_v <= 1'h1;
      view__laneMaskSewSelect_9_pipe_pipe_v <= view__laneMaskSewSelect_9_pipe_v;
      lsuLastPipe_pipe_v_9 <= 1'h1;
      maskLastPipe_pipe_v_9 <= 1'h1;
      pipe_v_29 <= 1'h1;
      sinkVec_releasePipe_pipe_v_40 <= sinkVec_sinkWire_40_ready & sinkVec_sinkWire_40_valid;
      if (sinkVec_validSource_40_valid ^ sinkVec_releasePipe_pipe_out_40_valid)
        sinkVec_tokenCheck_counter_40 <= sinkVec_tokenCheck_counter_40 + sinkVec_tokenCheck_counterChange_40;
      if (sinkVec_shifterValid_40) begin
        sinkVec_shifterReg_40_0_valid <= sinkVec_validSource_40_valid;
        sinkVec_shifterReg_40_0_bits_vs <= sinkVec_validSource_40_bits_vs;
        sinkVec_shifterReg_40_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_40_0_bits_offset <= sinkVec_validSource_40_bits_offset;
        sinkVec_shifterReg_40_0_bits_instructionIndex <= sinkVec_validSource_40_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_41 <= sinkVec_sinkWire_41_ready & sinkVec_sinkWire_41_valid;
      if (sinkVec_validSource_41_valid ^ sinkVec_releasePipe_pipe_out_41_valid)
        sinkVec_tokenCheck_counter_41 <= sinkVec_tokenCheck_counter_41 + sinkVec_tokenCheck_counterChange_41;
      if (sinkVec_shifterValid_41) begin
        sinkVec_shifterReg_41_0_valid <= sinkVec_validSource_41_valid;
        sinkVec_shifterReg_41_0_bits_vs <= sinkVec_validSource_41_bits_vs;
        sinkVec_shifterReg_41_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_41_0_bits_offset <= sinkVec_validSource_41_bits_offset;
        sinkVec_shifterReg_41_0_bits_instructionIndex <= sinkVec_validSource_41_bits_instructionIndex;
      end
      maskUnitFirst_20 <= tryToRead_20 & ~(sinkWire_20_ready & sinkWire_20_valid) ^ maskUnitFirst_20;
      accessDataValid_pipe_v_20 <= sinkVec_20_0_ready & sinkVec_20_0_valid;
      accessDataValid_pipe_pipe_v_20 <= accessDataValid_pipe_v_20;
      if (shifterValid_36) begin
        shifterReg_36_0_valid <= accessDataSource_20_valid;
        shifterReg_36_0_bits <= accessDataSource_20_bits;
      end
      accessDataValid_pipe_v_21 <= sinkVec_20_1_ready & sinkVec_20_1_valid;
      accessDataValid_pipe_pipe_v_21 <= accessDataValid_pipe_v_21;
      if (shifterValid_37) begin
        shifterReg_37_0_valid <= accessDataSource_21_valid;
        shifterReg_37_0_bits <= accessDataSource_21_bits;
      end
      sinkVec_releasePipe_pipe_v_42 <= sinkVec_sinkWire_42_ready & sinkVec_sinkWire_42_valid;
      if (sinkVec_validSource_42_valid ^ sinkVec_releasePipe_pipe_out_42_valid)
        sinkVec_tokenCheck_counter_42 <= sinkVec_tokenCheck_counter_42 + sinkVec_tokenCheck_counterChange_42;
      if (sinkVec_shifterValid_42) begin
        sinkVec_shifterReg_42_0_valid <= sinkVec_validSource_42_valid;
        sinkVec_shifterReg_42_0_bits_vd <= sinkVec_validSource_42_bits_vd;
        sinkVec_shifterReg_42_0_bits_offset <= sinkVec_validSource_42_bits_offset;
        sinkVec_shifterReg_42_0_bits_mask <= sinkVec_validSource_42_bits_mask;
        sinkVec_shifterReg_42_0_bits_data <= sinkVec_validSource_42_bits_data;
        sinkVec_shifterReg_42_0_bits_instructionIndex <= sinkVec_validSource_42_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_43 <= sinkVec_sinkWire_43_ready & sinkVec_sinkWire_43_valid;
      if (sinkVec_validSource_43_valid ^ sinkVec_releasePipe_pipe_out_43_valid)
        sinkVec_tokenCheck_counter_43 <= sinkVec_tokenCheck_counter_43 + sinkVec_tokenCheck_counterChange_43;
      if (sinkVec_shifterValid_43) begin
        sinkVec_shifterReg_43_0_valid <= sinkVec_validSource_43_valid;
        sinkVec_shifterReg_43_0_bits_vd <= sinkVec_validSource_43_bits_vd;
        sinkVec_shifterReg_43_0_bits_offset <= sinkVec_validSource_43_bits_offset;
        sinkVec_shifterReg_43_0_bits_mask <= sinkVec_validSource_43_bits_mask;
        sinkVec_shifterReg_43_0_bits_data <= sinkVec_validSource_43_bits_data;
        sinkVec_shifterReg_43_0_bits_last <= sinkVec_validSource_43_bits_last;
        sinkVec_shifterReg_43_0_bits_instructionIndex <= sinkVec_validSource_43_bits_instructionIndex;
      end
      maskUnitFirst_21 <= tryToRead_21 & ~(sinkWire_21_ready & sinkWire_21_valid) ^ maskUnitFirst_21;
      view__writeRelease_10_pipe_v <= sinkVec_21_0_ready & sinkVec_21_0_valid;
      pipe_v_30 <= sinkVec_21_1_ready & sinkVec_21_1_valid;
      instructionFinishedPipe_pipe_v_10 <= 1'h1;
      pipe_v_31 <= 1'h1;
      pipe_pipe_v_10 <= pipe_v_31;
      view__laneMaskSelect_10_pipe_v <= 1'h1;
      view__laneMaskSelect_10_pipe_pipe_v <= view__laneMaskSelect_10_pipe_v;
      view__laneMaskSewSelect_10_pipe_v <= 1'h1;
      view__laneMaskSewSelect_10_pipe_pipe_v <= view__laneMaskSewSelect_10_pipe_v;
      lsuLastPipe_pipe_v_10 <= 1'h1;
      maskLastPipe_pipe_v_10 <= 1'h1;
      pipe_v_32 <= 1'h1;
      sinkVec_releasePipe_pipe_v_44 <= sinkVec_sinkWire_44_ready & sinkVec_sinkWire_44_valid;
      if (sinkVec_validSource_44_valid ^ sinkVec_releasePipe_pipe_out_44_valid)
        sinkVec_tokenCheck_counter_44 <= sinkVec_tokenCheck_counter_44 + sinkVec_tokenCheck_counterChange_44;
      if (sinkVec_shifterValid_44) begin
        sinkVec_shifterReg_44_0_valid <= sinkVec_validSource_44_valid;
        sinkVec_shifterReg_44_0_bits_vs <= sinkVec_validSource_44_bits_vs;
        sinkVec_shifterReg_44_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_44_0_bits_offset <= sinkVec_validSource_44_bits_offset;
        sinkVec_shifterReg_44_0_bits_instructionIndex <= sinkVec_validSource_44_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_45 <= sinkVec_sinkWire_45_ready & sinkVec_sinkWire_45_valid;
      if (sinkVec_validSource_45_valid ^ sinkVec_releasePipe_pipe_out_45_valid)
        sinkVec_tokenCheck_counter_45 <= sinkVec_tokenCheck_counter_45 + sinkVec_tokenCheck_counterChange_45;
      if (sinkVec_shifterValid_45) begin
        sinkVec_shifterReg_45_0_valid <= sinkVec_validSource_45_valid;
        sinkVec_shifterReg_45_0_bits_vs <= sinkVec_validSource_45_bits_vs;
        sinkVec_shifterReg_45_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_45_0_bits_offset <= sinkVec_validSource_45_bits_offset;
        sinkVec_shifterReg_45_0_bits_instructionIndex <= sinkVec_validSource_45_bits_instructionIndex;
      end
      maskUnitFirst_22 <= tryToRead_22 & ~(sinkWire_22_ready & sinkWire_22_valid) ^ maskUnitFirst_22;
      accessDataValid_pipe_v_22 <= sinkVec_22_0_ready & sinkVec_22_0_valid;
      accessDataValid_pipe_pipe_v_22 <= accessDataValid_pipe_v_22;
      if (shifterValid_38) begin
        shifterReg_38_0_valid <= accessDataSource_22_valid;
        shifterReg_38_0_bits <= accessDataSource_22_bits;
      end
      accessDataValid_pipe_v_23 <= sinkVec_22_1_ready & sinkVec_22_1_valid;
      accessDataValid_pipe_pipe_v_23 <= accessDataValid_pipe_v_23;
      if (shifterValid_39) begin
        shifterReg_39_0_valid <= accessDataSource_23_valid;
        shifterReg_39_0_bits <= accessDataSource_23_bits;
      end
      sinkVec_releasePipe_pipe_v_46 <= sinkVec_sinkWire_46_ready & sinkVec_sinkWire_46_valid;
      if (sinkVec_validSource_46_valid ^ sinkVec_releasePipe_pipe_out_46_valid)
        sinkVec_tokenCheck_counter_46 <= sinkVec_tokenCheck_counter_46 + sinkVec_tokenCheck_counterChange_46;
      if (sinkVec_shifterValid_46) begin
        sinkVec_shifterReg_46_0_valid <= sinkVec_validSource_46_valid;
        sinkVec_shifterReg_46_0_bits_vd <= sinkVec_validSource_46_bits_vd;
        sinkVec_shifterReg_46_0_bits_offset <= sinkVec_validSource_46_bits_offset;
        sinkVec_shifterReg_46_0_bits_mask <= sinkVec_validSource_46_bits_mask;
        sinkVec_shifterReg_46_0_bits_data <= sinkVec_validSource_46_bits_data;
        sinkVec_shifterReg_46_0_bits_instructionIndex <= sinkVec_validSource_46_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_47 <= sinkVec_sinkWire_47_ready & sinkVec_sinkWire_47_valid;
      if (sinkVec_validSource_47_valid ^ sinkVec_releasePipe_pipe_out_47_valid)
        sinkVec_tokenCheck_counter_47 <= sinkVec_tokenCheck_counter_47 + sinkVec_tokenCheck_counterChange_47;
      if (sinkVec_shifterValid_47) begin
        sinkVec_shifterReg_47_0_valid <= sinkVec_validSource_47_valid;
        sinkVec_shifterReg_47_0_bits_vd <= sinkVec_validSource_47_bits_vd;
        sinkVec_shifterReg_47_0_bits_offset <= sinkVec_validSource_47_bits_offset;
        sinkVec_shifterReg_47_0_bits_mask <= sinkVec_validSource_47_bits_mask;
        sinkVec_shifterReg_47_0_bits_data <= sinkVec_validSource_47_bits_data;
        sinkVec_shifterReg_47_0_bits_last <= sinkVec_validSource_47_bits_last;
        sinkVec_shifterReg_47_0_bits_instructionIndex <= sinkVec_validSource_47_bits_instructionIndex;
      end
      maskUnitFirst_23 <= tryToRead_23 & ~(sinkWire_23_ready & sinkWire_23_valid) ^ maskUnitFirst_23;
      view__writeRelease_11_pipe_v <= sinkVec_23_0_ready & sinkVec_23_0_valid;
      pipe_v_33 <= sinkVec_23_1_ready & sinkVec_23_1_valid;
      instructionFinishedPipe_pipe_v_11 <= 1'h1;
      pipe_v_34 <= 1'h1;
      pipe_pipe_v_11 <= pipe_v_34;
      view__laneMaskSelect_11_pipe_v <= 1'h1;
      view__laneMaskSelect_11_pipe_pipe_v <= view__laneMaskSelect_11_pipe_v;
      view__laneMaskSewSelect_11_pipe_v <= 1'h1;
      view__laneMaskSewSelect_11_pipe_pipe_v <= view__laneMaskSewSelect_11_pipe_v;
      lsuLastPipe_pipe_v_11 <= 1'h1;
      maskLastPipe_pipe_v_11 <= 1'h1;
      pipe_v_35 <= 1'h1;
      sinkVec_releasePipe_pipe_v_48 <= sinkVec_sinkWire_48_ready & sinkVec_sinkWire_48_valid;
      if (sinkVec_validSource_48_valid ^ sinkVec_releasePipe_pipe_out_48_valid)
        sinkVec_tokenCheck_counter_48 <= sinkVec_tokenCheck_counter_48 + sinkVec_tokenCheck_counterChange_48;
      if (sinkVec_shifterValid_48) begin
        sinkVec_shifterReg_48_0_valid <= sinkVec_validSource_48_valid;
        sinkVec_shifterReg_48_0_bits_vs <= sinkVec_validSource_48_bits_vs;
        sinkVec_shifterReg_48_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_48_0_bits_offset <= sinkVec_validSource_48_bits_offset;
        sinkVec_shifterReg_48_0_bits_instructionIndex <= sinkVec_validSource_48_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_49 <= sinkVec_sinkWire_49_ready & sinkVec_sinkWire_49_valid;
      if (sinkVec_validSource_49_valid ^ sinkVec_releasePipe_pipe_out_49_valid)
        sinkVec_tokenCheck_counter_49 <= sinkVec_tokenCheck_counter_49 + sinkVec_tokenCheck_counterChange_49;
      if (sinkVec_shifterValid_49) begin
        sinkVec_shifterReg_49_0_valid <= sinkVec_validSource_49_valid;
        sinkVec_shifterReg_49_0_bits_vs <= sinkVec_validSource_49_bits_vs;
        sinkVec_shifterReg_49_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_49_0_bits_offset <= sinkVec_validSource_49_bits_offset;
        sinkVec_shifterReg_49_0_bits_instructionIndex <= sinkVec_validSource_49_bits_instructionIndex;
      end
      maskUnitFirst_24 <= tryToRead_24 & ~(sinkWire_24_ready & sinkWire_24_valid) ^ maskUnitFirst_24;
      accessDataValid_pipe_v_24 <= sinkVec_24_0_ready & sinkVec_24_0_valid;
      accessDataValid_pipe_pipe_v_24 <= accessDataValid_pipe_v_24;
      if (shifterValid_40) begin
        shifterReg_40_0_valid <= accessDataSource_24_valid;
        shifterReg_40_0_bits <= accessDataSource_24_bits;
      end
      accessDataValid_pipe_v_25 <= sinkVec_24_1_ready & sinkVec_24_1_valid;
      accessDataValid_pipe_pipe_v_25 <= accessDataValid_pipe_v_25;
      if (shifterValid_41) begin
        shifterReg_41_0_valid <= accessDataSource_25_valid;
        shifterReg_41_0_bits <= accessDataSource_25_bits;
      end
      sinkVec_releasePipe_pipe_v_50 <= sinkVec_sinkWire_50_ready & sinkVec_sinkWire_50_valid;
      if (sinkVec_validSource_50_valid ^ sinkVec_releasePipe_pipe_out_50_valid)
        sinkVec_tokenCheck_counter_50 <= sinkVec_tokenCheck_counter_50 + sinkVec_tokenCheck_counterChange_50;
      if (sinkVec_shifterValid_50) begin
        sinkVec_shifterReg_50_0_valid <= sinkVec_validSource_50_valid;
        sinkVec_shifterReg_50_0_bits_vd <= sinkVec_validSource_50_bits_vd;
        sinkVec_shifterReg_50_0_bits_offset <= sinkVec_validSource_50_bits_offset;
        sinkVec_shifterReg_50_0_bits_mask <= sinkVec_validSource_50_bits_mask;
        sinkVec_shifterReg_50_0_bits_data <= sinkVec_validSource_50_bits_data;
        sinkVec_shifterReg_50_0_bits_instructionIndex <= sinkVec_validSource_50_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_51 <= sinkVec_sinkWire_51_ready & sinkVec_sinkWire_51_valid;
      if (sinkVec_validSource_51_valid ^ sinkVec_releasePipe_pipe_out_51_valid)
        sinkVec_tokenCheck_counter_51 <= sinkVec_tokenCheck_counter_51 + sinkVec_tokenCheck_counterChange_51;
      if (sinkVec_shifterValid_51) begin
        sinkVec_shifterReg_51_0_valid <= sinkVec_validSource_51_valid;
        sinkVec_shifterReg_51_0_bits_vd <= sinkVec_validSource_51_bits_vd;
        sinkVec_shifterReg_51_0_bits_offset <= sinkVec_validSource_51_bits_offset;
        sinkVec_shifterReg_51_0_bits_mask <= sinkVec_validSource_51_bits_mask;
        sinkVec_shifterReg_51_0_bits_data <= sinkVec_validSource_51_bits_data;
        sinkVec_shifterReg_51_0_bits_last <= sinkVec_validSource_51_bits_last;
        sinkVec_shifterReg_51_0_bits_instructionIndex <= sinkVec_validSource_51_bits_instructionIndex;
      end
      maskUnitFirst_25 <= tryToRead_25 & ~(sinkWire_25_ready & sinkWire_25_valid) ^ maskUnitFirst_25;
      view__writeRelease_12_pipe_v <= sinkVec_25_0_ready & sinkVec_25_0_valid;
      pipe_v_36 <= sinkVec_25_1_ready & sinkVec_25_1_valid;
      instructionFinishedPipe_pipe_v_12 <= 1'h1;
      pipe_v_37 <= 1'h1;
      pipe_pipe_v_12 <= pipe_v_37;
      view__laneMaskSelect_12_pipe_v <= 1'h1;
      view__laneMaskSelect_12_pipe_pipe_v <= view__laneMaskSelect_12_pipe_v;
      view__laneMaskSewSelect_12_pipe_v <= 1'h1;
      view__laneMaskSewSelect_12_pipe_pipe_v <= view__laneMaskSewSelect_12_pipe_v;
      lsuLastPipe_pipe_v_12 <= 1'h1;
      maskLastPipe_pipe_v_12 <= 1'h1;
      pipe_v_38 <= 1'h1;
      sinkVec_releasePipe_pipe_v_52 <= sinkVec_sinkWire_52_ready & sinkVec_sinkWire_52_valid;
      if (sinkVec_validSource_52_valid ^ sinkVec_releasePipe_pipe_out_52_valid)
        sinkVec_tokenCheck_counter_52 <= sinkVec_tokenCheck_counter_52 + sinkVec_tokenCheck_counterChange_52;
      if (sinkVec_shifterValid_52) begin
        sinkVec_shifterReg_52_0_valid <= sinkVec_validSource_52_valid;
        sinkVec_shifterReg_52_0_bits_vs <= sinkVec_validSource_52_bits_vs;
        sinkVec_shifterReg_52_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_52_0_bits_offset <= sinkVec_validSource_52_bits_offset;
        sinkVec_shifterReg_52_0_bits_instructionIndex <= sinkVec_validSource_52_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_53 <= sinkVec_sinkWire_53_ready & sinkVec_sinkWire_53_valid;
      if (sinkVec_validSource_53_valid ^ sinkVec_releasePipe_pipe_out_53_valid)
        sinkVec_tokenCheck_counter_53 <= sinkVec_tokenCheck_counter_53 + sinkVec_tokenCheck_counterChange_53;
      if (sinkVec_shifterValid_53) begin
        sinkVec_shifterReg_53_0_valid <= sinkVec_validSource_53_valid;
        sinkVec_shifterReg_53_0_bits_vs <= sinkVec_validSource_53_bits_vs;
        sinkVec_shifterReg_53_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_53_0_bits_offset <= sinkVec_validSource_53_bits_offset;
        sinkVec_shifterReg_53_0_bits_instructionIndex <= sinkVec_validSource_53_bits_instructionIndex;
      end
      maskUnitFirst_26 <= tryToRead_26 & ~(sinkWire_26_ready & sinkWire_26_valid) ^ maskUnitFirst_26;
      accessDataValid_pipe_v_26 <= sinkVec_26_0_ready & sinkVec_26_0_valid;
      accessDataValid_pipe_pipe_v_26 <= accessDataValid_pipe_v_26;
      if (shifterValid_42) begin
        shifterReg_42_0_valid <= accessDataSource_26_valid;
        shifterReg_42_0_bits <= accessDataSource_26_bits;
      end
      accessDataValid_pipe_v_27 <= sinkVec_26_1_ready & sinkVec_26_1_valid;
      accessDataValid_pipe_pipe_v_27 <= accessDataValid_pipe_v_27;
      if (shifterValid_43) begin
        shifterReg_43_0_valid <= accessDataSource_27_valid;
        shifterReg_43_0_bits <= accessDataSource_27_bits;
      end
      sinkVec_releasePipe_pipe_v_54 <= sinkVec_sinkWire_54_ready & sinkVec_sinkWire_54_valid;
      if (sinkVec_validSource_54_valid ^ sinkVec_releasePipe_pipe_out_54_valid)
        sinkVec_tokenCheck_counter_54 <= sinkVec_tokenCheck_counter_54 + sinkVec_tokenCheck_counterChange_54;
      if (sinkVec_shifterValid_54) begin
        sinkVec_shifterReg_54_0_valid <= sinkVec_validSource_54_valid;
        sinkVec_shifterReg_54_0_bits_vd <= sinkVec_validSource_54_bits_vd;
        sinkVec_shifterReg_54_0_bits_offset <= sinkVec_validSource_54_bits_offset;
        sinkVec_shifterReg_54_0_bits_mask <= sinkVec_validSource_54_bits_mask;
        sinkVec_shifterReg_54_0_bits_data <= sinkVec_validSource_54_bits_data;
        sinkVec_shifterReg_54_0_bits_instructionIndex <= sinkVec_validSource_54_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_55 <= sinkVec_sinkWire_55_ready & sinkVec_sinkWire_55_valid;
      if (sinkVec_validSource_55_valid ^ sinkVec_releasePipe_pipe_out_55_valid)
        sinkVec_tokenCheck_counter_55 <= sinkVec_tokenCheck_counter_55 + sinkVec_tokenCheck_counterChange_55;
      if (sinkVec_shifterValid_55) begin
        sinkVec_shifterReg_55_0_valid <= sinkVec_validSource_55_valid;
        sinkVec_shifterReg_55_0_bits_vd <= sinkVec_validSource_55_bits_vd;
        sinkVec_shifterReg_55_0_bits_offset <= sinkVec_validSource_55_bits_offset;
        sinkVec_shifterReg_55_0_bits_mask <= sinkVec_validSource_55_bits_mask;
        sinkVec_shifterReg_55_0_bits_data <= sinkVec_validSource_55_bits_data;
        sinkVec_shifterReg_55_0_bits_last <= sinkVec_validSource_55_bits_last;
        sinkVec_shifterReg_55_0_bits_instructionIndex <= sinkVec_validSource_55_bits_instructionIndex;
      end
      maskUnitFirst_27 <= tryToRead_27 & ~(sinkWire_27_ready & sinkWire_27_valid) ^ maskUnitFirst_27;
      view__writeRelease_13_pipe_v <= sinkVec_27_0_ready & sinkVec_27_0_valid;
      pipe_v_39 <= sinkVec_27_1_ready & sinkVec_27_1_valid;
      instructionFinishedPipe_pipe_v_13 <= 1'h1;
      pipe_v_40 <= 1'h1;
      pipe_pipe_v_13 <= pipe_v_40;
      view__laneMaskSelect_13_pipe_v <= 1'h1;
      view__laneMaskSelect_13_pipe_pipe_v <= view__laneMaskSelect_13_pipe_v;
      view__laneMaskSewSelect_13_pipe_v <= 1'h1;
      view__laneMaskSewSelect_13_pipe_pipe_v <= view__laneMaskSewSelect_13_pipe_v;
      lsuLastPipe_pipe_v_13 <= 1'h1;
      maskLastPipe_pipe_v_13 <= 1'h1;
      pipe_v_41 <= 1'h1;
      sinkVec_releasePipe_pipe_v_56 <= sinkVec_sinkWire_56_ready & sinkVec_sinkWire_56_valid;
      if (sinkVec_validSource_56_valid ^ sinkVec_releasePipe_pipe_out_56_valid)
        sinkVec_tokenCheck_counter_56 <= sinkVec_tokenCheck_counter_56 + sinkVec_tokenCheck_counterChange_56;
      if (sinkVec_shifterValid_56) begin
        sinkVec_shifterReg_56_0_valid <= sinkVec_validSource_56_valid;
        sinkVec_shifterReg_56_0_bits_vs <= sinkVec_validSource_56_bits_vs;
        sinkVec_shifterReg_56_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_56_0_bits_offset <= sinkVec_validSource_56_bits_offset;
        sinkVec_shifterReg_56_0_bits_instructionIndex <= sinkVec_validSource_56_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_57 <= sinkVec_sinkWire_57_ready & sinkVec_sinkWire_57_valid;
      if (sinkVec_validSource_57_valid ^ sinkVec_releasePipe_pipe_out_57_valid)
        sinkVec_tokenCheck_counter_57 <= sinkVec_tokenCheck_counter_57 + sinkVec_tokenCheck_counterChange_57;
      if (sinkVec_shifterValid_57) begin
        sinkVec_shifterReg_57_0_valid <= sinkVec_validSource_57_valid;
        sinkVec_shifterReg_57_0_bits_vs <= sinkVec_validSource_57_bits_vs;
        sinkVec_shifterReg_57_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_57_0_bits_offset <= sinkVec_validSource_57_bits_offset;
        sinkVec_shifterReg_57_0_bits_instructionIndex <= sinkVec_validSource_57_bits_instructionIndex;
      end
      maskUnitFirst_28 <= tryToRead_28 & ~(sinkWire_28_ready & sinkWire_28_valid) ^ maskUnitFirst_28;
      accessDataValid_pipe_v_28 <= sinkVec_28_0_ready & sinkVec_28_0_valid;
      accessDataValid_pipe_pipe_v_28 <= accessDataValid_pipe_v_28;
      if (shifterValid_44) begin
        shifterReg_44_0_valid <= accessDataSource_28_valid;
        shifterReg_44_0_bits <= accessDataSource_28_bits;
      end
      accessDataValid_pipe_v_29 <= sinkVec_28_1_ready & sinkVec_28_1_valid;
      accessDataValid_pipe_pipe_v_29 <= accessDataValid_pipe_v_29;
      if (shifterValid_45) begin
        shifterReg_45_0_valid <= accessDataSource_29_valid;
        shifterReg_45_0_bits <= accessDataSource_29_bits;
      end
      sinkVec_releasePipe_pipe_v_58 <= sinkVec_sinkWire_58_ready & sinkVec_sinkWire_58_valid;
      if (sinkVec_validSource_58_valid ^ sinkVec_releasePipe_pipe_out_58_valid)
        sinkVec_tokenCheck_counter_58 <= sinkVec_tokenCheck_counter_58 + sinkVec_tokenCheck_counterChange_58;
      if (sinkVec_shifterValid_58) begin
        sinkVec_shifterReg_58_0_valid <= sinkVec_validSource_58_valid;
        sinkVec_shifterReg_58_0_bits_vd <= sinkVec_validSource_58_bits_vd;
        sinkVec_shifterReg_58_0_bits_offset <= sinkVec_validSource_58_bits_offset;
        sinkVec_shifterReg_58_0_bits_mask <= sinkVec_validSource_58_bits_mask;
        sinkVec_shifterReg_58_0_bits_data <= sinkVec_validSource_58_bits_data;
        sinkVec_shifterReg_58_0_bits_instructionIndex <= sinkVec_validSource_58_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_59 <= sinkVec_sinkWire_59_ready & sinkVec_sinkWire_59_valid;
      if (sinkVec_validSource_59_valid ^ sinkVec_releasePipe_pipe_out_59_valid)
        sinkVec_tokenCheck_counter_59 <= sinkVec_tokenCheck_counter_59 + sinkVec_tokenCheck_counterChange_59;
      if (sinkVec_shifterValid_59) begin
        sinkVec_shifterReg_59_0_valid <= sinkVec_validSource_59_valid;
        sinkVec_shifterReg_59_0_bits_vd <= sinkVec_validSource_59_bits_vd;
        sinkVec_shifterReg_59_0_bits_offset <= sinkVec_validSource_59_bits_offset;
        sinkVec_shifterReg_59_0_bits_mask <= sinkVec_validSource_59_bits_mask;
        sinkVec_shifterReg_59_0_bits_data <= sinkVec_validSource_59_bits_data;
        sinkVec_shifterReg_59_0_bits_last <= sinkVec_validSource_59_bits_last;
        sinkVec_shifterReg_59_0_bits_instructionIndex <= sinkVec_validSource_59_bits_instructionIndex;
      end
      maskUnitFirst_29 <= tryToRead_29 & ~(sinkWire_29_ready & sinkWire_29_valid) ^ maskUnitFirst_29;
      view__writeRelease_14_pipe_v <= sinkVec_29_0_ready & sinkVec_29_0_valid;
      pipe_v_42 <= sinkVec_29_1_ready & sinkVec_29_1_valid;
      instructionFinishedPipe_pipe_v_14 <= 1'h1;
      pipe_v_43 <= 1'h1;
      pipe_pipe_v_14 <= pipe_v_43;
      view__laneMaskSelect_14_pipe_v <= 1'h1;
      view__laneMaskSelect_14_pipe_pipe_v <= view__laneMaskSelect_14_pipe_v;
      view__laneMaskSewSelect_14_pipe_v <= 1'h1;
      view__laneMaskSewSelect_14_pipe_pipe_v <= view__laneMaskSewSelect_14_pipe_v;
      lsuLastPipe_pipe_v_14 <= 1'h1;
      maskLastPipe_pipe_v_14 <= 1'h1;
      pipe_v_44 <= 1'h1;
      sinkVec_releasePipe_pipe_v_60 <= sinkVec_sinkWire_60_ready & sinkVec_sinkWire_60_valid;
      if (sinkVec_validSource_60_valid ^ sinkVec_releasePipe_pipe_out_60_valid)
        sinkVec_tokenCheck_counter_60 <= sinkVec_tokenCheck_counter_60 + sinkVec_tokenCheck_counterChange_60;
      if (sinkVec_shifterValid_60) begin
        sinkVec_shifterReg_60_0_valid <= sinkVec_validSource_60_valid;
        sinkVec_shifterReg_60_0_bits_vs <= sinkVec_validSource_60_bits_vs;
        sinkVec_shifterReg_60_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_60_0_bits_offset <= sinkVec_validSource_60_bits_offset;
        sinkVec_shifterReg_60_0_bits_instructionIndex <= sinkVec_validSource_60_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_61 <= sinkVec_sinkWire_61_ready & sinkVec_sinkWire_61_valid;
      if (sinkVec_validSource_61_valid ^ sinkVec_releasePipe_pipe_out_61_valid)
        sinkVec_tokenCheck_counter_61 <= sinkVec_tokenCheck_counter_61 + sinkVec_tokenCheck_counterChange_61;
      if (sinkVec_shifterValid_61) begin
        sinkVec_shifterReg_61_0_valid <= sinkVec_validSource_61_valid;
        sinkVec_shifterReg_61_0_bits_vs <= sinkVec_validSource_61_bits_vs;
        sinkVec_shifterReg_61_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_61_0_bits_offset <= sinkVec_validSource_61_bits_offset;
        sinkVec_shifterReg_61_0_bits_instructionIndex <= sinkVec_validSource_61_bits_instructionIndex;
      end
      maskUnitFirst_30 <= tryToRead_30 & ~(sinkWire_30_ready & sinkWire_30_valid) ^ maskUnitFirst_30;
      accessDataValid_pipe_v_30 <= sinkVec_30_0_ready & sinkVec_30_0_valid;
      accessDataValid_pipe_pipe_v_30 <= accessDataValid_pipe_v_30;
      if (shifterValid_46) begin
        shifterReg_46_0_valid <= accessDataSource_30_valid;
        shifterReg_46_0_bits <= accessDataSource_30_bits;
      end
      accessDataValid_pipe_v_31 <= sinkVec_30_1_ready & sinkVec_30_1_valid;
      accessDataValid_pipe_pipe_v_31 <= accessDataValid_pipe_v_31;
      if (shifterValid_47) begin
        shifterReg_47_0_valid <= accessDataSource_31_valid;
        shifterReg_47_0_bits <= accessDataSource_31_bits;
      end
      sinkVec_releasePipe_pipe_v_62 <= sinkVec_sinkWire_62_ready & sinkVec_sinkWire_62_valid;
      if (sinkVec_validSource_62_valid ^ sinkVec_releasePipe_pipe_out_62_valid)
        sinkVec_tokenCheck_counter_62 <= sinkVec_tokenCheck_counter_62 + sinkVec_tokenCheck_counterChange_62;
      if (sinkVec_shifterValid_62) begin
        sinkVec_shifterReg_62_0_valid <= sinkVec_validSource_62_valid;
        sinkVec_shifterReg_62_0_bits_vd <= sinkVec_validSource_62_bits_vd;
        sinkVec_shifterReg_62_0_bits_offset <= sinkVec_validSource_62_bits_offset;
        sinkVec_shifterReg_62_0_bits_mask <= sinkVec_validSource_62_bits_mask;
        sinkVec_shifterReg_62_0_bits_data <= sinkVec_validSource_62_bits_data;
        sinkVec_shifterReg_62_0_bits_instructionIndex <= sinkVec_validSource_62_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_63 <= sinkVec_sinkWire_63_ready & sinkVec_sinkWire_63_valid;
      if (sinkVec_validSource_63_valid ^ sinkVec_releasePipe_pipe_out_63_valid)
        sinkVec_tokenCheck_counter_63 <= sinkVec_tokenCheck_counter_63 + sinkVec_tokenCheck_counterChange_63;
      if (sinkVec_shifterValid_63) begin
        sinkVec_shifterReg_63_0_valid <= sinkVec_validSource_63_valid;
        sinkVec_shifterReg_63_0_bits_vd <= sinkVec_validSource_63_bits_vd;
        sinkVec_shifterReg_63_0_bits_offset <= sinkVec_validSource_63_bits_offset;
        sinkVec_shifterReg_63_0_bits_mask <= sinkVec_validSource_63_bits_mask;
        sinkVec_shifterReg_63_0_bits_data <= sinkVec_validSource_63_bits_data;
        sinkVec_shifterReg_63_0_bits_last <= sinkVec_validSource_63_bits_last;
        sinkVec_shifterReg_63_0_bits_instructionIndex <= sinkVec_validSource_63_bits_instructionIndex;
      end
      maskUnitFirst_31 <= tryToRead_31 & ~(sinkWire_31_ready & sinkWire_31_valid) ^ maskUnitFirst_31;
      view__writeRelease_15_pipe_v <= sinkVec_31_0_ready & sinkVec_31_0_valid;
      pipe_v_45 <= sinkVec_31_1_ready & sinkVec_31_1_valid;
      instructionFinishedPipe_pipe_v_15 <= 1'h1;
      pipe_v_46 <= 1'h1;
      pipe_pipe_v_15 <= pipe_v_46;
      view__laneMaskSelect_15_pipe_v <= 1'h1;
      view__laneMaskSelect_15_pipe_pipe_v <= view__laneMaskSelect_15_pipe_v;
      view__laneMaskSewSelect_15_pipe_v <= 1'h1;
      view__laneMaskSewSelect_15_pipe_pipe_v <= view__laneMaskSewSelect_15_pipe_v;
      lsuLastPipe_pipe_v_15 <= 1'h1;
      maskLastPipe_pipe_v_15 <= 1'h1;
      pipe_v_47 <= 1'h1;
      pipe_v_48 <= _laneVec_0_readBusPort_0_enqRelease;
      if (shifterValid_48) begin
        shifterReg_48_0_valid <= _laneVec_0_readBusPort_0_deq_valid;
        shifterReg_48_0_bits_data <= _laneVec_0_readBusPort_0_deq_bits_data;
      end
      pipe_v_49 <= _laneVec_0_writeBusPort_0_enqRelease;
      if (shifterValid_49) begin
        shifterReg_49_0_valid <= _laneVec_0_writeBusPort_0_deq_valid;
        shifterReg_49_0_bits_data <= _laneVec_0_writeBusPort_0_deq_bits_data;
        shifterReg_49_0_bits_mask <= _laneVec_0_writeBusPort_0_deq_bits_mask;
        shifterReg_49_0_bits_instructionIndex <= _laneVec_0_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_49_0_bits_counter <= _laneVec_0_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_50 <= _laneVec_0_readBusPort_1_enqRelease;
      if (shifterValid_50) begin
        shifterReg_50_0_valid <= _laneVec_1_readBusPort_0_deq_valid;
        shifterReg_50_0_bits_data <= _laneVec_1_readBusPort_0_deq_bits_data;
      end
      pipe_v_51 <= _laneVec_1_writeBusPort_0_enqRelease;
      if (shifterValid_51) begin
        shifterReg_51_0_valid <= _laneVec_0_writeBusPort_1_deq_valid;
        shifterReg_51_0_bits_data <= _laneVec_0_writeBusPort_1_deq_bits_data;
        shifterReg_51_0_bits_mask <= _laneVec_0_writeBusPort_1_deq_bits_mask;
        shifterReg_51_0_bits_instructionIndex <= _laneVec_0_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_51_0_bits_counter <= _laneVec_0_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_52 <= _laneVec_1_readBusPort_0_enqRelease;
      if (shifterValid_52) begin
        shifterReg_52_0_valid <= _laneVec_2_readBusPort_0_deq_valid;
        shifterReg_52_0_bits_data <= _laneVec_2_readBusPort_0_deq_bits_data;
      end
      pipe_v_53 <= _laneVec_2_writeBusPort_0_enqRelease;
      if (shifterValid_53) begin
        shifterReg_53_0_valid <= _laneVec_1_writeBusPort_0_deq_valid;
        shifterReg_53_0_bits_data <= _laneVec_1_writeBusPort_0_deq_bits_data;
        shifterReg_53_0_bits_mask <= _laneVec_1_writeBusPort_0_deq_bits_mask;
        shifterReg_53_0_bits_instructionIndex <= _laneVec_1_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_53_0_bits_counter <= _laneVec_1_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_54 <= _laneVec_1_readBusPort_1_enqRelease;
      if (shifterValid_54) begin
        shifterReg_54_0_valid <= _laneVec_3_readBusPort_0_deq_valid;
        shifterReg_54_0_bits_data <= _laneVec_3_readBusPort_0_deq_bits_data;
      end
      pipe_v_55 <= _laneVec_3_writeBusPort_0_enqRelease;
      if (shifterValid_55) begin
        shifterReg_55_0_valid <= _laneVec_1_writeBusPort_1_deq_valid;
        shifterReg_55_0_bits_data <= _laneVec_1_writeBusPort_1_deq_bits_data;
        shifterReg_55_0_bits_mask <= _laneVec_1_writeBusPort_1_deq_bits_mask;
        shifterReg_55_0_bits_instructionIndex <= _laneVec_1_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_55_0_bits_counter <= _laneVec_1_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_56 <= _laneVec_2_readBusPort_0_enqRelease;
      if (shifterValid_56) begin
        shifterReg_56_0_valid <= _laneVec_4_readBusPort_0_deq_valid;
        shifterReg_56_0_bits_data <= _laneVec_4_readBusPort_0_deq_bits_data;
      end
      pipe_v_57 <= _laneVec_4_writeBusPort_0_enqRelease;
      if (shifterValid_57) begin
        shifterReg_57_0_valid <= _laneVec_2_writeBusPort_0_deq_valid;
        shifterReg_57_0_bits_data <= _laneVec_2_writeBusPort_0_deq_bits_data;
        shifterReg_57_0_bits_mask <= _laneVec_2_writeBusPort_0_deq_bits_mask;
        shifterReg_57_0_bits_instructionIndex <= _laneVec_2_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_57_0_bits_counter <= _laneVec_2_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_58 <= _laneVec_2_readBusPort_1_enqRelease;
      if (shifterValid_58) begin
        shifterReg_58_0_valid <= _laneVec_5_readBusPort_0_deq_valid;
        shifterReg_58_0_bits_data <= _laneVec_5_readBusPort_0_deq_bits_data;
      end
      pipe_v_59 <= _laneVec_5_writeBusPort_0_enqRelease;
      if (shifterValid_59) begin
        shifterReg_59_0_valid <= _laneVec_2_writeBusPort_1_deq_valid;
        shifterReg_59_0_bits_data <= _laneVec_2_writeBusPort_1_deq_bits_data;
        shifterReg_59_0_bits_mask <= _laneVec_2_writeBusPort_1_deq_bits_mask;
        shifterReg_59_0_bits_instructionIndex <= _laneVec_2_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_59_0_bits_counter <= _laneVec_2_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_60 <= _laneVec_3_readBusPort_0_enqRelease;
      if (shifterValid_60) begin
        shifterReg_60_0_valid <= _laneVec_6_readBusPort_0_deq_valid;
        shifterReg_60_0_bits_data <= _laneVec_6_readBusPort_0_deq_bits_data;
      end
      pipe_v_61 <= _laneVec_6_writeBusPort_0_enqRelease;
      if (shifterValid_61) begin
        shifterReg_61_0_valid <= _laneVec_3_writeBusPort_0_deq_valid;
        shifterReg_61_0_bits_data <= _laneVec_3_writeBusPort_0_deq_bits_data;
        shifterReg_61_0_bits_mask <= _laneVec_3_writeBusPort_0_deq_bits_mask;
        shifterReg_61_0_bits_instructionIndex <= _laneVec_3_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_61_0_bits_counter <= _laneVec_3_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_62 <= _laneVec_3_readBusPort_1_enqRelease;
      if (shifterValid_62) begin
        shifterReg_62_0_valid <= _laneVec_7_readBusPort_0_deq_valid;
        shifterReg_62_0_bits_data <= _laneVec_7_readBusPort_0_deq_bits_data;
      end
      pipe_v_63 <= _laneVec_7_writeBusPort_0_enqRelease;
      if (shifterValid_63) begin
        shifterReg_63_0_valid <= _laneVec_3_writeBusPort_1_deq_valid;
        shifterReg_63_0_bits_data <= _laneVec_3_writeBusPort_1_deq_bits_data;
        shifterReg_63_0_bits_mask <= _laneVec_3_writeBusPort_1_deq_bits_mask;
        shifterReg_63_0_bits_instructionIndex <= _laneVec_3_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_63_0_bits_counter <= _laneVec_3_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_64 <= _laneVec_4_readBusPort_0_enqRelease;
      if (shifterValid_64) begin
        shifterReg_64_0_valid <= _laneVec_8_readBusPort_0_deq_valid;
        shifterReg_64_0_bits_data <= _laneVec_8_readBusPort_0_deq_bits_data;
      end
      pipe_v_65 <= _laneVec_8_writeBusPort_0_enqRelease;
      if (shifterValid_65) begin
        shifterReg_65_0_valid <= _laneVec_4_writeBusPort_0_deq_valid;
        shifterReg_65_0_bits_data <= _laneVec_4_writeBusPort_0_deq_bits_data;
        shifterReg_65_0_bits_mask <= _laneVec_4_writeBusPort_0_deq_bits_mask;
        shifterReg_65_0_bits_instructionIndex <= _laneVec_4_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_65_0_bits_counter <= _laneVec_4_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_66 <= _laneVec_4_readBusPort_1_enqRelease;
      if (shifterValid_66) begin
        shifterReg_66_0_valid <= _laneVec_9_readBusPort_0_deq_valid;
        shifterReg_66_0_bits_data <= _laneVec_9_readBusPort_0_deq_bits_data;
      end
      pipe_v_67 <= _laneVec_9_writeBusPort_0_enqRelease;
      if (shifterValid_67) begin
        shifterReg_67_0_valid <= _laneVec_4_writeBusPort_1_deq_valid;
        shifterReg_67_0_bits_data <= _laneVec_4_writeBusPort_1_deq_bits_data;
        shifterReg_67_0_bits_mask <= _laneVec_4_writeBusPort_1_deq_bits_mask;
        shifterReg_67_0_bits_instructionIndex <= _laneVec_4_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_67_0_bits_counter <= _laneVec_4_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_68 <= _laneVec_5_readBusPort_0_enqRelease;
      if (shifterValid_68) begin
        shifterReg_68_0_valid <= _laneVec_10_readBusPort_0_deq_valid;
        shifterReg_68_0_bits_data <= _laneVec_10_readBusPort_0_deq_bits_data;
      end
      pipe_v_69 <= _laneVec_10_writeBusPort_0_enqRelease;
      if (shifterValid_69) begin
        shifterReg_69_0_valid <= _laneVec_5_writeBusPort_0_deq_valid;
        shifterReg_69_0_bits_data <= _laneVec_5_writeBusPort_0_deq_bits_data;
        shifterReg_69_0_bits_mask <= _laneVec_5_writeBusPort_0_deq_bits_mask;
        shifterReg_69_0_bits_instructionIndex <= _laneVec_5_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_69_0_bits_counter <= _laneVec_5_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_70 <= _laneVec_5_readBusPort_1_enqRelease;
      if (shifterValid_70) begin
        shifterReg_70_0_valid <= _laneVec_11_readBusPort_0_deq_valid;
        shifterReg_70_0_bits_data <= _laneVec_11_readBusPort_0_deq_bits_data;
      end
      pipe_v_71 <= _laneVec_11_writeBusPort_0_enqRelease;
      if (shifterValid_71) begin
        shifterReg_71_0_valid <= _laneVec_5_writeBusPort_1_deq_valid;
        shifterReg_71_0_bits_data <= _laneVec_5_writeBusPort_1_deq_bits_data;
        shifterReg_71_0_bits_mask <= _laneVec_5_writeBusPort_1_deq_bits_mask;
        shifterReg_71_0_bits_instructionIndex <= _laneVec_5_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_71_0_bits_counter <= _laneVec_5_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_72 <= _laneVec_6_readBusPort_0_enqRelease;
      if (shifterValid_72) begin
        shifterReg_72_0_valid <= _laneVec_12_readBusPort_0_deq_valid;
        shifterReg_72_0_bits_data <= _laneVec_12_readBusPort_0_deq_bits_data;
      end
      pipe_v_73 <= _laneVec_12_writeBusPort_0_enqRelease;
      if (shifterValid_73) begin
        shifterReg_73_0_valid <= _laneVec_6_writeBusPort_0_deq_valid;
        shifterReg_73_0_bits_data <= _laneVec_6_writeBusPort_0_deq_bits_data;
        shifterReg_73_0_bits_mask <= _laneVec_6_writeBusPort_0_deq_bits_mask;
        shifterReg_73_0_bits_instructionIndex <= _laneVec_6_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_73_0_bits_counter <= _laneVec_6_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_74 <= _laneVec_6_readBusPort_1_enqRelease;
      if (shifterValid_74) begin
        shifterReg_74_0_valid <= _laneVec_13_readBusPort_0_deq_valid;
        shifterReg_74_0_bits_data <= _laneVec_13_readBusPort_0_deq_bits_data;
      end
      pipe_v_75 <= _laneVec_13_writeBusPort_0_enqRelease;
      if (shifterValid_75) begin
        shifterReg_75_0_valid <= _laneVec_6_writeBusPort_1_deq_valid;
        shifterReg_75_0_bits_data <= _laneVec_6_writeBusPort_1_deq_bits_data;
        shifterReg_75_0_bits_mask <= _laneVec_6_writeBusPort_1_deq_bits_mask;
        shifterReg_75_0_bits_instructionIndex <= _laneVec_6_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_75_0_bits_counter <= _laneVec_6_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_76 <= _laneVec_7_readBusPort_0_enqRelease;
      if (shifterValid_76) begin
        shifterReg_76_0_valid <= _laneVec_14_readBusPort_0_deq_valid;
        shifterReg_76_0_bits_data <= _laneVec_14_readBusPort_0_deq_bits_data;
      end
      pipe_v_77 <= _laneVec_14_writeBusPort_0_enqRelease;
      if (shifterValid_77) begin
        shifterReg_77_0_valid <= _laneVec_7_writeBusPort_0_deq_valid;
        shifterReg_77_0_bits_data <= _laneVec_7_writeBusPort_0_deq_bits_data;
        shifterReg_77_0_bits_mask <= _laneVec_7_writeBusPort_0_deq_bits_mask;
        shifterReg_77_0_bits_instructionIndex <= _laneVec_7_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_77_0_bits_counter <= _laneVec_7_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_78 <= _laneVec_7_readBusPort_1_enqRelease;
      if (shifterValid_78) begin
        shifterReg_78_0_valid <= _laneVec_15_readBusPort_0_deq_valid;
        shifterReg_78_0_bits_data <= _laneVec_15_readBusPort_0_deq_bits_data;
      end
      pipe_v_79 <= _laneVec_15_writeBusPort_0_enqRelease;
      if (shifterValid_79) begin
        shifterReg_79_0_valid <= _laneVec_7_writeBusPort_1_deq_valid;
        shifterReg_79_0_bits_data <= _laneVec_7_writeBusPort_1_deq_bits_data;
        shifterReg_79_0_bits_mask <= _laneVec_7_writeBusPort_1_deq_bits_mask;
        shifterReg_79_0_bits_instructionIndex <= _laneVec_7_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_79_0_bits_counter <= _laneVec_7_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_80 <= _laneVec_8_readBusPort_0_enqRelease;
      if (shifterValid_80) begin
        shifterReg_80_0_valid <= _laneVec_0_readBusPort_1_deq_valid;
        shifterReg_80_0_bits_data <= _laneVec_0_readBusPort_1_deq_bits_data;
      end
      pipe_v_81 <= _laneVec_0_writeBusPort_1_enqRelease;
      if (shifterValid_81) begin
        shifterReg_81_0_valid <= _laneVec_8_writeBusPort_0_deq_valid;
        shifterReg_81_0_bits_data <= _laneVec_8_writeBusPort_0_deq_bits_data;
        shifterReg_81_0_bits_mask <= _laneVec_8_writeBusPort_0_deq_bits_mask;
        shifterReg_81_0_bits_instructionIndex <= _laneVec_8_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_81_0_bits_counter <= _laneVec_8_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_82 <= _laneVec_8_readBusPort_1_enqRelease;
      if (shifterValid_82) begin
        shifterReg_82_0_valid <= _laneVec_1_readBusPort_1_deq_valid;
        shifterReg_82_0_bits_data <= _laneVec_1_readBusPort_1_deq_bits_data;
      end
      pipe_v_83 <= _laneVec_1_writeBusPort_1_enqRelease;
      if (shifterValid_83) begin
        shifterReg_83_0_valid <= _laneVec_8_writeBusPort_1_deq_valid;
        shifterReg_83_0_bits_data <= _laneVec_8_writeBusPort_1_deq_bits_data;
        shifterReg_83_0_bits_mask <= _laneVec_8_writeBusPort_1_deq_bits_mask;
        shifterReg_83_0_bits_instructionIndex <= _laneVec_8_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_83_0_bits_counter <= _laneVec_8_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_84 <= _laneVec_9_readBusPort_0_enqRelease;
      if (shifterValid_84) begin
        shifterReg_84_0_valid <= _laneVec_2_readBusPort_1_deq_valid;
        shifterReg_84_0_bits_data <= _laneVec_2_readBusPort_1_deq_bits_data;
      end
      pipe_v_85 <= _laneVec_2_writeBusPort_1_enqRelease;
      if (shifterValid_85) begin
        shifterReg_85_0_valid <= _laneVec_9_writeBusPort_0_deq_valid;
        shifterReg_85_0_bits_data <= _laneVec_9_writeBusPort_0_deq_bits_data;
        shifterReg_85_0_bits_mask <= _laneVec_9_writeBusPort_0_deq_bits_mask;
        shifterReg_85_0_bits_instructionIndex <= _laneVec_9_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_85_0_bits_counter <= _laneVec_9_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_86 <= _laneVec_9_readBusPort_1_enqRelease;
      if (shifterValid_86) begin
        shifterReg_86_0_valid <= _laneVec_3_readBusPort_1_deq_valid;
        shifterReg_86_0_bits_data <= _laneVec_3_readBusPort_1_deq_bits_data;
      end
      pipe_v_87 <= _laneVec_3_writeBusPort_1_enqRelease;
      if (shifterValid_87) begin
        shifterReg_87_0_valid <= _laneVec_9_writeBusPort_1_deq_valid;
        shifterReg_87_0_bits_data <= _laneVec_9_writeBusPort_1_deq_bits_data;
        shifterReg_87_0_bits_mask <= _laneVec_9_writeBusPort_1_deq_bits_mask;
        shifterReg_87_0_bits_instructionIndex <= _laneVec_9_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_87_0_bits_counter <= _laneVec_9_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_88 <= _laneVec_10_readBusPort_0_enqRelease;
      if (shifterValid_88) begin
        shifterReg_88_0_valid <= _laneVec_4_readBusPort_1_deq_valid;
        shifterReg_88_0_bits_data <= _laneVec_4_readBusPort_1_deq_bits_data;
      end
      pipe_v_89 <= _laneVec_4_writeBusPort_1_enqRelease;
      if (shifterValid_89) begin
        shifterReg_89_0_valid <= _laneVec_10_writeBusPort_0_deq_valid;
        shifterReg_89_0_bits_data <= _laneVec_10_writeBusPort_0_deq_bits_data;
        shifterReg_89_0_bits_mask <= _laneVec_10_writeBusPort_0_deq_bits_mask;
        shifterReg_89_0_bits_instructionIndex <= _laneVec_10_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_89_0_bits_counter <= _laneVec_10_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_90 <= _laneVec_10_readBusPort_1_enqRelease;
      if (shifterValid_90) begin
        shifterReg_90_0_valid <= _laneVec_5_readBusPort_1_deq_valid;
        shifterReg_90_0_bits_data <= _laneVec_5_readBusPort_1_deq_bits_data;
      end
      pipe_v_91 <= _laneVec_5_writeBusPort_1_enqRelease;
      if (shifterValid_91) begin
        shifterReg_91_0_valid <= _laneVec_10_writeBusPort_1_deq_valid;
        shifterReg_91_0_bits_data <= _laneVec_10_writeBusPort_1_deq_bits_data;
        shifterReg_91_0_bits_mask <= _laneVec_10_writeBusPort_1_deq_bits_mask;
        shifterReg_91_0_bits_instructionIndex <= _laneVec_10_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_91_0_bits_counter <= _laneVec_10_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_92 <= _laneVec_11_readBusPort_0_enqRelease;
      if (shifterValid_92) begin
        shifterReg_92_0_valid <= _laneVec_6_readBusPort_1_deq_valid;
        shifterReg_92_0_bits_data <= _laneVec_6_readBusPort_1_deq_bits_data;
      end
      pipe_v_93 <= _laneVec_6_writeBusPort_1_enqRelease;
      if (shifterValid_93) begin
        shifterReg_93_0_valid <= _laneVec_11_writeBusPort_0_deq_valid;
        shifterReg_93_0_bits_data <= _laneVec_11_writeBusPort_0_deq_bits_data;
        shifterReg_93_0_bits_mask <= _laneVec_11_writeBusPort_0_deq_bits_mask;
        shifterReg_93_0_bits_instructionIndex <= _laneVec_11_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_93_0_bits_counter <= _laneVec_11_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_94 <= _laneVec_11_readBusPort_1_enqRelease;
      if (shifterValid_94) begin
        shifterReg_94_0_valid <= _laneVec_7_readBusPort_1_deq_valid;
        shifterReg_94_0_bits_data <= _laneVec_7_readBusPort_1_deq_bits_data;
      end
      pipe_v_95 <= _laneVec_7_writeBusPort_1_enqRelease;
      if (shifterValid_95) begin
        shifterReg_95_0_valid <= _laneVec_11_writeBusPort_1_deq_valid;
        shifterReg_95_0_bits_data <= _laneVec_11_writeBusPort_1_deq_bits_data;
        shifterReg_95_0_bits_mask <= _laneVec_11_writeBusPort_1_deq_bits_mask;
        shifterReg_95_0_bits_instructionIndex <= _laneVec_11_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_95_0_bits_counter <= _laneVec_11_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_96 <= _laneVec_12_readBusPort_0_enqRelease;
      if (shifterValid_96) begin
        shifterReg_96_0_valid <= _laneVec_8_readBusPort_1_deq_valid;
        shifterReg_96_0_bits_data <= _laneVec_8_readBusPort_1_deq_bits_data;
      end
      pipe_v_97 <= _laneVec_8_writeBusPort_1_enqRelease;
      if (shifterValid_97) begin
        shifterReg_97_0_valid <= _laneVec_12_writeBusPort_0_deq_valid;
        shifterReg_97_0_bits_data <= _laneVec_12_writeBusPort_0_deq_bits_data;
        shifterReg_97_0_bits_mask <= _laneVec_12_writeBusPort_0_deq_bits_mask;
        shifterReg_97_0_bits_instructionIndex <= _laneVec_12_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_97_0_bits_counter <= _laneVec_12_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_98 <= _laneVec_12_readBusPort_1_enqRelease;
      if (shifterValid_98) begin
        shifterReg_98_0_valid <= _laneVec_9_readBusPort_1_deq_valid;
        shifterReg_98_0_bits_data <= _laneVec_9_readBusPort_1_deq_bits_data;
      end
      pipe_v_99 <= _laneVec_9_writeBusPort_1_enqRelease;
      if (shifterValid_99) begin
        shifterReg_99_0_valid <= _laneVec_12_writeBusPort_1_deq_valid;
        shifterReg_99_0_bits_data <= _laneVec_12_writeBusPort_1_deq_bits_data;
        shifterReg_99_0_bits_mask <= _laneVec_12_writeBusPort_1_deq_bits_mask;
        shifterReg_99_0_bits_instructionIndex <= _laneVec_12_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_99_0_bits_counter <= _laneVec_12_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_100 <= _laneVec_13_readBusPort_0_enqRelease;
      if (shifterValid_100) begin
        shifterReg_100_0_valid <= _laneVec_10_readBusPort_1_deq_valid;
        shifterReg_100_0_bits_data <= _laneVec_10_readBusPort_1_deq_bits_data;
      end
      pipe_v_101 <= _laneVec_10_writeBusPort_1_enqRelease;
      if (shifterValid_101) begin
        shifterReg_101_0_valid <= _laneVec_13_writeBusPort_0_deq_valid;
        shifterReg_101_0_bits_data <= _laneVec_13_writeBusPort_0_deq_bits_data;
        shifterReg_101_0_bits_mask <= _laneVec_13_writeBusPort_0_deq_bits_mask;
        shifterReg_101_0_bits_instructionIndex <= _laneVec_13_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_101_0_bits_counter <= _laneVec_13_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_102 <= _laneVec_13_readBusPort_1_enqRelease;
      if (shifterValid_102) begin
        shifterReg_102_0_valid <= _laneVec_11_readBusPort_1_deq_valid;
        shifterReg_102_0_bits_data <= _laneVec_11_readBusPort_1_deq_bits_data;
      end
      pipe_v_103 <= _laneVec_11_writeBusPort_1_enqRelease;
      if (shifterValid_103) begin
        shifterReg_103_0_valid <= _laneVec_13_writeBusPort_1_deq_valid;
        shifterReg_103_0_bits_data <= _laneVec_13_writeBusPort_1_deq_bits_data;
        shifterReg_103_0_bits_mask <= _laneVec_13_writeBusPort_1_deq_bits_mask;
        shifterReg_103_0_bits_instructionIndex <= _laneVec_13_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_103_0_bits_counter <= _laneVec_13_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_104 <= _laneVec_14_readBusPort_0_enqRelease;
      if (shifterValid_104) begin
        shifterReg_104_0_valid <= _laneVec_12_readBusPort_1_deq_valid;
        shifterReg_104_0_bits_data <= _laneVec_12_readBusPort_1_deq_bits_data;
      end
      pipe_v_105 <= _laneVec_12_writeBusPort_1_enqRelease;
      if (shifterValid_105) begin
        shifterReg_105_0_valid <= _laneVec_14_writeBusPort_0_deq_valid;
        shifterReg_105_0_bits_data <= _laneVec_14_writeBusPort_0_deq_bits_data;
        shifterReg_105_0_bits_mask <= _laneVec_14_writeBusPort_0_deq_bits_mask;
        shifterReg_105_0_bits_instructionIndex <= _laneVec_14_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_105_0_bits_counter <= _laneVec_14_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_106 <= _laneVec_14_readBusPort_1_enqRelease;
      if (shifterValid_106) begin
        shifterReg_106_0_valid <= _laneVec_13_readBusPort_1_deq_valid;
        shifterReg_106_0_bits_data <= _laneVec_13_readBusPort_1_deq_bits_data;
      end
      pipe_v_107 <= _laneVec_13_writeBusPort_1_enqRelease;
      if (shifterValid_107) begin
        shifterReg_107_0_valid <= _laneVec_14_writeBusPort_1_deq_valid;
        shifterReg_107_0_bits_data <= _laneVec_14_writeBusPort_1_deq_bits_data;
        shifterReg_107_0_bits_mask <= _laneVec_14_writeBusPort_1_deq_bits_mask;
        shifterReg_107_0_bits_instructionIndex <= _laneVec_14_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_107_0_bits_counter <= _laneVec_14_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_108 <= _laneVec_15_readBusPort_0_enqRelease;
      if (shifterValid_108) begin
        shifterReg_108_0_valid <= _laneVec_14_readBusPort_1_deq_valid;
        shifterReg_108_0_bits_data <= _laneVec_14_readBusPort_1_deq_bits_data;
      end
      pipe_v_109 <= _laneVec_14_writeBusPort_1_enqRelease;
      if (shifterValid_109) begin
        shifterReg_109_0_valid <= _laneVec_15_writeBusPort_0_deq_valid;
        shifterReg_109_0_bits_data <= _laneVec_15_writeBusPort_0_deq_bits_data;
        shifterReg_109_0_bits_mask <= _laneVec_15_writeBusPort_0_deq_bits_mask;
        shifterReg_109_0_bits_instructionIndex <= _laneVec_15_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_109_0_bits_counter <= _laneVec_15_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_110 <= _laneVec_15_readBusPort_1_enqRelease;
      if (shifterValid_110) begin
        shifterReg_110_0_valid <= _laneVec_15_readBusPort_1_deq_valid;
        shifterReg_110_0_bits_data <= _laneVec_15_readBusPort_1_deq_bits_data;
      end
      pipe_v_111 <= _laneVec_15_writeBusPort_1_enqRelease;
      if (shifterValid_111) begin
        shifterReg_111_0_valid <= _laneVec_15_writeBusPort_1_deq_valid;
        shifterReg_111_0_bits_data <= _laneVec_15_writeBusPort_1_deq_bits_data;
        shifterReg_111_0_bits_mask <= _laneVec_15_writeBusPort_1_deq_bits_mask;
        shifterReg_111_0_bits_instructionIndex <= _laneVec_15_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_111_0_bits_counter <= _laneVec_15_writeBusPort_1_deq_bits_counter;
      end
    end
    instructionFinishedPipe_pipe_b <= _laneVec_0_instructionFinished;
    pipe_b_1 <= _maskUnit_laneMaskInput_0;
    if (pipe_v_1)
      pipe_pipe_b <= pipe_b_1;
    view__laneMaskSelect_0_pipe_b <= _laneVec_0_maskSelect;
    if (view__laneMaskSelect_0_pipe_v)
      view__laneMaskSelect_0_pipe_pipe_b <= view__laneMaskSelect_0_pipe_b;
    view__laneMaskSewSelect_0_pipe_b <= _laneVec_0_maskSelectSew;
    if (view__laneMaskSewSelect_0_pipe_v)
      view__laneMaskSewSelect_0_pipe_pipe_b <= view__laneMaskSewSelect_0_pipe_b;
    lsuLastPipe_pipe_b <= _lsu_lastReport;
    maskLastPipe_pipe_b <= _maskUnit_lastReport;
    pipe_b_2 <= writeCounter;
    instructionFinishedPipe_pipe_b_1 <= _laneVec_1_instructionFinished;
    pipe_b_4 <= _maskUnit_laneMaskInput_1;
    if (pipe_v_4)
      pipe_pipe_b_1 <= pipe_b_4;
    view__laneMaskSelect_1_pipe_b <= _laneVec_1_maskSelect;
    if (view__laneMaskSelect_1_pipe_v)
      view__laneMaskSelect_1_pipe_pipe_b <= view__laneMaskSelect_1_pipe_b;
    view__laneMaskSewSelect_1_pipe_b <= _laneVec_1_maskSelectSew;
    if (view__laneMaskSewSelect_1_pipe_v)
      view__laneMaskSewSelect_1_pipe_pipe_b <= view__laneMaskSewSelect_1_pipe_b;
    lsuLastPipe_pipe_b_1 <= _lsu_lastReport;
    maskLastPipe_pipe_b_1 <= _maskUnit_lastReport;
    pipe_b_5 <= writeCounter_1;
    instructionFinishedPipe_pipe_b_2 <= _laneVec_2_instructionFinished;
    pipe_b_7 <= _maskUnit_laneMaskInput_2;
    if (pipe_v_7)
      pipe_pipe_b_2 <= pipe_b_7;
    view__laneMaskSelect_2_pipe_b <= _laneVec_2_maskSelect;
    if (view__laneMaskSelect_2_pipe_v)
      view__laneMaskSelect_2_pipe_pipe_b <= view__laneMaskSelect_2_pipe_b;
    view__laneMaskSewSelect_2_pipe_b <= _laneVec_2_maskSelectSew;
    if (view__laneMaskSewSelect_2_pipe_v)
      view__laneMaskSewSelect_2_pipe_pipe_b <= view__laneMaskSewSelect_2_pipe_b;
    lsuLastPipe_pipe_b_2 <= _lsu_lastReport;
    maskLastPipe_pipe_b_2 <= _maskUnit_lastReport;
    pipe_b_8 <= writeCounter_2;
    instructionFinishedPipe_pipe_b_3 <= _laneVec_3_instructionFinished;
    pipe_b_10 <= _maskUnit_laneMaskInput_3;
    if (pipe_v_10)
      pipe_pipe_b_3 <= pipe_b_10;
    view__laneMaskSelect_3_pipe_b <= _laneVec_3_maskSelect;
    if (view__laneMaskSelect_3_pipe_v)
      view__laneMaskSelect_3_pipe_pipe_b <= view__laneMaskSelect_3_pipe_b;
    view__laneMaskSewSelect_3_pipe_b <= _laneVec_3_maskSelectSew;
    if (view__laneMaskSewSelect_3_pipe_v)
      view__laneMaskSewSelect_3_pipe_pipe_b <= view__laneMaskSewSelect_3_pipe_b;
    lsuLastPipe_pipe_b_3 <= _lsu_lastReport;
    maskLastPipe_pipe_b_3 <= _maskUnit_lastReport;
    pipe_b_11 <= writeCounter_3;
    instructionFinishedPipe_pipe_b_4 <= _laneVec_4_instructionFinished;
    pipe_b_13 <= _maskUnit_laneMaskInput_4;
    if (pipe_v_13)
      pipe_pipe_b_4 <= pipe_b_13;
    view__laneMaskSelect_4_pipe_b <= _laneVec_4_maskSelect;
    if (view__laneMaskSelect_4_pipe_v)
      view__laneMaskSelect_4_pipe_pipe_b <= view__laneMaskSelect_4_pipe_b;
    view__laneMaskSewSelect_4_pipe_b <= _laneVec_4_maskSelectSew;
    if (view__laneMaskSewSelect_4_pipe_v)
      view__laneMaskSewSelect_4_pipe_pipe_b <= view__laneMaskSewSelect_4_pipe_b;
    lsuLastPipe_pipe_b_4 <= _lsu_lastReport;
    maskLastPipe_pipe_b_4 <= _maskUnit_lastReport;
    pipe_b_14 <= writeCounter_4;
    instructionFinishedPipe_pipe_b_5 <= _laneVec_5_instructionFinished;
    pipe_b_16 <= _maskUnit_laneMaskInput_5;
    if (pipe_v_16)
      pipe_pipe_b_5 <= pipe_b_16;
    view__laneMaskSelect_5_pipe_b <= _laneVec_5_maskSelect;
    if (view__laneMaskSelect_5_pipe_v)
      view__laneMaskSelect_5_pipe_pipe_b <= view__laneMaskSelect_5_pipe_b;
    view__laneMaskSewSelect_5_pipe_b <= _laneVec_5_maskSelectSew;
    if (view__laneMaskSewSelect_5_pipe_v)
      view__laneMaskSewSelect_5_pipe_pipe_b <= view__laneMaskSewSelect_5_pipe_b;
    lsuLastPipe_pipe_b_5 <= _lsu_lastReport;
    maskLastPipe_pipe_b_5 <= _maskUnit_lastReport;
    pipe_b_17 <= writeCounter_5;
    instructionFinishedPipe_pipe_b_6 <= _laneVec_6_instructionFinished;
    pipe_b_19 <= _maskUnit_laneMaskInput_6;
    if (pipe_v_19)
      pipe_pipe_b_6 <= pipe_b_19;
    view__laneMaskSelect_6_pipe_b <= _laneVec_6_maskSelect;
    if (view__laneMaskSelect_6_pipe_v)
      view__laneMaskSelect_6_pipe_pipe_b <= view__laneMaskSelect_6_pipe_b;
    view__laneMaskSewSelect_6_pipe_b <= _laneVec_6_maskSelectSew;
    if (view__laneMaskSewSelect_6_pipe_v)
      view__laneMaskSewSelect_6_pipe_pipe_b <= view__laneMaskSewSelect_6_pipe_b;
    lsuLastPipe_pipe_b_6 <= _lsu_lastReport;
    maskLastPipe_pipe_b_6 <= _maskUnit_lastReport;
    pipe_b_20 <= writeCounter_6;
    instructionFinishedPipe_pipe_b_7 <= _laneVec_7_instructionFinished;
    pipe_b_22 <= _maskUnit_laneMaskInput_7;
    if (pipe_v_22)
      pipe_pipe_b_7 <= pipe_b_22;
    view__laneMaskSelect_7_pipe_b <= _laneVec_7_maskSelect;
    if (view__laneMaskSelect_7_pipe_v)
      view__laneMaskSelect_7_pipe_pipe_b <= view__laneMaskSelect_7_pipe_b;
    view__laneMaskSewSelect_7_pipe_b <= _laneVec_7_maskSelectSew;
    if (view__laneMaskSewSelect_7_pipe_v)
      view__laneMaskSewSelect_7_pipe_pipe_b <= view__laneMaskSewSelect_7_pipe_b;
    lsuLastPipe_pipe_b_7 <= _lsu_lastReport;
    maskLastPipe_pipe_b_7 <= _maskUnit_lastReport;
    pipe_b_23 <= writeCounter_7;
    instructionFinishedPipe_pipe_b_8 <= _laneVec_8_instructionFinished;
    pipe_b_25 <= _maskUnit_laneMaskInput_8;
    if (pipe_v_25)
      pipe_pipe_b_8 <= pipe_b_25;
    view__laneMaskSelect_8_pipe_b <= _laneVec_8_maskSelect;
    if (view__laneMaskSelect_8_pipe_v)
      view__laneMaskSelect_8_pipe_pipe_b <= view__laneMaskSelect_8_pipe_b;
    view__laneMaskSewSelect_8_pipe_b <= _laneVec_8_maskSelectSew;
    if (view__laneMaskSewSelect_8_pipe_v)
      view__laneMaskSewSelect_8_pipe_pipe_b <= view__laneMaskSewSelect_8_pipe_b;
    lsuLastPipe_pipe_b_8 <= _lsu_lastReport;
    maskLastPipe_pipe_b_8 <= _maskUnit_lastReport;
    pipe_b_26 <= writeCounter_8;
    instructionFinishedPipe_pipe_b_9 <= _laneVec_9_instructionFinished;
    pipe_b_28 <= _maskUnit_laneMaskInput_9;
    if (pipe_v_28)
      pipe_pipe_b_9 <= pipe_b_28;
    view__laneMaskSelect_9_pipe_b <= _laneVec_9_maskSelect;
    if (view__laneMaskSelect_9_pipe_v)
      view__laneMaskSelect_9_pipe_pipe_b <= view__laneMaskSelect_9_pipe_b;
    view__laneMaskSewSelect_9_pipe_b <= _laneVec_9_maskSelectSew;
    if (view__laneMaskSewSelect_9_pipe_v)
      view__laneMaskSewSelect_9_pipe_pipe_b <= view__laneMaskSewSelect_9_pipe_b;
    lsuLastPipe_pipe_b_9 <= _lsu_lastReport;
    maskLastPipe_pipe_b_9 <= _maskUnit_lastReport;
    pipe_b_29 <= writeCounter_9;
    instructionFinishedPipe_pipe_b_10 <= _laneVec_10_instructionFinished;
    pipe_b_31 <= _maskUnit_laneMaskInput_10;
    if (pipe_v_31)
      pipe_pipe_b_10 <= pipe_b_31;
    view__laneMaskSelect_10_pipe_b <= _laneVec_10_maskSelect;
    if (view__laneMaskSelect_10_pipe_v)
      view__laneMaskSelect_10_pipe_pipe_b <= view__laneMaskSelect_10_pipe_b;
    view__laneMaskSewSelect_10_pipe_b <= _laneVec_10_maskSelectSew;
    if (view__laneMaskSewSelect_10_pipe_v)
      view__laneMaskSewSelect_10_pipe_pipe_b <= view__laneMaskSewSelect_10_pipe_b;
    lsuLastPipe_pipe_b_10 <= _lsu_lastReport;
    maskLastPipe_pipe_b_10 <= _maskUnit_lastReport;
    pipe_b_32 <= writeCounter_10;
    instructionFinishedPipe_pipe_b_11 <= _laneVec_11_instructionFinished;
    pipe_b_34 <= _maskUnit_laneMaskInput_11;
    if (pipe_v_34)
      pipe_pipe_b_11 <= pipe_b_34;
    view__laneMaskSelect_11_pipe_b <= _laneVec_11_maskSelect;
    if (view__laneMaskSelect_11_pipe_v)
      view__laneMaskSelect_11_pipe_pipe_b <= view__laneMaskSelect_11_pipe_b;
    view__laneMaskSewSelect_11_pipe_b <= _laneVec_11_maskSelectSew;
    if (view__laneMaskSewSelect_11_pipe_v)
      view__laneMaskSewSelect_11_pipe_pipe_b <= view__laneMaskSewSelect_11_pipe_b;
    lsuLastPipe_pipe_b_11 <= _lsu_lastReport;
    maskLastPipe_pipe_b_11 <= _maskUnit_lastReport;
    pipe_b_35 <= writeCounter_11;
    instructionFinishedPipe_pipe_b_12 <= _laneVec_12_instructionFinished;
    pipe_b_37 <= _maskUnit_laneMaskInput_12;
    if (pipe_v_37)
      pipe_pipe_b_12 <= pipe_b_37;
    view__laneMaskSelect_12_pipe_b <= _laneVec_12_maskSelect;
    if (view__laneMaskSelect_12_pipe_v)
      view__laneMaskSelect_12_pipe_pipe_b <= view__laneMaskSelect_12_pipe_b;
    view__laneMaskSewSelect_12_pipe_b <= _laneVec_12_maskSelectSew;
    if (view__laneMaskSewSelect_12_pipe_v)
      view__laneMaskSewSelect_12_pipe_pipe_b <= view__laneMaskSewSelect_12_pipe_b;
    lsuLastPipe_pipe_b_12 <= _lsu_lastReport;
    maskLastPipe_pipe_b_12 <= _maskUnit_lastReport;
    pipe_b_38 <= writeCounter_12;
    instructionFinishedPipe_pipe_b_13 <= _laneVec_13_instructionFinished;
    pipe_b_40 <= _maskUnit_laneMaskInput_13;
    if (pipe_v_40)
      pipe_pipe_b_13 <= pipe_b_40;
    view__laneMaskSelect_13_pipe_b <= _laneVec_13_maskSelect;
    if (view__laneMaskSelect_13_pipe_v)
      view__laneMaskSelect_13_pipe_pipe_b <= view__laneMaskSelect_13_pipe_b;
    view__laneMaskSewSelect_13_pipe_b <= _laneVec_13_maskSelectSew;
    if (view__laneMaskSewSelect_13_pipe_v)
      view__laneMaskSewSelect_13_pipe_pipe_b <= view__laneMaskSewSelect_13_pipe_b;
    lsuLastPipe_pipe_b_13 <= _lsu_lastReport;
    maskLastPipe_pipe_b_13 <= _maskUnit_lastReport;
    pipe_b_41 <= writeCounter_13;
    instructionFinishedPipe_pipe_b_14 <= _laneVec_14_instructionFinished;
    pipe_b_43 <= _maskUnit_laneMaskInput_14;
    if (pipe_v_43)
      pipe_pipe_b_14 <= pipe_b_43;
    view__laneMaskSelect_14_pipe_b <= _laneVec_14_maskSelect;
    if (view__laneMaskSelect_14_pipe_v)
      view__laneMaskSelect_14_pipe_pipe_b <= view__laneMaskSelect_14_pipe_b;
    view__laneMaskSewSelect_14_pipe_b <= _laneVec_14_maskSelectSew;
    if (view__laneMaskSewSelect_14_pipe_v)
      view__laneMaskSewSelect_14_pipe_pipe_b <= view__laneMaskSewSelect_14_pipe_b;
    lsuLastPipe_pipe_b_14 <= _lsu_lastReport;
    maskLastPipe_pipe_b_14 <= _maskUnit_lastReport;
    pipe_b_44 <= writeCounter_14;
    instructionFinishedPipe_pipe_b_15 <= _laneVec_15_instructionFinished;
    pipe_b_46 <= _maskUnit_laneMaskInput_15;
    if (pipe_v_46)
      pipe_pipe_b_15 <= pipe_b_46;
    view__laneMaskSelect_15_pipe_b <= _laneVec_15_maskSelect;
    if (view__laneMaskSelect_15_pipe_v)
      view__laneMaskSelect_15_pipe_pipe_b <= view__laneMaskSelect_15_pipe_b;
    view__laneMaskSewSelect_15_pipe_b <= _laneVec_15_maskSelectSew;
    if (view__laneMaskSewSelect_15_pipe_v)
      view__laneMaskSewSelect_15_pipe_pipe_b <= view__laneMaskSewSelect_15_pipe_b;
    lsuLastPipe_pipe_b_15 <= _lsu_lastReport;
    maskLastPipe_pipe_b_15 <= _maskUnit_lastReport;
    pipe_b_47 <= writeCounter_15;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:336];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h151; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        instructionCounter = _RANDOM[9'h0][2:0];
        responseCounter = _RANDOM[9'h0][5:3];
        requestReg_valid = _RANDOM[9'h0][6];
        requestReg_bits_issue_instruction = {_RANDOM[9'h0][31:7], _RANDOM[9'h1][6:0]};
        requestReg_bits_issue_rs1Data = {_RANDOM[9'h1][31:7], _RANDOM[9'h2][6:0]};
        requestReg_bits_issue_rs2Data = {_RANDOM[9'h2][31:7], _RANDOM[9'h3][6:0]};
        requestReg_bits_issue_vtype = {_RANDOM[9'h3][31:7], _RANDOM[9'h4][6:0]};
        requestReg_bits_issue_vl = {_RANDOM[9'h4][31:7], _RANDOM[9'h5][6:0]};
        requestReg_bits_issue_vstart = {_RANDOM[9'h5][31:7], _RANDOM[9'h6][6:0]};
        requestReg_bits_issue_vcsr = {_RANDOM[9'h6][31:7], _RANDOM[9'h7][6:0]};
        requestReg_bits_decodeResult_orderReduce = _RANDOM[9'h7][7];
        requestReg_bits_decodeResult_floatMul = _RANDOM[9'h7][8];
        requestReg_bits_decodeResult_fpExecutionType = _RANDOM[9'h7][10:9];
        requestReg_bits_decodeResult_float = _RANDOM[9'h7][11];
        requestReg_bits_decodeResult_specialSlot = _RANDOM[9'h7][12];
        requestReg_bits_decodeResult_topUop = _RANDOM[9'h7][17:13];
        requestReg_bits_decodeResult_popCount = _RANDOM[9'h7][18];
        requestReg_bits_decodeResult_ffo = _RANDOM[9'h7][19];
        requestReg_bits_decodeResult_average = _RANDOM[9'h7][20];
        requestReg_bits_decodeResult_reverse = _RANDOM[9'h7][21];
        requestReg_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h7][22];
        requestReg_bits_decodeResult_scheduler = _RANDOM[9'h7][23];
        requestReg_bits_decodeResult_sReadVD = _RANDOM[9'h7][24];
        requestReg_bits_decodeResult_vtype = _RANDOM[9'h7][25];
        requestReg_bits_decodeResult_sWrite = _RANDOM[9'h7][26];
        requestReg_bits_decodeResult_crossRead = _RANDOM[9'h7][27];
        requestReg_bits_decodeResult_crossWrite = _RANDOM[9'h7][28];
        requestReg_bits_decodeResult_maskUnit = _RANDOM[9'h7][29];
        requestReg_bits_decodeResult_special = _RANDOM[9'h7][30];
        requestReg_bits_decodeResult_saturate = _RANDOM[9'h7][31];
        requestReg_bits_decodeResult_vwmacc = _RANDOM[9'h8][0];
        requestReg_bits_decodeResult_readOnly = _RANDOM[9'h8][1];
        requestReg_bits_decodeResult_maskSource = _RANDOM[9'h8][2];
        requestReg_bits_decodeResult_maskDestination = _RANDOM[9'h8][3];
        requestReg_bits_decodeResult_maskLogic = _RANDOM[9'h8][4];
        requestReg_bits_decodeResult_uop = _RANDOM[9'h8][8:5];
        requestReg_bits_decodeResult_iota = _RANDOM[9'h8][9];
        requestReg_bits_decodeResult_mv = _RANDOM[9'h8][10];
        requestReg_bits_decodeResult_extend = _RANDOM[9'h8][11];
        requestReg_bits_decodeResult_unOrderWrite = _RANDOM[9'h8][12];
        requestReg_bits_decodeResult_compress = _RANDOM[9'h8][13];
        requestReg_bits_decodeResult_gather16 = _RANDOM[9'h8][14];
        requestReg_bits_decodeResult_gather = _RANDOM[9'h8][15];
        requestReg_bits_decodeResult_slid = _RANDOM[9'h8][16];
        requestReg_bits_decodeResult_targetRd = _RANDOM[9'h8][17];
        requestReg_bits_decodeResult_widenReduce = _RANDOM[9'h8][18];
        requestReg_bits_decodeResult_red = _RANDOM[9'h8][19];
        requestReg_bits_decodeResult_nr = _RANDOM[9'h8][20];
        requestReg_bits_decodeResult_itype = _RANDOM[9'h8][21];
        requestReg_bits_decodeResult_unsigned1 = _RANDOM[9'h8][22];
        requestReg_bits_decodeResult_unsigned0 = _RANDOM[9'h8][23];
        requestReg_bits_decodeResult_other = _RANDOM[9'h8][24];
        requestReg_bits_decodeResult_multiCycle = _RANDOM[9'h8][25];
        requestReg_bits_decodeResult_divider = _RANDOM[9'h8][26];
        requestReg_bits_decodeResult_multiplier = _RANDOM[9'h8][27];
        requestReg_bits_decodeResult_shift = _RANDOM[9'h8][28];
        requestReg_bits_decodeResult_adder = _RANDOM[9'h8][29];
        requestReg_bits_decodeResult_logic = _RANDOM[9'h8][30];
        requestReg_bits_instructionIndex = {_RANDOM[9'h8][31], _RANDOM[9'h9][1:0]};
        requestReg_bits_vdIsV0 = _RANDOM[9'h9][2];
        requestReg_bits_writeByte = _RANDOM[9'h9][14:3];
        slots_0_record_instructionIndex = _RANDOM[9'hA][18:16];
        slots_0_record_isLoadStore = _RANDOM[9'hA][19];
        slots_0_record_maskType = _RANDOM[9'hA][20];
        slots_0_state_wLast = _RANDOM[9'hA][21];
        slots_0_state_idle = _RANDOM[9'hA][22];
        slots_0_state_wMaskUnitLast = _RANDOM[9'hA][23];
        slots_0_state_wVRFWrite = _RANDOM[9'hA][24];
        slots_0_state_sCommit = _RANDOM[9'hA][25];
        slots_0_endTag_0 = _RANDOM[9'hA][26];
        slots_0_endTag_1 = _RANDOM[9'hA][27];
        slots_0_endTag_2 = _RANDOM[9'hA][28];
        slots_0_endTag_3 = _RANDOM[9'hA][29];
        slots_0_endTag_4 = _RANDOM[9'hA][30];
        slots_0_endTag_5 = _RANDOM[9'hA][31];
        slots_0_endTag_6 = _RANDOM[9'hB][0];
        slots_0_endTag_7 = _RANDOM[9'hB][1];
        slots_0_endTag_8 = _RANDOM[9'hB][2];
        slots_0_endTag_9 = _RANDOM[9'hB][3];
        slots_0_endTag_10 = _RANDOM[9'hB][4];
        slots_0_endTag_11 = _RANDOM[9'hB][5];
        slots_0_endTag_12 = _RANDOM[9'hB][6];
        slots_0_endTag_13 = _RANDOM[9'hB][7];
        slots_0_endTag_14 = _RANDOM[9'hB][8];
        slots_0_endTag_15 = _RANDOM[9'hB][9];
        slots_0_endTag_16 = _RANDOM[9'hB][10];
        slots_0_vxsat = _RANDOM[9'hB][11];
        slots_1_record_instructionIndex = _RANDOM[9'hB][14:12];
        slots_1_record_isLoadStore = _RANDOM[9'hB][15];
        slots_1_record_maskType = _RANDOM[9'hB][16];
        slots_1_state_wLast = _RANDOM[9'hB][17];
        slots_1_state_idle = _RANDOM[9'hB][18];
        slots_1_state_wMaskUnitLast = _RANDOM[9'hB][19];
        slots_1_state_wVRFWrite = _RANDOM[9'hB][20];
        slots_1_state_sCommit = _RANDOM[9'hB][21];
        slots_1_endTag_0 = _RANDOM[9'hB][22];
        slots_1_endTag_1 = _RANDOM[9'hB][23];
        slots_1_endTag_2 = _RANDOM[9'hB][24];
        slots_1_endTag_3 = _RANDOM[9'hB][25];
        slots_1_endTag_4 = _RANDOM[9'hB][26];
        slots_1_endTag_5 = _RANDOM[9'hB][27];
        slots_1_endTag_6 = _RANDOM[9'hB][28];
        slots_1_endTag_7 = _RANDOM[9'hB][29];
        slots_1_endTag_8 = _RANDOM[9'hB][30];
        slots_1_endTag_9 = _RANDOM[9'hB][31];
        slots_1_endTag_10 = _RANDOM[9'hC][0];
        slots_1_endTag_11 = _RANDOM[9'hC][1];
        slots_1_endTag_12 = _RANDOM[9'hC][2];
        slots_1_endTag_13 = _RANDOM[9'hC][3];
        slots_1_endTag_14 = _RANDOM[9'hC][4];
        slots_1_endTag_15 = _RANDOM[9'hC][5];
        slots_1_endTag_16 = _RANDOM[9'hC][6];
        slots_1_vxsat = _RANDOM[9'hC][7];
        slots_2_record_instructionIndex = _RANDOM[9'hC][10:8];
        slots_2_record_isLoadStore = _RANDOM[9'hC][11];
        slots_2_record_maskType = _RANDOM[9'hC][12];
        slots_2_state_wLast = _RANDOM[9'hC][13];
        slots_2_state_idle = _RANDOM[9'hC][14];
        slots_2_state_wMaskUnitLast = _RANDOM[9'hC][15];
        slots_2_state_wVRFWrite = _RANDOM[9'hC][16];
        slots_2_state_sCommit = _RANDOM[9'hC][17];
        slots_2_endTag_0 = _RANDOM[9'hC][18];
        slots_2_endTag_1 = _RANDOM[9'hC][19];
        slots_2_endTag_2 = _RANDOM[9'hC][20];
        slots_2_endTag_3 = _RANDOM[9'hC][21];
        slots_2_endTag_4 = _RANDOM[9'hC][22];
        slots_2_endTag_5 = _RANDOM[9'hC][23];
        slots_2_endTag_6 = _RANDOM[9'hC][24];
        slots_2_endTag_7 = _RANDOM[9'hC][25];
        slots_2_endTag_8 = _RANDOM[9'hC][26];
        slots_2_endTag_9 = _RANDOM[9'hC][27];
        slots_2_endTag_10 = _RANDOM[9'hC][28];
        slots_2_endTag_11 = _RANDOM[9'hC][29];
        slots_2_endTag_12 = _RANDOM[9'hC][30];
        slots_2_endTag_13 = _RANDOM[9'hC][31];
        slots_2_endTag_14 = _RANDOM[9'hD][0];
        slots_2_endTag_15 = _RANDOM[9'hD][1];
        slots_2_endTag_16 = _RANDOM[9'hD][2];
        slots_2_vxsat = _RANDOM[9'hD][3];
        slots_3_record_instructionIndex = _RANDOM[9'hD][6:4];
        slots_3_record_isLoadStore = _RANDOM[9'hD][7];
        slots_3_record_maskType = _RANDOM[9'hD][8];
        slots_3_state_wLast = _RANDOM[9'hD][9];
        slots_3_state_idle = _RANDOM[9'hD][10];
        slots_3_state_wMaskUnitLast = _RANDOM[9'hD][11];
        slots_3_state_wVRFWrite = _RANDOM[9'hD][12];
        slots_3_state_sCommit = _RANDOM[9'hD][13];
        slots_3_endTag_0 = _RANDOM[9'hD][14];
        slots_3_endTag_1 = _RANDOM[9'hD][15];
        slots_3_endTag_2 = _RANDOM[9'hD][16];
        slots_3_endTag_3 = _RANDOM[9'hD][17];
        slots_3_endTag_4 = _RANDOM[9'hD][18];
        slots_3_endTag_5 = _RANDOM[9'hD][19];
        slots_3_endTag_6 = _RANDOM[9'hD][20];
        slots_3_endTag_7 = _RANDOM[9'hD][21];
        slots_3_endTag_8 = _RANDOM[9'hD][22];
        slots_3_endTag_9 = _RANDOM[9'hD][23];
        slots_3_endTag_10 = _RANDOM[9'hD][24];
        slots_3_endTag_11 = _RANDOM[9'hD][25];
        slots_3_endTag_12 = _RANDOM[9'hD][26];
        slots_3_endTag_13 = _RANDOM[9'hD][27];
        slots_3_endTag_14 = _RANDOM[9'hD][28];
        slots_3_endTag_15 = _RANDOM[9'hD][29];
        slots_3_endTag_16 = _RANDOM[9'hD][30];
        slots_3_vxsat = _RANDOM[9'hD][31];
        slots_writeRD = _RANDOM[9'hE][0];
        slots_float = _RANDOM[9'hE][1];
        slots_vd = _RANDOM[9'hE][6:2];
        releasePipe_pipe_v = _RANDOM[9'hE][7];
        tokenCheck_counter = _RANDOM[9'hE][10:8];
        shifterReg_0_valid = _RANDOM[9'hE][11];
        shifterReg_0_bits_instructionIndex = _RANDOM[9'hE][14:12];
        shifterReg_0_bits_decodeResult_orderReduce = _RANDOM[9'hE][15];
        shifterReg_0_bits_decodeResult_floatMul = _RANDOM[9'hE][16];
        shifterReg_0_bits_decodeResult_fpExecutionType = _RANDOM[9'hE][18:17];
        shifterReg_0_bits_decodeResult_float = _RANDOM[9'hE][19];
        shifterReg_0_bits_decodeResult_specialSlot = _RANDOM[9'hE][20];
        shifterReg_0_bits_decodeResult_topUop = _RANDOM[9'hE][25:21];
        shifterReg_0_bits_decodeResult_popCount = _RANDOM[9'hE][26];
        shifterReg_0_bits_decodeResult_ffo = _RANDOM[9'hE][27];
        shifterReg_0_bits_decodeResult_average = _RANDOM[9'hE][28];
        shifterReg_0_bits_decodeResult_reverse = _RANDOM[9'hE][29];
        shifterReg_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'hE][30];
        shifterReg_0_bits_decodeResult_scheduler = _RANDOM[9'hE][31];
        shifterReg_0_bits_decodeResult_sReadVD = _RANDOM[9'hF][0];
        shifterReg_0_bits_decodeResult_vtype = _RANDOM[9'hF][1];
        shifterReg_0_bits_decodeResult_sWrite = _RANDOM[9'hF][2];
        shifterReg_0_bits_decodeResult_crossRead = _RANDOM[9'hF][3];
        shifterReg_0_bits_decodeResult_crossWrite = _RANDOM[9'hF][4];
        shifterReg_0_bits_decodeResult_maskUnit = _RANDOM[9'hF][5];
        shifterReg_0_bits_decodeResult_special = _RANDOM[9'hF][6];
        shifterReg_0_bits_decodeResult_saturate = _RANDOM[9'hF][7];
        shifterReg_0_bits_decodeResult_vwmacc = _RANDOM[9'hF][8];
        shifterReg_0_bits_decodeResult_readOnly = _RANDOM[9'hF][9];
        shifterReg_0_bits_decodeResult_maskSource = _RANDOM[9'hF][10];
        shifterReg_0_bits_decodeResult_maskDestination = _RANDOM[9'hF][11];
        shifterReg_0_bits_decodeResult_maskLogic = _RANDOM[9'hF][12];
        shifterReg_0_bits_decodeResult_uop = _RANDOM[9'hF][16:13];
        shifterReg_0_bits_decodeResult_iota = _RANDOM[9'hF][17];
        shifterReg_0_bits_decodeResult_mv = _RANDOM[9'hF][18];
        shifterReg_0_bits_decodeResult_extend = _RANDOM[9'hF][19];
        shifterReg_0_bits_decodeResult_unOrderWrite = _RANDOM[9'hF][20];
        shifterReg_0_bits_decodeResult_compress = _RANDOM[9'hF][21];
        shifterReg_0_bits_decodeResult_gather16 = _RANDOM[9'hF][22];
        shifterReg_0_bits_decodeResult_gather = _RANDOM[9'hF][23];
        shifterReg_0_bits_decodeResult_slid = _RANDOM[9'hF][24];
        shifterReg_0_bits_decodeResult_targetRd = _RANDOM[9'hF][25];
        shifterReg_0_bits_decodeResult_widenReduce = _RANDOM[9'hF][26];
        shifterReg_0_bits_decodeResult_red = _RANDOM[9'hF][27];
        shifterReg_0_bits_decodeResult_nr = _RANDOM[9'hF][28];
        shifterReg_0_bits_decodeResult_itype = _RANDOM[9'hF][29];
        shifterReg_0_bits_decodeResult_unsigned1 = _RANDOM[9'hF][30];
        shifterReg_0_bits_decodeResult_unsigned0 = _RANDOM[9'hF][31];
        shifterReg_0_bits_decodeResult_other = _RANDOM[9'h10][0];
        shifterReg_0_bits_decodeResult_multiCycle = _RANDOM[9'h10][1];
        shifterReg_0_bits_decodeResult_divider = _RANDOM[9'h10][2];
        shifterReg_0_bits_decodeResult_multiplier = _RANDOM[9'h10][3];
        shifterReg_0_bits_decodeResult_shift = _RANDOM[9'h10][4];
        shifterReg_0_bits_decodeResult_adder = _RANDOM[9'h10][5];
        shifterReg_0_bits_decodeResult_logic = _RANDOM[9'h10][6];
        shifterReg_0_bits_loadStore = _RANDOM[9'h10][7];
        shifterReg_0_bits_issueInst = _RANDOM[9'h10][8];
        shifterReg_0_bits_store = _RANDOM[9'h10][9];
        shifterReg_0_bits_special = _RANDOM[9'h10][10];
        shifterReg_0_bits_lsWholeReg = _RANDOM[9'h10][11];
        shifterReg_0_bits_vs1 = _RANDOM[9'h10][16:12];
        shifterReg_0_bits_vs2 = _RANDOM[9'h10][21:17];
        shifterReg_0_bits_vd = _RANDOM[9'h10][26:22];
        shifterReg_0_bits_loadStoreEEW = _RANDOM[9'h10][28:27];
        shifterReg_0_bits_mask = _RANDOM[9'h10][29];
        shifterReg_0_bits_segment = {_RANDOM[9'h10][31:30], _RANDOM[9'h11][0]};
        shifterReg_0_bits_readFromScalar = {_RANDOM[9'h11][31:1], _RANDOM[9'h12][0]};
        shifterReg_0_bits_csrInterface_vl = _RANDOM[9'h12][12:1];
        shifterReg_0_bits_csrInterface_vStart = _RANDOM[9'h12][24:13];
        shifterReg_0_bits_csrInterface_vlmul = _RANDOM[9'h12][27:25];
        shifterReg_0_bits_csrInterface_vSew = _RANDOM[9'h12][29:28];
        shifterReg_0_bits_csrInterface_vxrm = _RANDOM[9'h12][31:30];
        shifterReg_0_bits_csrInterface_vta = _RANDOM[9'h13][0];
        shifterReg_0_bits_csrInterface_vma = _RANDOM[9'h13][1];
        releasePipe_pipe_v_1 = _RANDOM[9'h13][2];
        tokenCheck_counter_1 = _RANDOM[9'h13][5:3];
        shifterReg_1_0_valid = _RANDOM[9'h13][6];
        shifterReg_1_0_bits_instructionIndex = _RANDOM[9'h13][9:7];
        shifterReg_1_0_bits_decodeResult_orderReduce = _RANDOM[9'h13][10];
        shifterReg_1_0_bits_decodeResult_floatMul = _RANDOM[9'h13][11];
        shifterReg_1_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h13][13:12];
        shifterReg_1_0_bits_decodeResult_float = _RANDOM[9'h13][14];
        shifterReg_1_0_bits_decodeResult_specialSlot = _RANDOM[9'h13][15];
        shifterReg_1_0_bits_decodeResult_topUop = _RANDOM[9'h13][20:16];
        shifterReg_1_0_bits_decodeResult_popCount = _RANDOM[9'h13][21];
        shifterReg_1_0_bits_decodeResult_ffo = _RANDOM[9'h13][22];
        shifterReg_1_0_bits_decodeResult_average = _RANDOM[9'h13][23];
        shifterReg_1_0_bits_decodeResult_reverse = _RANDOM[9'h13][24];
        shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h13][25];
        shifterReg_1_0_bits_decodeResult_scheduler = _RANDOM[9'h13][26];
        shifterReg_1_0_bits_decodeResult_sReadVD = _RANDOM[9'h13][27];
        shifterReg_1_0_bits_decodeResult_vtype = _RANDOM[9'h13][28];
        shifterReg_1_0_bits_decodeResult_sWrite = _RANDOM[9'h13][29];
        shifterReg_1_0_bits_decodeResult_crossRead = _RANDOM[9'h13][30];
        shifterReg_1_0_bits_decodeResult_crossWrite = _RANDOM[9'h13][31];
        shifterReg_1_0_bits_decodeResult_maskUnit = _RANDOM[9'h14][0];
        shifterReg_1_0_bits_decodeResult_special = _RANDOM[9'h14][1];
        shifterReg_1_0_bits_decodeResult_saturate = _RANDOM[9'h14][2];
        shifterReg_1_0_bits_decodeResult_vwmacc = _RANDOM[9'h14][3];
        shifterReg_1_0_bits_decodeResult_readOnly = _RANDOM[9'h14][4];
        shifterReg_1_0_bits_decodeResult_maskSource = _RANDOM[9'h14][5];
        shifterReg_1_0_bits_decodeResult_maskDestination = _RANDOM[9'h14][6];
        shifterReg_1_0_bits_decodeResult_maskLogic = _RANDOM[9'h14][7];
        shifterReg_1_0_bits_decodeResult_uop = _RANDOM[9'h14][11:8];
        shifterReg_1_0_bits_decodeResult_iota = _RANDOM[9'h14][12];
        shifterReg_1_0_bits_decodeResult_mv = _RANDOM[9'h14][13];
        shifterReg_1_0_bits_decodeResult_extend = _RANDOM[9'h14][14];
        shifterReg_1_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h14][15];
        shifterReg_1_0_bits_decodeResult_compress = _RANDOM[9'h14][16];
        shifterReg_1_0_bits_decodeResult_gather16 = _RANDOM[9'h14][17];
        shifterReg_1_0_bits_decodeResult_gather = _RANDOM[9'h14][18];
        shifterReg_1_0_bits_decodeResult_slid = _RANDOM[9'h14][19];
        shifterReg_1_0_bits_decodeResult_targetRd = _RANDOM[9'h14][20];
        shifterReg_1_0_bits_decodeResult_widenReduce = _RANDOM[9'h14][21];
        shifterReg_1_0_bits_decodeResult_red = _RANDOM[9'h14][22];
        shifterReg_1_0_bits_decodeResult_nr = _RANDOM[9'h14][23];
        shifterReg_1_0_bits_decodeResult_itype = _RANDOM[9'h14][24];
        shifterReg_1_0_bits_decodeResult_unsigned1 = _RANDOM[9'h14][25];
        shifterReg_1_0_bits_decodeResult_unsigned0 = _RANDOM[9'h14][26];
        shifterReg_1_0_bits_decodeResult_other = _RANDOM[9'h14][27];
        shifterReg_1_0_bits_decodeResult_multiCycle = _RANDOM[9'h14][28];
        shifterReg_1_0_bits_decodeResult_divider = _RANDOM[9'h14][29];
        shifterReg_1_0_bits_decodeResult_multiplier = _RANDOM[9'h14][30];
        shifterReg_1_0_bits_decodeResult_shift = _RANDOM[9'h14][31];
        shifterReg_1_0_bits_decodeResult_adder = _RANDOM[9'h15][0];
        shifterReg_1_0_bits_decodeResult_logic = _RANDOM[9'h15][1];
        shifterReg_1_0_bits_loadStore = _RANDOM[9'h15][2];
        shifterReg_1_0_bits_issueInst = _RANDOM[9'h15][3];
        shifterReg_1_0_bits_store = _RANDOM[9'h15][4];
        shifterReg_1_0_bits_special = _RANDOM[9'h15][5];
        shifterReg_1_0_bits_lsWholeReg = _RANDOM[9'h15][6];
        shifterReg_1_0_bits_vs1 = _RANDOM[9'h15][11:7];
        shifterReg_1_0_bits_vs2 = _RANDOM[9'h15][16:12];
        shifterReg_1_0_bits_vd = _RANDOM[9'h15][21:17];
        shifterReg_1_0_bits_loadStoreEEW = _RANDOM[9'h15][23:22];
        shifterReg_1_0_bits_mask = _RANDOM[9'h15][24];
        shifterReg_1_0_bits_segment = _RANDOM[9'h15][27:25];
        shifterReg_1_0_bits_readFromScalar = {_RANDOM[9'h15][31:28], _RANDOM[9'h16][27:0]};
        shifterReg_1_0_bits_csrInterface_vl = {_RANDOM[9'h16][31:28], _RANDOM[9'h17][7:0]};
        shifterReg_1_0_bits_csrInterface_vStart = _RANDOM[9'h17][19:8];
        shifterReg_1_0_bits_csrInterface_vlmul = _RANDOM[9'h17][22:20];
        shifterReg_1_0_bits_csrInterface_vSew = _RANDOM[9'h17][24:23];
        shifterReg_1_0_bits_csrInterface_vxrm = _RANDOM[9'h17][26:25];
        shifterReg_1_0_bits_csrInterface_vta = _RANDOM[9'h17][27];
        shifterReg_1_0_bits_csrInterface_vma = _RANDOM[9'h17][28];
        releasePipe_pipe_v_2 = _RANDOM[9'h17][29];
        tokenCheck_counter_2 = {_RANDOM[9'h17][31:30], _RANDOM[9'h18][0]};
        shifterReg_2_0_valid = _RANDOM[9'h18][1];
        shifterReg_2_0_bits_instructionIndex = _RANDOM[9'h18][4:2];
        shifterReg_2_0_bits_decodeResult_orderReduce = _RANDOM[9'h18][5];
        shifterReg_2_0_bits_decodeResult_floatMul = _RANDOM[9'h18][6];
        shifterReg_2_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h18][8:7];
        shifterReg_2_0_bits_decodeResult_float = _RANDOM[9'h18][9];
        shifterReg_2_0_bits_decodeResult_specialSlot = _RANDOM[9'h18][10];
        shifterReg_2_0_bits_decodeResult_topUop = _RANDOM[9'h18][15:11];
        shifterReg_2_0_bits_decodeResult_popCount = _RANDOM[9'h18][16];
        shifterReg_2_0_bits_decodeResult_ffo = _RANDOM[9'h18][17];
        shifterReg_2_0_bits_decodeResult_average = _RANDOM[9'h18][18];
        shifterReg_2_0_bits_decodeResult_reverse = _RANDOM[9'h18][19];
        shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h18][20];
        shifterReg_2_0_bits_decodeResult_scheduler = _RANDOM[9'h18][21];
        shifterReg_2_0_bits_decodeResult_sReadVD = _RANDOM[9'h18][22];
        shifterReg_2_0_bits_decodeResult_vtype = _RANDOM[9'h18][23];
        shifterReg_2_0_bits_decodeResult_sWrite = _RANDOM[9'h18][24];
        shifterReg_2_0_bits_decodeResult_crossRead = _RANDOM[9'h18][25];
        shifterReg_2_0_bits_decodeResult_crossWrite = _RANDOM[9'h18][26];
        shifterReg_2_0_bits_decodeResult_maskUnit = _RANDOM[9'h18][27];
        shifterReg_2_0_bits_decodeResult_special = _RANDOM[9'h18][28];
        shifterReg_2_0_bits_decodeResult_saturate = _RANDOM[9'h18][29];
        shifterReg_2_0_bits_decodeResult_vwmacc = _RANDOM[9'h18][30];
        shifterReg_2_0_bits_decodeResult_readOnly = _RANDOM[9'h18][31];
        shifterReg_2_0_bits_decodeResult_maskSource = _RANDOM[9'h19][0];
        shifterReg_2_0_bits_decodeResult_maskDestination = _RANDOM[9'h19][1];
        shifterReg_2_0_bits_decodeResult_maskLogic = _RANDOM[9'h19][2];
        shifterReg_2_0_bits_decodeResult_uop = _RANDOM[9'h19][6:3];
        shifterReg_2_0_bits_decodeResult_iota = _RANDOM[9'h19][7];
        shifterReg_2_0_bits_decodeResult_mv = _RANDOM[9'h19][8];
        shifterReg_2_0_bits_decodeResult_extend = _RANDOM[9'h19][9];
        shifterReg_2_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h19][10];
        shifterReg_2_0_bits_decodeResult_compress = _RANDOM[9'h19][11];
        shifterReg_2_0_bits_decodeResult_gather16 = _RANDOM[9'h19][12];
        shifterReg_2_0_bits_decodeResult_gather = _RANDOM[9'h19][13];
        shifterReg_2_0_bits_decodeResult_slid = _RANDOM[9'h19][14];
        shifterReg_2_0_bits_decodeResult_targetRd = _RANDOM[9'h19][15];
        shifterReg_2_0_bits_decodeResult_widenReduce = _RANDOM[9'h19][16];
        shifterReg_2_0_bits_decodeResult_red = _RANDOM[9'h19][17];
        shifterReg_2_0_bits_decodeResult_nr = _RANDOM[9'h19][18];
        shifterReg_2_0_bits_decodeResult_itype = _RANDOM[9'h19][19];
        shifterReg_2_0_bits_decodeResult_unsigned1 = _RANDOM[9'h19][20];
        shifterReg_2_0_bits_decodeResult_unsigned0 = _RANDOM[9'h19][21];
        shifterReg_2_0_bits_decodeResult_other = _RANDOM[9'h19][22];
        shifterReg_2_0_bits_decodeResult_multiCycle = _RANDOM[9'h19][23];
        shifterReg_2_0_bits_decodeResult_divider = _RANDOM[9'h19][24];
        shifterReg_2_0_bits_decodeResult_multiplier = _RANDOM[9'h19][25];
        shifterReg_2_0_bits_decodeResult_shift = _RANDOM[9'h19][26];
        shifterReg_2_0_bits_decodeResult_adder = _RANDOM[9'h19][27];
        shifterReg_2_0_bits_decodeResult_logic = _RANDOM[9'h19][28];
        shifterReg_2_0_bits_loadStore = _RANDOM[9'h19][29];
        shifterReg_2_0_bits_issueInst = _RANDOM[9'h19][30];
        shifterReg_2_0_bits_store = _RANDOM[9'h19][31];
        shifterReg_2_0_bits_special = _RANDOM[9'h1A][0];
        shifterReg_2_0_bits_lsWholeReg = _RANDOM[9'h1A][1];
        shifterReg_2_0_bits_vs1 = _RANDOM[9'h1A][6:2];
        shifterReg_2_0_bits_vs2 = _RANDOM[9'h1A][11:7];
        shifterReg_2_0_bits_vd = _RANDOM[9'h1A][16:12];
        shifterReg_2_0_bits_loadStoreEEW = _RANDOM[9'h1A][18:17];
        shifterReg_2_0_bits_mask = _RANDOM[9'h1A][19];
        shifterReg_2_0_bits_segment = _RANDOM[9'h1A][22:20];
        shifterReg_2_0_bits_readFromScalar = {_RANDOM[9'h1A][31:23], _RANDOM[9'h1B][22:0]};
        shifterReg_2_0_bits_csrInterface_vl = {_RANDOM[9'h1B][31:23], _RANDOM[9'h1C][2:0]};
        shifterReg_2_0_bits_csrInterface_vStart = _RANDOM[9'h1C][14:3];
        shifterReg_2_0_bits_csrInterface_vlmul = _RANDOM[9'h1C][17:15];
        shifterReg_2_0_bits_csrInterface_vSew = _RANDOM[9'h1C][19:18];
        shifterReg_2_0_bits_csrInterface_vxrm = _RANDOM[9'h1C][21:20];
        shifterReg_2_0_bits_csrInterface_vta = _RANDOM[9'h1C][22];
        shifterReg_2_0_bits_csrInterface_vma = _RANDOM[9'h1C][23];
        releasePipe_pipe_v_3 = _RANDOM[9'h1C][24];
        tokenCheck_counter_3 = _RANDOM[9'h1C][27:25];
        shifterReg_3_0_valid = _RANDOM[9'h1C][28];
        shifterReg_3_0_bits_instructionIndex = _RANDOM[9'h1C][31:29];
        shifterReg_3_0_bits_decodeResult_orderReduce = _RANDOM[9'h1D][0];
        shifterReg_3_0_bits_decodeResult_floatMul = _RANDOM[9'h1D][1];
        shifterReg_3_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h1D][3:2];
        shifterReg_3_0_bits_decodeResult_float = _RANDOM[9'h1D][4];
        shifterReg_3_0_bits_decodeResult_specialSlot = _RANDOM[9'h1D][5];
        shifterReg_3_0_bits_decodeResult_topUop = _RANDOM[9'h1D][10:6];
        shifterReg_3_0_bits_decodeResult_popCount = _RANDOM[9'h1D][11];
        shifterReg_3_0_bits_decodeResult_ffo = _RANDOM[9'h1D][12];
        shifterReg_3_0_bits_decodeResult_average = _RANDOM[9'h1D][13];
        shifterReg_3_0_bits_decodeResult_reverse = _RANDOM[9'h1D][14];
        shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h1D][15];
        shifterReg_3_0_bits_decodeResult_scheduler = _RANDOM[9'h1D][16];
        shifterReg_3_0_bits_decodeResult_sReadVD = _RANDOM[9'h1D][17];
        shifterReg_3_0_bits_decodeResult_vtype = _RANDOM[9'h1D][18];
        shifterReg_3_0_bits_decodeResult_sWrite = _RANDOM[9'h1D][19];
        shifterReg_3_0_bits_decodeResult_crossRead = _RANDOM[9'h1D][20];
        shifterReg_3_0_bits_decodeResult_crossWrite = _RANDOM[9'h1D][21];
        shifterReg_3_0_bits_decodeResult_maskUnit = _RANDOM[9'h1D][22];
        shifterReg_3_0_bits_decodeResult_special = _RANDOM[9'h1D][23];
        shifterReg_3_0_bits_decodeResult_saturate = _RANDOM[9'h1D][24];
        shifterReg_3_0_bits_decodeResult_vwmacc = _RANDOM[9'h1D][25];
        shifterReg_3_0_bits_decodeResult_readOnly = _RANDOM[9'h1D][26];
        shifterReg_3_0_bits_decodeResult_maskSource = _RANDOM[9'h1D][27];
        shifterReg_3_0_bits_decodeResult_maskDestination = _RANDOM[9'h1D][28];
        shifterReg_3_0_bits_decodeResult_maskLogic = _RANDOM[9'h1D][29];
        shifterReg_3_0_bits_decodeResult_uop = {_RANDOM[9'h1D][31:30], _RANDOM[9'h1E][1:0]};
        shifterReg_3_0_bits_decodeResult_iota = _RANDOM[9'h1E][2];
        shifterReg_3_0_bits_decodeResult_mv = _RANDOM[9'h1E][3];
        shifterReg_3_0_bits_decodeResult_extend = _RANDOM[9'h1E][4];
        shifterReg_3_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h1E][5];
        shifterReg_3_0_bits_decodeResult_compress = _RANDOM[9'h1E][6];
        shifterReg_3_0_bits_decodeResult_gather16 = _RANDOM[9'h1E][7];
        shifterReg_3_0_bits_decodeResult_gather = _RANDOM[9'h1E][8];
        shifterReg_3_0_bits_decodeResult_slid = _RANDOM[9'h1E][9];
        shifterReg_3_0_bits_decodeResult_targetRd = _RANDOM[9'h1E][10];
        shifterReg_3_0_bits_decodeResult_widenReduce = _RANDOM[9'h1E][11];
        shifterReg_3_0_bits_decodeResult_red = _RANDOM[9'h1E][12];
        shifterReg_3_0_bits_decodeResult_nr = _RANDOM[9'h1E][13];
        shifterReg_3_0_bits_decodeResult_itype = _RANDOM[9'h1E][14];
        shifterReg_3_0_bits_decodeResult_unsigned1 = _RANDOM[9'h1E][15];
        shifterReg_3_0_bits_decodeResult_unsigned0 = _RANDOM[9'h1E][16];
        shifterReg_3_0_bits_decodeResult_other = _RANDOM[9'h1E][17];
        shifterReg_3_0_bits_decodeResult_multiCycle = _RANDOM[9'h1E][18];
        shifterReg_3_0_bits_decodeResult_divider = _RANDOM[9'h1E][19];
        shifterReg_3_0_bits_decodeResult_multiplier = _RANDOM[9'h1E][20];
        shifterReg_3_0_bits_decodeResult_shift = _RANDOM[9'h1E][21];
        shifterReg_3_0_bits_decodeResult_adder = _RANDOM[9'h1E][22];
        shifterReg_3_0_bits_decodeResult_logic = _RANDOM[9'h1E][23];
        shifterReg_3_0_bits_loadStore = _RANDOM[9'h1E][24];
        shifterReg_3_0_bits_issueInst = _RANDOM[9'h1E][25];
        shifterReg_3_0_bits_store = _RANDOM[9'h1E][26];
        shifterReg_3_0_bits_special = _RANDOM[9'h1E][27];
        shifterReg_3_0_bits_lsWholeReg = _RANDOM[9'h1E][28];
        shifterReg_3_0_bits_vs1 = {_RANDOM[9'h1E][31:29], _RANDOM[9'h1F][1:0]};
        shifterReg_3_0_bits_vs2 = _RANDOM[9'h1F][6:2];
        shifterReg_3_0_bits_vd = _RANDOM[9'h1F][11:7];
        shifterReg_3_0_bits_loadStoreEEW = _RANDOM[9'h1F][13:12];
        shifterReg_3_0_bits_mask = _RANDOM[9'h1F][14];
        shifterReg_3_0_bits_segment = _RANDOM[9'h1F][17:15];
        shifterReg_3_0_bits_readFromScalar = {_RANDOM[9'h1F][31:18], _RANDOM[9'h20][17:0]};
        shifterReg_3_0_bits_csrInterface_vl = _RANDOM[9'h20][29:18];
        shifterReg_3_0_bits_csrInterface_vStart = {_RANDOM[9'h20][31:30], _RANDOM[9'h21][9:0]};
        shifterReg_3_0_bits_csrInterface_vlmul = _RANDOM[9'h21][12:10];
        shifterReg_3_0_bits_csrInterface_vSew = _RANDOM[9'h21][14:13];
        shifterReg_3_0_bits_csrInterface_vxrm = _RANDOM[9'h21][16:15];
        shifterReg_3_0_bits_csrInterface_vta = _RANDOM[9'h21][17];
        shifterReg_3_0_bits_csrInterface_vma = _RANDOM[9'h21][18];
        releasePipe_pipe_v_4 = _RANDOM[9'h21][19];
        tokenCheck_counter_4 = _RANDOM[9'h21][22:20];
        shifterReg_4_0_valid = _RANDOM[9'h21][23];
        shifterReg_4_0_bits_instructionIndex = _RANDOM[9'h21][26:24];
        shifterReg_4_0_bits_decodeResult_orderReduce = _RANDOM[9'h21][27];
        shifterReg_4_0_bits_decodeResult_floatMul = _RANDOM[9'h21][28];
        shifterReg_4_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h21][30:29];
        shifterReg_4_0_bits_decodeResult_float = _RANDOM[9'h21][31];
        shifterReg_4_0_bits_decodeResult_specialSlot = _RANDOM[9'h22][0];
        shifterReg_4_0_bits_decodeResult_topUop = _RANDOM[9'h22][5:1];
        shifterReg_4_0_bits_decodeResult_popCount = _RANDOM[9'h22][6];
        shifterReg_4_0_bits_decodeResult_ffo = _RANDOM[9'h22][7];
        shifterReg_4_0_bits_decodeResult_average = _RANDOM[9'h22][8];
        shifterReg_4_0_bits_decodeResult_reverse = _RANDOM[9'h22][9];
        shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h22][10];
        shifterReg_4_0_bits_decodeResult_scheduler = _RANDOM[9'h22][11];
        shifterReg_4_0_bits_decodeResult_sReadVD = _RANDOM[9'h22][12];
        shifterReg_4_0_bits_decodeResult_vtype = _RANDOM[9'h22][13];
        shifterReg_4_0_bits_decodeResult_sWrite = _RANDOM[9'h22][14];
        shifterReg_4_0_bits_decodeResult_crossRead = _RANDOM[9'h22][15];
        shifterReg_4_0_bits_decodeResult_crossWrite = _RANDOM[9'h22][16];
        shifterReg_4_0_bits_decodeResult_maskUnit = _RANDOM[9'h22][17];
        shifterReg_4_0_bits_decodeResult_special = _RANDOM[9'h22][18];
        shifterReg_4_0_bits_decodeResult_saturate = _RANDOM[9'h22][19];
        shifterReg_4_0_bits_decodeResult_vwmacc = _RANDOM[9'h22][20];
        shifterReg_4_0_bits_decodeResult_readOnly = _RANDOM[9'h22][21];
        shifterReg_4_0_bits_decodeResult_maskSource = _RANDOM[9'h22][22];
        shifterReg_4_0_bits_decodeResult_maskDestination = _RANDOM[9'h22][23];
        shifterReg_4_0_bits_decodeResult_maskLogic = _RANDOM[9'h22][24];
        shifterReg_4_0_bits_decodeResult_uop = _RANDOM[9'h22][28:25];
        shifterReg_4_0_bits_decodeResult_iota = _RANDOM[9'h22][29];
        shifterReg_4_0_bits_decodeResult_mv = _RANDOM[9'h22][30];
        shifterReg_4_0_bits_decodeResult_extend = _RANDOM[9'h22][31];
        shifterReg_4_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h23][0];
        shifterReg_4_0_bits_decodeResult_compress = _RANDOM[9'h23][1];
        shifterReg_4_0_bits_decodeResult_gather16 = _RANDOM[9'h23][2];
        shifterReg_4_0_bits_decodeResult_gather = _RANDOM[9'h23][3];
        shifterReg_4_0_bits_decodeResult_slid = _RANDOM[9'h23][4];
        shifterReg_4_0_bits_decodeResult_targetRd = _RANDOM[9'h23][5];
        shifterReg_4_0_bits_decodeResult_widenReduce = _RANDOM[9'h23][6];
        shifterReg_4_0_bits_decodeResult_red = _RANDOM[9'h23][7];
        shifterReg_4_0_bits_decodeResult_nr = _RANDOM[9'h23][8];
        shifterReg_4_0_bits_decodeResult_itype = _RANDOM[9'h23][9];
        shifterReg_4_0_bits_decodeResult_unsigned1 = _RANDOM[9'h23][10];
        shifterReg_4_0_bits_decodeResult_unsigned0 = _RANDOM[9'h23][11];
        shifterReg_4_0_bits_decodeResult_other = _RANDOM[9'h23][12];
        shifterReg_4_0_bits_decodeResult_multiCycle = _RANDOM[9'h23][13];
        shifterReg_4_0_bits_decodeResult_divider = _RANDOM[9'h23][14];
        shifterReg_4_0_bits_decodeResult_multiplier = _RANDOM[9'h23][15];
        shifterReg_4_0_bits_decodeResult_shift = _RANDOM[9'h23][16];
        shifterReg_4_0_bits_decodeResult_adder = _RANDOM[9'h23][17];
        shifterReg_4_0_bits_decodeResult_logic = _RANDOM[9'h23][18];
        shifterReg_4_0_bits_loadStore = _RANDOM[9'h23][19];
        shifterReg_4_0_bits_issueInst = _RANDOM[9'h23][20];
        shifterReg_4_0_bits_store = _RANDOM[9'h23][21];
        shifterReg_4_0_bits_special = _RANDOM[9'h23][22];
        shifterReg_4_0_bits_lsWholeReg = _RANDOM[9'h23][23];
        shifterReg_4_0_bits_vs1 = _RANDOM[9'h23][28:24];
        shifterReg_4_0_bits_vs2 = {_RANDOM[9'h23][31:29], _RANDOM[9'h24][1:0]};
        shifterReg_4_0_bits_vd = _RANDOM[9'h24][6:2];
        shifterReg_4_0_bits_loadStoreEEW = _RANDOM[9'h24][8:7];
        shifterReg_4_0_bits_mask = _RANDOM[9'h24][9];
        shifterReg_4_0_bits_segment = _RANDOM[9'h24][12:10];
        shifterReg_4_0_bits_readFromScalar = {_RANDOM[9'h24][31:13], _RANDOM[9'h25][12:0]};
        shifterReg_4_0_bits_csrInterface_vl = _RANDOM[9'h25][24:13];
        shifterReg_4_0_bits_csrInterface_vStart = {_RANDOM[9'h25][31:25], _RANDOM[9'h26][4:0]};
        shifterReg_4_0_bits_csrInterface_vlmul = _RANDOM[9'h26][7:5];
        shifterReg_4_0_bits_csrInterface_vSew = _RANDOM[9'h26][9:8];
        shifterReg_4_0_bits_csrInterface_vxrm = _RANDOM[9'h26][11:10];
        shifterReg_4_0_bits_csrInterface_vta = _RANDOM[9'h26][12];
        shifterReg_4_0_bits_csrInterface_vma = _RANDOM[9'h26][13];
        releasePipe_pipe_v_5 = _RANDOM[9'h26][14];
        tokenCheck_counter_5 = _RANDOM[9'h26][17:15];
        shifterReg_5_0_valid = _RANDOM[9'h26][18];
        shifterReg_5_0_bits_instructionIndex = _RANDOM[9'h26][21:19];
        shifterReg_5_0_bits_decodeResult_orderReduce = _RANDOM[9'h26][22];
        shifterReg_5_0_bits_decodeResult_floatMul = _RANDOM[9'h26][23];
        shifterReg_5_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h26][25:24];
        shifterReg_5_0_bits_decodeResult_float = _RANDOM[9'h26][26];
        shifterReg_5_0_bits_decodeResult_specialSlot = _RANDOM[9'h26][27];
        shifterReg_5_0_bits_decodeResult_topUop = {_RANDOM[9'h26][31:28], _RANDOM[9'h27][0]};
        shifterReg_5_0_bits_decodeResult_popCount = _RANDOM[9'h27][1];
        shifterReg_5_0_bits_decodeResult_ffo = _RANDOM[9'h27][2];
        shifterReg_5_0_bits_decodeResult_average = _RANDOM[9'h27][3];
        shifterReg_5_0_bits_decodeResult_reverse = _RANDOM[9'h27][4];
        shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h27][5];
        shifterReg_5_0_bits_decodeResult_scheduler = _RANDOM[9'h27][6];
        shifterReg_5_0_bits_decodeResult_sReadVD = _RANDOM[9'h27][7];
        shifterReg_5_0_bits_decodeResult_vtype = _RANDOM[9'h27][8];
        shifterReg_5_0_bits_decodeResult_sWrite = _RANDOM[9'h27][9];
        shifterReg_5_0_bits_decodeResult_crossRead = _RANDOM[9'h27][10];
        shifterReg_5_0_bits_decodeResult_crossWrite = _RANDOM[9'h27][11];
        shifterReg_5_0_bits_decodeResult_maskUnit = _RANDOM[9'h27][12];
        shifterReg_5_0_bits_decodeResult_special = _RANDOM[9'h27][13];
        shifterReg_5_0_bits_decodeResult_saturate = _RANDOM[9'h27][14];
        shifterReg_5_0_bits_decodeResult_vwmacc = _RANDOM[9'h27][15];
        shifterReg_5_0_bits_decodeResult_readOnly = _RANDOM[9'h27][16];
        shifterReg_5_0_bits_decodeResult_maskSource = _RANDOM[9'h27][17];
        shifterReg_5_0_bits_decodeResult_maskDestination = _RANDOM[9'h27][18];
        shifterReg_5_0_bits_decodeResult_maskLogic = _RANDOM[9'h27][19];
        shifterReg_5_0_bits_decodeResult_uop = _RANDOM[9'h27][23:20];
        shifterReg_5_0_bits_decodeResult_iota = _RANDOM[9'h27][24];
        shifterReg_5_0_bits_decodeResult_mv = _RANDOM[9'h27][25];
        shifterReg_5_0_bits_decodeResult_extend = _RANDOM[9'h27][26];
        shifterReg_5_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h27][27];
        shifterReg_5_0_bits_decodeResult_compress = _RANDOM[9'h27][28];
        shifterReg_5_0_bits_decodeResult_gather16 = _RANDOM[9'h27][29];
        shifterReg_5_0_bits_decodeResult_gather = _RANDOM[9'h27][30];
        shifterReg_5_0_bits_decodeResult_slid = _RANDOM[9'h27][31];
        shifterReg_5_0_bits_decodeResult_targetRd = _RANDOM[9'h28][0];
        shifterReg_5_0_bits_decodeResult_widenReduce = _RANDOM[9'h28][1];
        shifterReg_5_0_bits_decodeResult_red = _RANDOM[9'h28][2];
        shifterReg_5_0_bits_decodeResult_nr = _RANDOM[9'h28][3];
        shifterReg_5_0_bits_decodeResult_itype = _RANDOM[9'h28][4];
        shifterReg_5_0_bits_decodeResult_unsigned1 = _RANDOM[9'h28][5];
        shifterReg_5_0_bits_decodeResult_unsigned0 = _RANDOM[9'h28][6];
        shifterReg_5_0_bits_decodeResult_other = _RANDOM[9'h28][7];
        shifterReg_5_0_bits_decodeResult_multiCycle = _RANDOM[9'h28][8];
        shifterReg_5_0_bits_decodeResult_divider = _RANDOM[9'h28][9];
        shifterReg_5_0_bits_decodeResult_multiplier = _RANDOM[9'h28][10];
        shifterReg_5_0_bits_decodeResult_shift = _RANDOM[9'h28][11];
        shifterReg_5_0_bits_decodeResult_adder = _RANDOM[9'h28][12];
        shifterReg_5_0_bits_decodeResult_logic = _RANDOM[9'h28][13];
        shifterReg_5_0_bits_loadStore = _RANDOM[9'h28][14];
        shifterReg_5_0_bits_issueInst = _RANDOM[9'h28][15];
        shifterReg_5_0_bits_store = _RANDOM[9'h28][16];
        shifterReg_5_0_bits_special = _RANDOM[9'h28][17];
        shifterReg_5_0_bits_lsWholeReg = _RANDOM[9'h28][18];
        shifterReg_5_0_bits_vs1 = _RANDOM[9'h28][23:19];
        shifterReg_5_0_bits_vs2 = _RANDOM[9'h28][28:24];
        shifterReg_5_0_bits_vd = {_RANDOM[9'h28][31:29], _RANDOM[9'h29][1:0]};
        shifterReg_5_0_bits_loadStoreEEW = _RANDOM[9'h29][3:2];
        shifterReg_5_0_bits_mask = _RANDOM[9'h29][4];
        shifterReg_5_0_bits_segment = _RANDOM[9'h29][7:5];
        shifterReg_5_0_bits_readFromScalar = {_RANDOM[9'h29][31:8], _RANDOM[9'h2A][7:0]};
        shifterReg_5_0_bits_csrInterface_vl = _RANDOM[9'h2A][19:8];
        shifterReg_5_0_bits_csrInterface_vStart = _RANDOM[9'h2A][31:20];
        shifterReg_5_0_bits_csrInterface_vlmul = _RANDOM[9'h2B][2:0];
        shifterReg_5_0_bits_csrInterface_vSew = _RANDOM[9'h2B][4:3];
        shifterReg_5_0_bits_csrInterface_vxrm = _RANDOM[9'h2B][6:5];
        shifterReg_5_0_bits_csrInterface_vta = _RANDOM[9'h2B][7];
        shifterReg_5_0_bits_csrInterface_vma = _RANDOM[9'h2B][8];
        releasePipe_pipe_v_6 = _RANDOM[9'h2B][9];
        tokenCheck_counter_6 = _RANDOM[9'h2B][12:10];
        shifterReg_6_0_valid = _RANDOM[9'h2B][13];
        shifterReg_6_0_bits_instructionIndex = _RANDOM[9'h2B][16:14];
        shifterReg_6_0_bits_decodeResult_orderReduce = _RANDOM[9'h2B][17];
        shifterReg_6_0_bits_decodeResult_floatMul = _RANDOM[9'h2B][18];
        shifterReg_6_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h2B][20:19];
        shifterReg_6_0_bits_decodeResult_float = _RANDOM[9'h2B][21];
        shifterReg_6_0_bits_decodeResult_specialSlot = _RANDOM[9'h2B][22];
        shifterReg_6_0_bits_decodeResult_topUop = _RANDOM[9'h2B][27:23];
        shifterReg_6_0_bits_decodeResult_popCount = _RANDOM[9'h2B][28];
        shifterReg_6_0_bits_decodeResult_ffo = _RANDOM[9'h2B][29];
        shifterReg_6_0_bits_decodeResult_average = _RANDOM[9'h2B][30];
        shifterReg_6_0_bits_decodeResult_reverse = _RANDOM[9'h2B][31];
        shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h2C][0];
        shifterReg_6_0_bits_decodeResult_scheduler = _RANDOM[9'h2C][1];
        shifterReg_6_0_bits_decodeResult_sReadVD = _RANDOM[9'h2C][2];
        shifterReg_6_0_bits_decodeResult_vtype = _RANDOM[9'h2C][3];
        shifterReg_6_0_bits_decodeResult_sWrite = _RANDOM[9'h2C][4];
        shifterReg_6_0_bits_decodeResult_crossRead = _RANDOM[9'h2C][5];
        shifterReg_6_0_bits_decodeResult_crossWrite = _RANDOM[9'h2C][6];
        shifterReg_6_0_bits_decodeResult_maskUnit = _RANDOM[9'h2C][7];
        shifterReg_6_0_bits_decodeResult_special = _RANDOM[9'h2C][8];
        shifterReg_6_0_bits_decodeResult_saturate = _RANDOM[9'h2C][9];
        shifterReg_6_0_bits_decodeResult_vwmacc = _RANDOM[9'h2C][10];
        shifterReg_6_0_bits_decodeResult_readOnly = _RANDOM[9'h2C][11];
        shifterReg_6_0_bits_decodeResult_maskSource = _RANDOM[9'h2C][12];
        shifterReg_6_0_bits_decodeResult_maskDestination = _RANDOM[9'h2C][13];
        shifterReg_6_0_bits_decodeResult_maskLogic = _RANDOM[9'h2C][14];
        shifterReg_6_0_bits_decodeResult_uop = _RANDOM[9'h2C][18:15];
        shifterReg_6_0_bits_decodeResult_iota = _RANDOM[9'h2C][19];
        shifterReg_6_0_bits_decodeResult_mv = _RANDOM[9'h2C][20];
        shifterReg_6_0_bits_decodeResult_extend = _RANDOM[9'h2C][21];
        shifterReg_6_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h2C][22];
        shifterReg_6_0_bits_decodeResult_compress = _RANDOM[9'h2C][23];
        shifterReg_6_0_bits_decodeResult_gather16 = _RANDOM[9'h2C][24];
        shifterReg_6_0_bits_decodeResult_gather = _RANDOM[9'h2C][25];
        shifterReg_6_0_bits_decodeResult_slid = _RANDOM[9'h2C][26];
        shifterReg_6_0_bits_decodeResult_targetRd = _RANDOM[9'h2C][27];
        shifterReg_6_0_bits_decodeResult_widenReduce = _RANDOM[9'h2C][28];
        shifterReg_6_0_bits_decodeResult_red = _RANDOM[9'h2C][29];
        shifterReg_6_0_bits_decodeResult_nr = _RANDOM[9'h2C][30];
        shifterReg_6_0_bits_decodeResult_itype = _RANDOM[9'h2C][31];
        shifterReg_6_0_bits_decodeResult_unsigned1 = _RANDOM[9'h2D][0];
        shifterReg_6_0_bits_decodeResult_unsigned0 = _RANDOM[9'h2D][1];
        shifterReg_6_0_bits_decodeResult_other = _RANDOM[9'h2D][2];
        shifterReg_6_0_bits_decodeResult_multiCycle = _RANDOM[9'h2D][3];
        shifterReg_6_0_bits_decodeResult_divider = _RANDOM[9'h2D][4];
        shifterReg_6_0_bits_decodeResult_multiplier = _RANDOM[9'h2D][5];
        shifterReg_6_0_bits_decodeResult_shift = _RANDOM[9'h2D][6];
        shifterReg_6_0_bits_decodeResult_adder = _RANDOM[9'h2D][7];
        shifterReg_6_0_bits_decodeResult_logic = _RANDOM[9'h2D][8];
        shifterReg_6_0_bits_loadStore = _RANDOM[9'h2D][9];
        shifterReg_6_0_bits_issueInst = _RANDOM[9'h2D][10];
        shifterReg_6_0_bits_store = _RANDOM[9'h2D][11];
        shifterReg_6_0_bits_special = _RANDOM[9'h2D][12];
        shifterReg_6_0_bits_lsWholeReg = _RANDOM[9'h2D][13];
        shifterReg_6_0_bits_vs1 = _RANDOM[9'h2D][18:14];
        shifterReg_6_0_bits_vs2 = _RANDOM[9'h2D][23:19];
        shifterReg_6_0_bits_vd = _RANDOM[9'h2D][28:24];
        shifterReg_6_0_bits_loadStoreEEW = _RANDOM[9'h2D][30:29];
        shifterReg_6_0_bits_mask = _RANDOM[9'h2D][31];
        shifterReg_6_0_bits_segment = _RANDOM[9'h2E][2:0];
        shifterReg_6_0_bits_readFromScalar = {_RANDOM[9'h2E][31:3], _RANDOM[9'h2F][2:0]};
        shifterReg_6_0_bits_csrInterface_vl = _RANDOM[9'h2F][14:3];
        shifterReg_6_0_bits_csrInterface_vStart = _RANDOM[9'h2F][26:15];
        shifterReg_6_0_bits_csrInterface_vlmul = _RANDOM[9'h2F][29:27];
        shifterReg_6_0_bits_csrInterface_vSew = _RANDOM[9'h2F][31:30];
        shifterReg_6_0_bits_csrInterface_vxrm = _RANDOM[9'h30][1:0];
        shifterReg_6_0_bits_csrInterface_vta = _RANDOM[9'h30][2];
        shifterReg_6_0_bits_csrInterface_vma = _RANDOM[9'h30][3];
        releasePipe_pipe_v_7 = _RANDOM[9'h30][4];
        tokenCheck_counter_7 = _RANDOM[9'h30][7:5];
        shifterReg_7_0_valid = _RANDOM[9'h30][8];
        shifterReg_7_0_bits_instructionIndex = _RANDOM[9'h30][11:9];
        shifterReg_7_0_bits_decodeResult_orderReduce = _RANDOM[9'h30][12];
        shifterReg_7_0_bits_decodeResult_floatMul = _RANDOM[9'h30][13];
        shifterReg_7_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h30][15:14];
        shifterReg_7_0_bits_decodeResult_float = _RANDOM[9'h30][16];
        shifterReg_7_0_bits_decodeResult_specialSlot = _RANDOM[9'h30][17];
        shifterReg_7_0_bits_decodeResult_topUop = _RANDOM[9'h30][22:18];
        shifterReg_7_0_bits_decodeResult_popCount = _RANDOM[9'h30][23];
        shifterReg_7_0_bits_decodeResult_ffo = _RANDOM[9'h30][24];
        shifterReg_7_0_bits_decodeResult_average = _RANDOM[9'h30][25];
        shifterReg_7_0_bits_decodeResult_reverse = _RANDOM[9'h30][26];
        shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h30][27];
        shifterReg_7_0_bits_decodeResult_scheduler = _RANDOM[9'h30][28];
        shifterReg_7_0_bits_decodeResult_sReadVD = _RANDOM[9'h30][29];
        shifterReg_7_0_bits_decodeResult_vtype = _RANDOM[9'h30][30];
        shifterReg_7_0_bits_decodeResult_sWrite = _RANDOM[9'h30][31];
        shifterReg_7_0_bits_decodeResult_crossRead = _RANDOM[9'h31][0];
        shifterReg_7_0_bits_decodeResult_crossWrite = _RANDOM[9'h31][1];
        shifterReg_7_0_bits_decodeResult_maskUnit = _RANDOM[9'h31][2];
        shifterReg_7_0_bits_decodeResult_special = _RANDOM[9'h31][3];
        shifterReg_7_0_bits_decodeResult_saturate = _RANDOM[9'h31][4];
        shifterReg_7_0_bits_decodeResult_vwmacc = _RANDOM[9'h31][5];
        shifterReg_7_0_bits_decodeResult_readOnly = _RANDOM[9'h31][6];
        shifterReg_7_0_bits_decodeResult_maskSource = _RANDOM[9'h31][7];
        shifterReg_7_0_bits_decodeResult_maskDestination = _RANDOM[9'h31][8];
        shifterReg_7_0_bits_decodeResult_maskLogic = _RANDOM[9'h31][9];
        shifterReg_7_0_bits_decodeResult_uop = _RANDOM[9'h31][13:10];
        shifterReg_7_0_bits_decodeResult_iota = _RANDOM[9'h31][14];
        shifterReg_7_0_bits_decodeResult_mv = _RANDOM[9'h31][15];
        shifterReg_7_0_bits_decodeResult_extend = _RANDOM[9'h31][16];
        shifterReg_7_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h31][17];
        shifterReg_7_0_bits_decodeResult_compress = _RANDOM[9'h31][18];
        shifterReg_7_0_bits_decodeResult_gather16 = _RANDOM[9'h31][19];
        shifterReg_7_0_bits_decodeResult_gather = _RANDOM[9'h31][20];
        shifterReg_7_0_bits_decodeResult_slid = _RANDOM[9'h31][21];
        shifterReg_7_0_bits_decodeResult_targetRd = _RANDOM[9'h31][22];
        shifterReg_7_0_bits_decodeResult_widenReduce = _RANDOM[9'h31][23];
        shifterReg_7_0_bits_decodeResult_red = _RANDOM[9'h31][24];
        shifterReg_7_0_bits_decodeResult_nr = _RANDOM[9'h31][25];
        shifterReg_7_0_bits_decodeResult_itype = _RANDOM[9'h31][26];
        shifterReg_7_0_bits_decodeResult_unsigned1 = _RANDOM[9'h31][27];
        shifterReg_7_0_bits_decodeResult_unsigned0 = _RANDOM[9'h31][28];
        shifterReg_7_0_bits_decodeResult_other = _RANDOM[9'h31][29];
        shifterReg_7_0_bits_decodeResult_multiCycle = _RANDOM[9'h31][30];
        shifterReg_7_0_bits_decodeResult_divider = _RANDOM[9'h31][31];
        shifterReg_7_0_bits_decodeResult_multiplier = _RANDOM[9'h32][0];
        shifterReg_7_0_bits_decodeResult_shift = _RANDOM[9'h32][1];
        shifterReg_7_0_bits_decodeResult_adder = _RANDOM[9'h32][2];
        shifterReg_7_0_bits_decodeResult_logic = _RANDOM[9'h32][3];
        shifterReg_7_0_bits_loadStore = _RANDOM[9'h32][4];
        shifterReg_7_0_bits_issueInst = _RANDOM[9'h32][5];
        shifterReg_7_0_bits_store = _RANDOM[9'h32][6];
        shifterReg_7_0_bits_special = _RANDOM[9'h32][7];
        shifterReg_7_0_bits_lsWholeReg = _RANDOM[9'h32][8];
        shifterReg_7_0_bits_vs1 = _RANDOM[9'h32][13:9];
        shifterReg_7_0_bits_vs2 = _RANDOM[9'h32][18:14];
        shifterReg_7_0_bits_vd = _RANDOM[9'h32][23:19];
        shifterReg_7_0_bits_loadStoreEEW = _RANDOM[9'h32][25:24];
        shifterReg_7_0_bits_mask = _RANDOM[9'h32][26];
        shifterReg_7_0_bits_segment = _RANDOM[9'h32][29:27];
        shifterReg_7_0_bits_readFromScalar = {_RANDOM[9'h32][31:30], _RANDOM[9'h33][29:0]};
        shifterReg_7_0_bits_csrInterface_vl = {_RANDOM[9'h33][31:30], _RANDOM[9'h34][9:0]};
        shifterReg_7_0_bits_csrInterface_vStart = _RANDOM[9'h34][21:10];
        shifterReg_7_0_bits_csrInterface_vlmul = _RANDOM[9'h34][24:22];
        shifterReg_7_0_bits_csrInterface_vSew = _RANDOM[9'h34][26:25];
        shifterReg_7_0_bits_csrInterface_vxrm = _RANDOM[9'h34][28:27];
        shifterReg_7_0_bits_csrInterface_vta = _RANDOM[9'h34][29];
        shifterReg_7_0_bits_csrInterface_vma = _RANDOM[9'h34][30];
        releasePipe_pipe_v_8 = _RANDOM[9'h34][31];
        tokenCheck_counter_8 = _RANDOM[9'h35][2:0];
        shifterReg_8_0_valid = _RANDOM[9'h35][3];
        shifterReg_8_0_bits_instructionIndex = _RANDOM[9'h35][6:4];
        shifterReg_8_0_bits_decodeResult_orderReduce = _RANDOM[9'h35][7];
        shifterReg_8_0_bits_decodeResult_floatMul = _RANDOM[9'h35][8];
        shifterReg_8_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h35][10:9];
        shifterReg_8_0_bits_decodeResult_float = _RANDOM[9'h35][11];
        shifterReg_8_0_bits_decodeResult_specialSlot = _RANDOM[9'h35][12];
        shifterReg_8_0_bits_decodeResult_topUop = _RANDOM[9'h35][17:13];
        shifterReg_8_0_bits_decodeResult_popCount = _RANDOM[9'h35][18];
        shifterReg_8_0_bits_decodeResult_ffo = _RANDOM[9'h35][19];
        shifterReg_8_0_bits_decodeResult_average = _RANDOM[9'h35][20];
        shifterReg_8_0_bits_decodeResult_reverse = _RANDOM[9'h35][21];
        shifterReg_8_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h35][22];
        shifterReg_8_0_bits_decodeResult_scheduler = _RANDOM[9'h35][23];
        shifterReg_8_0_bits_decodeResult_sReadVD = _RANDOM[9'h35][24];
        shifterReg_8_0_bits_decodeResult_vtype = _RANDOM[9'h35][25];
        shifterReg_8_0_bits_decodeResult_sWrite = _RANDOM[9'h35][26];
        shifterReg_8_0_bits_decodeResult_crossRead = _RANDOM[9'h35][27];
        shifterReg_8_0_bits_decodeResult_crossWrite = _RANDOM[9'h35][28];
        shifterReg_8_0_bits_decodeResult_maskUnit = _RANDOM[9'h35][29];
        shifterReg_8_0_bits_decodeResult_special = _RANDOM[9'h35][30];
        shifterReg_8_0_bits_decodeResult_saturate = _RANDOM[9'h35][31];
        shifterReg_8_0_bits_decodeResult_vwmacc = _RANDOM[9'h36][0];
        shifterReg_8_0_bits_decodeResult_readOnly = _RANDOM[9'h36][1];
        shifterReg_8_0_bits_decodeResult_maskSource = _RANDOM[9'h36][2];
        shifterReg_8_0_bits_decodeResult_maskDestination = _RANDOM[9'h36][3];
        shifterReg_8_0_bits_decodeResult_maskLogic = _RANDOM[9'h36][4];
        shifterReg_8_0_bits_decodeResult_uop = _RANDOM[9'h36][8:5];
        shifterReg_8_0_bits_decodeResult_iota = _RANDOM[9'h36][9];
        shifterReg_8_0_bits_decodeResult_mv = _RANDOM[9'h36][10];
        shifterReg_8_0_bits_decodeResult_extend = _RANDOM[9'h36][11];
        shifterReg_8_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h36][12];
        shifterReg_8_0_bits_decodeResult_compress = _RANDOM[9'h36][13];
        shifterReg_8_0_bits_decodeResult_gather16 = _RANDOM[9'h36][14];
        shifterReg_8_0_bits_decodeResult_gather = _RANDOM[9'h36][15];
        shifterReg_8_0_bits_decodeResult_slid = _RANDOM[9'h36][16];
        shifterReg_8_0_bits_decodeResult_targetRd = _RANDOM[9'h36][17];
        shifterReg_8_0_bits_decodeResult_widenReduce = _RANDOM[9'h36][18];
        shifterReg_8_0_bits_decodeResult_red = _RANDOM[9'h36][19];
        shifterReg_8_0_bits_decodeResult_nr = _RANDOM[9'h36][20];
        shifterReg_8_0_bits_decodeResult_itype = _RANDOM[9'h36][21];
        shifterReg_8_0_bits_decodeResult_unsigned1 = _RANDOM[9'h36][22];
        shifterReg_8_0_bits_decodeResult_unsigned0 = _RANDOM[9'h36][23];
        shifterReg_8_0_bits_decodeResult_other = _RANDOM[9'h36][24];
        shifterReg_8_0_bits_decodeResult_multiCycle = _RANDOM[9'h36][25];
        shifterReg_8_0_bits_decodeResult_divider = _RANDOM[9'h36][26];
        shifterReg_8_0_bits_decodeResult_multiplier = _RANDOM[9'h36][27];
        shifterReg_8_0_bits_decodeResult_shift = _RANDOM[9'h36][28];
        shifterReg_8_0_bits_decodeResult_adder = _RANDOM[9'h36][29];
        shifterReg_8_0_bits_decodeResult_logic = _RANDOM[9'h36][30];
        shifterReg_8_0_bits_loadStore = _RANDOM[9'h36][31];
        shifterReg_8_0_bits_issueInst = _RANDOM[9'h37][0];
        shifterReg_8_0_bits_store = _RANDOM[9'h37][1];
        shifterReg_8_0_bits_special = _RANDOM[9'h37][2];
        shifterReg_8_0_bits_lsWholeReg = _RANDOM[9'h37][3];
        shifterReg_8_0_bits_vs1 = _RANDOM[9'h37][8:4];
        shifterReg_8_0_bits_vs2 = _RANDOM[9'h37][13:9];
        shifterReg_8_0_bits_vd = _RANDOM[9'h37][18:14];
        shifterReg_8_0_bits_loadStoreEEW = _RANDOM[9'h37][20:19];
        shifterReg_8_0_bits_mask = _RANDOM[9'h37][21];
        shifterReg_8_0_bits_segment = _RANDOM[9'h37][24:22];
        shifterReg_8_0_bits_readFromScalar = {_RANDOM[9'h37][31:25], _RANDOM[9'h38][24:0]};
        shifterReg_8_0_bits_csrInterface_vl = {_RANDOM[9'h38][31:25], _RANDOM[9'h39][4:0]};
        shifterReg_8_0_bits_csrInterface_vStart = _RANDOM[9'h39][16:5];
        shifterReg_8_0_bits_csrInterface_vlmul = _RANDOM[9'h39][19:17];
        shifterReg_8_0_bits_csrInterface_vSew = _RANDOM[9'h39][21:20];
        shifterReg_8_0_bits_csrInterface_vxrm = _RANDOM[9'h39][23:22];
        shifterReg_8_0_bits_csrInterface_vta = _RANDOM[9'h39][24];
        shifterReg_8_0_bits_csrInterface_vma = _RANDOM[9'h39][25];
        releasePipe_pipe_v_9 = _RANDOM[9'h39][26];
        tokenCheck_counter_9 = _RANDOM[9'h39][29:27];
        shifterReg_9_0_valid = _RANDOM[9'h39][30];
        shifterReg_9_0_bits_instructionIndex = {_RANDOM[9'h39][31], _RANDOM[9'h3A][1:0]};
        shifterReg_9_0_bits_decodeResult_orderReduce = _RANDOM[9'h3A][2];
        shifterReg_9_0_bits_decodeResult_floatMul = _RANDOM[9'h3A][3];
        shifterReg_9_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h3A][5:4];
        shifterReg_9_0_bits_decodeResult_float = _RANDOM[9'h3A][6];
        shifterReg_9_0_bits_decodeResult_specialSlot = _RANDOM[9'h3A][7];
        shifterReg_9_0_bits_decodeResult_topUop = _RANDOM[9'h3A][12:8];
        shifterReg_9_0_bits_decodeResult_popCount = _RANDOM[9'h3A][13];
        shifterReg_9_0_bits_decodeResult_ffo = _RANDOM[9'h3A][14];
        shifterReg_9_0_bits_decodeResult_average = _RANDOM[9'h3A][15];
        shifterReg_9_0_bits_decodeResult_reverse = _RANDOM[9'h3A][16];
        shifterReg_9_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h3A][17];
        shifterReg_9_0_bits_decodeResult_scheduler = _RANDOM[9'h3A][18];
        shifterReg_9_0_bits_decodeResult_sReadVD = _RANDOM[9'h3A][19];
        shifterReg_9_0_bits_decodeResult_vtype = _RANDOM[9'h3A][20];
        shifterReg_9_0_bits_decodeResult_sWrite = _RANDOM[9'h3A][21];
        shifterReg_9_0_bits_decodeResult_crossRead = _RANDOM[9'h3A][22];
        shifterReg_9_0_bits_decodeResult_crossWrite = _RANDOM[9'h3A][23];
        shifterReg_9_0_bits_decodeResult_maskUnit = _RANDOM[9'h3A][24];
        shifterReg_9_0_bits_decodeResult_special = _RANDOM[9'h3A][25];
        shifterReg_9_0_bits_decodeResult_saturate = _RANDOM[9'h3A][26];
        shifterReg_9_0_bits_decodeResult_vwmacc = _RANDOM[9'h3A][27];
        shifterReg_9_0_bits_decodeResult_readOnly = _RANDOM[9'h3A][28];
        shifterReg_9_0_bits_decodeResult_maskSource = _RANDOM[9'h3A][29];
        shifterReg_9_0_bits_decodeResult_maskDestination = _RANDOM[9'h3A][30];
        shifterReg_9_0_bits_decodeResult_maskLogic = _RANDOM[9'h3A][31];
        shifterReg_9_0_bits_decodeResult_uop = _RANDOM[9'h3B][3:0];
        shifterReg_9_0_bits_decodeResult_iota = _RANDOM[9'h3B][4];
        shifterReg_9_0_bits_decodeResult_mv = _RANDOM[9'h3B][5];
        shifterReg_9_0_bits_decodeResult_extend = _RANDOM[9'h3B][6];
        shifterReg_9_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h3B][7];
        shifterReg_9_0_bits_decodeResult_compress = _RANDOM[9'h3B][8];
        shifterReg_9_0_bits_decodeResult_gather16 = _RANDOM[9'h3B][9];
        shifterReg_9_0_bits_decodeResult_gather = _RANDOM[9'h3B][10];
        shifterReg_9_0_bits_decodeResult_slid = _RANDOM[9'h3B][11];
        shifterReg_9_0_bits_decodeResult_targetRd = _RANDOM[9'h3B][12];
        shifterReg_9_0_bits_decodeResult_widenReduce = _RANDOM[9'h3B][13];
        shifterReg_9_0_bits_decodeResult_red = _RANDOM[9'h3B][14];
        shifterReg_9_0_bits_decodeResult_nr = _RANDOM[9'h3B][15];
        shifterReg_9_0_bits_decodeResult_itype = _RANDOM[9'h3B][16];
        shifterReg_9_0_bits_decodeResult_unsigned1 = _RANDOM[9'h3B][17];
        shifterReg_9_0_bits_decodeResult_unsigned0 = _RANDOM[9'h3B][18];
        shifterReg_9_0_bits_decodeResult_other = _RANDOM[9'h3B][19];
        shifterReg_9_0_bits_decodeResult_multiCycle = _RANDOM[9'h3B][20];
        shifterReg_9_0_bits_decodeResult_divider = _RANDOM[9'h3B][21];
        shifterReg_9_0_bits_decodeResult_multiplier = _RANDOM[9'h3B][22];
        shifterReg_9_0_bits_decodeResult_shift = _RANDOM[9'h3B][23];
        shifterReg_9_0_bits_decodeResult_adder = _RANDOM[9'h3B][24];
        shifterReg_9_0_bits_decodeResult_logic = _RANDOM[9'h3B][25];
        shifterReg_9_0_bits_loadStore = _RANDOM[9'h3B][26];
        shifterReg_9_0_bits_issueInst = _RANDOM[9'h3B][27];
        shifterReg_9_0_bits_store = _RANDOM[9'h3B][28];
        shifterReg_9_0_bits_special = _RANDOM[9'h3B][29];
        shifterReg_9_0_bits_lsWholeReg = _RANDOM[9'h3B][30];
        shifterReg_9_0_bits_vs1 = {_RANDOM[9'h3B][31], _RANDOM[9'h3C][3:0]};
        shifterReg_9_0_bits_vs2 = _RANDOM[9'h3C][8:4];
        shifterReg_9_0_bits_vd = _RANDOM[9'h3C][13:9];
        shifterReg_9_0_bits_loadStoreEEW = _RANDOM[9'h3C][15:14];
        shifterReg_9_0_bits_mask = _RANDOM[9'h3C][16];
        shifterReg_9_0_bits_segment = _RANDOM[9'h3C][19:17];
        shifterReg_9_0_bits_readFromScalar = {_RANDOM[9'h3C][31:20], _RANDOM[9'h3D][19:0]};
        shifterReg_9_0_bits_csrInterface_vl = _RANDOM[9'h3D][31:20];
        shifterReg_9_0_bits_csrInterface_vStart = _RANDOM[9'h3E][11:0];
        shifterReg_9_0_bits_csrInterface_vlmul = _RANDOM[9'h3E][14:12];
        shifterReg_9_0_bits_csrInterface_vSew = _RANDOM[9'h3E][16:15];
        shifterReg_9_0_bits_csrInterface_vxrm = _RANDOM[9'h3E][18:17];
        shifterReg_9_0_bits_csrInterface_vta = _RANDOM[9'h3E][19];
        shifterReg_9_0_bits_csrInterface_vma = _RANDOM[9'h3E][20];
        releasePipe_pipe_v_10 = _RANDOM[9'h3E][21];
        tokenCheck_counter_10 = _RANDOM[9'h3E][24:22];
        shifterReg_10_0_valid = _RANDOM[9'h3E][25];
        shifterReg_10_0_bits_instructionIndex = _RANDOM[9'h3E][28:26];
        shifterReg_10_0_bits_decodeResult_orderReduce = _RANDOM[9'h3E][29];
        shifterReg_10_0_bits_decodeResult_floatMul = _RANDOM[9'h3E][30];
        shifterReg_10_0_bits_decodeResult_fpExecutionType = {_RANDOM[9'h3E][31], _RANDOM[9'h3F][0]};
        shifterReg_10_0_bits_decodeResult_float = _RANDOM[9'h3F][1];
        shifterReg_10_0_bits_decodeResult_specialSlot = _RANDOM[9'h3F][2];
        shifterReg_10_0_bits_decodeResult_topUop = _RANDOM[9'h3F][7:3];
        shifterReg_10_0_bits_decodeResult_popCount = _RANDOM[9'h3F][8];
        shifterReg_10_0_bits_decodeResult_ffo = _RANDOM[9'h3F][9];
        shifterReg_10_0_bits_decodeResult_average = _RANDOM[9'h3F][10];
        shifterReg_10_0_bits_decodeResult_reverse = _RANDOM[9'h3F][11];
        shifterReg_10_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h3F][12];
        shifterReg_10_0_bits_decodeResult_scheduler = _RANDOM[9'h3F][13];
        shifterReg_10_0_bits_decodeResult_sReadVD = _RANDOM[9'h3F][14];
        shifterReg_10_0_bits_decodeResult_vtype = _RANDOM[9'h3F][15];
        shifterReg_10_0_bits_decodeResult_sWrite = _RANDOM[9'h3F][16];
        shifterReg_10_0_bits_decodeResult_crossRead = _RANDOM[9'h3F][17];
        shifterReg_10_0_bits_decodeResult_crossWrite = _RANDOM[9'h3F][18];
        shifterReg_10_0_bits_decodeResult_maskUnit = _RANDOM[9'h3F][19];
        shifterReg_10_0_bits_decodeResult_special = _RANDOM[9'h3F][20];
        shifterReg_10_0_bits_decodeResult_saturate = _RANDOM[9'h3F][21];
        shifterReg_10_0_bits_decodeResult_vwmacc = _RANDOM[9'h3F][22];
        shifterReg_10_0_bits_decodeResult_readOnly = _RANDOM[9'h3F][23];
        shifterReg_10_0_bits_decodeResult_maskSource = _RANDOM[9'h3F][24];
        shifterReg_10_0_bits_decodeResult_maskDestination = _RANDOM[9'h3F][25];
        shifterReg_10_0_bits_decodeResult_maskLogic = _RANDOM[9'h3F][26];
        shifterReg_10_0_bits_decodeResult_uop = _RANDOM[9'h3F][30:27];
        shifterReg_10_0_bits_decodeResult_iota = _RANDOM[9'h3F][31];
        shifterReg_10_0_bits_decodeResult_mv = _RANDOM[9'h40][0];
        shifterReg_10_0_bits_decodeResult_extend = _RANDOM[9'h40][1];
        shifterReg_10_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h40][2];
        shifterReg_10_0_bits_decodeResult_compress = _RANDOM[9'h40][3];
        shifterReg_10_0_bits_decodeResult_gather16 = _RANDOM[9'h40][4];
        shifterReg_10_0_bits_decodeResult_gather = _RANDOM[9'h40][5];
        shifterReg_10_0_bits_decodeResult_slid = _RANDOM[9'h40][6];
        shifterReg_10_0_bits_decodeResult_targetRd = _RANDOM[9'h40][7];
        shifterReg_10_0_bits_decodeResult_widenReduce = _RANDOM[9'h40][8];
        shifterReg_10_0_bits_decodeResult_red = _RANDOM[9'h40][9];
        shifterReg_10_0_bits_decodeResult_nr = _RANDOM[9'h40][10];
        shifterReg_10_0_bits_decodeResult_itype = _RANDOM[9'h40][11];
        shifterReg_10_0_bits_decodeResult_unsigned1 = _RANDOM[9'h40][12];
        shifterReg_10_0_bits_decodeResult_unsigned0 = _RANDOM[9'h40][13];
        shifterReg_10_0_bits_decodeResult_other = _RANDOM[9'h40][14];
        shifterReg_10_0_bits_decodeResult_multiCycle = _RANDOM[9'h40][15];
        shifterReg_10_0_bits_decodeResult_divider = _RANDOM[9'h40][16];
        shifterReg_10_0_bits_decodeResult_multiplier = _RANDOM[9'h40][17];
        shifterReg_10_0_bits_decodeResult_shift = _RANDOM[9'h40][18];
        shifterReg_10_0_bits_decodeResult_adder = _RANDOM[9'h40][19];
        shifterReg_10_0_bits_decodeResult_logic = _RANDOM[9'h40][20];
        shifterReg_10_0_bits_loadStore = _RANDOM[9'h40][21];
        shifterReg_10_0_bits_issueInst = _RANDOM[9'h40][22];
        shifterReg_10_0_bits_store = _RANDOM[9'h40][23];
        shifterReg_10_0_bits_special = _RANDOM[9'h40][24];
        shifterReg_10_0_bits_lsWholeReg = _RANDOM[9'h40][25];
        shifterReg_10_0_bits_vs1 = _RANDOM[9'h40][30:26];
        shifterReg_10_0_bits_vs2 = {_RANDOM[9'h40][31], _RANDOM[9'h41][3:0]};
        shifterReg_10_0_bits_vd = _RANDOM[9'h41][8:4];
        shifterReg_10_0_bits_loadStoreEEW = _RANDOM[9'h41][10:9];
        shifterReg_10_0_bits_mask = _RANDOM[9'h41][11];
        shifterReg_10_0_bits_segment = _RANDOM[9'h41][14:12];
        shifterReg_10_0_bits_readFromScalar = {_RANDOM[9'h41][31:15], _RANDOM[9'h42][14:0]};
        shifterReg_10_0_bits_csrInterface_vl = _RANDOM[9'h42][26:15];
        shifterReg_10_0_bits_csrInterface_vStart = {_RANDOM[9'h42][31:27], _RANDOM[9'h43][6:0]};
        shifterReg_10_0_bits_csrInterface_vlmul = _RANDOM[9'h43][9:7];
        shifterReg_10_0_bits_csrInterface_vSew = _RANDOM[9'h43][11:10];
        shifterReg_10_0_bits_csrInterface_vxrm = _RANDOM[9'h43][13:12];
        shifterReg_10_0_bits_csrInterface_vta = _RANDOM[9'h43][14];
        shifterReg_10_0_bits_csrInterface_vma = _RANDOM[9'h43][15];
        releasePipe_pipe_v_11 = _RANDOM[9'h43][16];
        tokenCheck_counter_11 = _RANDOM[9'h43][19:17];
        shifterReg_11_0_valid = _RANDOM[9'h43][20];
        shifterReg_11_0_bits_instructionIndex = _RANDOM[9'h43][23:21];
        shifterReg_11_0_bits_decodeResult_orderReduce = _RANDOM[9'h43][24];
        shifterReg_11_0_bits_decodeResult_floatMul = _RANDOM[9'h43][25];
        shifterReg_11_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h43][27:26];
        shifterReg_11_0_bits_decodeResult_float = _RANDOM[9'h43][28];
        shifterReg_11_0_bits_decodeResult_specialSlot = _RANDOM[9'h43][29];
        shifterReg_11_0_bits_decodeResult_topUop = {_RANDOM[9'h43][31:30], _RANDOM[9'h44][2:0]};
        shifterReg_11_0_bits_decodeResult_popCount = _RANDOM[9'h44][3];
        shifterReg_11_0_bits_decodeResult_ffo = _RANDOM[9'h44][4];
        shifterReg_11_0_bits_decodeResult_average = _RANDOM[9'h44][5];
        shifterReg_11_0_bits_decodeResult_reverse = _RANDOM[9'h44][6];
        shifterReg_11_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h44][7];
        shifterReg_11_0_bits_decodeResult_scheduler = _RANDOM[9'h44][8];
        shifterReg_11_0_bits_decodeResult_sReadVD = _RANDOM[9'h44][9];
        shifterReg_11_0_bits_decodeResult_vtype = _RANDOM[9'h44][10];
        shifterReg_11_0_bits_decodeResult_sWrite = _RANDOM[9'h44][11];
        shifterReg_11_0_bits_decodeResult_crossRead = _RANDOM[9'h44][12];
        shifterReg_11_0_bits_decodeResult_crossWrite = _RANDOM[9'h44][13];
        shifterReg_11_0_bits_decodeResult_maskUnit = _RANDOM[9'h44][14];
        shifterReg_11_0_bits_decodeResult_special = _RANDOM[9'h44][15];
        shifterReg_11_0_bits_decodeResult_saturate = _RANDOM[9'h44][16];
        shifterReg_11_0_bits_decodeResult_vwmacc = _RANDOM[9'h44][17];
        shifterReg_11_0_bits_decodeResult_readOnly = _RANDOM[9'h44][18];
        shifterReg_11_0_bits_decodeResult_maskSource = _RANDOM[9'h44][19];
        shifterReg_11_0_bits_decodeResult_maskDestination = _RANDOM[9'h44][20];
        shifterReg_11_0_bits_decodeResult_maskLogic = _RANDOM[9'h44][21];
        shifterReg_11_0_bits_decodeResult_uop = _RANDOM[9'h44][25:22];
        shifterReg_11_0_bits_decodeResult_iota = _RANDOM[9'h44][26];
        shifterReg_11_0_bits_decodeResult_mv = _RANDOM[9'h44][27];
        shifterReg_11_0_bits_decodeResult_extend = _RANDOM[9'h44][28];
        shifterReg_11_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h44][29];
        shifterReg_11_0_bits_decodeResult_compress = _RANDOM[9'h44][30];
        shifterReg_11_0_bits_decodeResult_gather16 = _RANDOM[9'h44][31];
        shifterReg_11_0_bits_decodeResult_gather = _RANDOM[9'h45][0];
        shifterReg_11_0_bits_decodeResult_slid = _RANDOM[9'h45][1];
        shifterReg_11_0_bits_decodeResult_targetRd = _RANDOM[9'h45][2];
        shifterReg_11_0_bits_decodeResult_widenReduce = _RANDOM[9'h45][3];
        shifterReg_11_0_bits_decodeResult_red = _RANDOM[9'h45][4];
        shifterReg_11_0_bits_decodeResult_nr = _RANDOM[9'h45][5];
        shifterReg_11_0_bits_decodeResult_itype = _RANDOM[9'h45][6];
        shifterReg_11_0_bits_decodeResult_unsigned1 = _RANDOM[9'h45][7];
        shifterReg_11_0_bits_decodeResult_unsigned0 = _RANDOM[9'h45][8];
        shifterReg_11_0_bits_decodeResult_other = _RANDOM[9'h45][9];
        shifterReg_11_0_bits_decodeResult_multiCycle = _RANDOM[9'h45][10];
        shifterReg_11_0_bits_decodeResult_divider = _RANDOM[9'h45][11];
        shifterReg_11_0_bits_decodeResult_multiplier = _RANDOM[9'h45][12];
        shifterReg_11_0_bits_decodeResult_shift = _RANDOM[9'h45][13];
        shifterReg_11_0_bits_decodeResult_adder = _RANDOM[9'h45][14];
        shifterReg_11_0_bits_decodeResult_logic = _RANDOM[9'h45][15];
        shifterReg_11_0_bits_loadStore = _RANDOM[9'h45][16];
        shifterReg_11_0_bits_issueInst = _RANDOM[9'h45][17];
        shifterReg_11_0_bits_store = _RANDOM[9'h45][18];
        shifterReg_11_0_bits_special = _RANDOM[9'h45][19];
        shifterReg_11_0_bits_lsWholeReg = _RANDOM[9'h45][20];
        shifterReg_11_0_bits_vs1 = _RANDOM[9'h45][25:21];
        shifterReg_11_0_bits_vs2 = _RANDOM[9'h45][30:26];
        shifterReg_11_0_bits_vd = {_RANDOM[9'h45][31], _RANDOM[9'h46][3:0]};
        shifterReg_11_0_bits_loadStoreEEW = _RANDOM[9'h46][5:4];
        shifterReg_11_0_bits_mask = _RANDOM[9'h46][6];
        shifterReg_11_0_bits_segment = _RANDOM[9'h46][9:7];
        shifterReg_11_0_bits_readFromScalar = {_RANDOM[9'h46][31:10], _RANDOM[9'h47][9:0]};
        shifterReg_11_0_bits_csrInterface_vl = _RANDOM[9'h47][21:10];
        shifterReg_11_0_bits_csrInterface_vStart = {_RANDOM[9'h47][31:22], _RANDOM[9'h48][1:0]};
        shifterReg_11_0_bits_csrInterface_vlmul = _RANDOM[9'h48][4:2];
        shifterReg_11_0_bits_csrInterface_vSew = _RANDOM[9'h48][6:5];
        shifterReg_11_0_bits_csrInterface_vxrm = _RANDOM[9'h48][8:7];
        shifterReg_11_0_bits_csrInterface_vta = _RANDOM[9'h48][9];
        shifterReg_11_0_bits_csrInterface_vma = _RANDOM[9'h48][10];
        releasePipe_pipe_v_12 = _RANDOM[9'h48][11];
        tokenCheck_counter_12 = _RANDOM[9'h48][14:12];
        shifterReg_12_0_valid = _RANDOM[9'h48][15];
        shifterReg_12_0_bits_instructionIndex = _RANDOM[9'h48][18:16];
        shifterReg_12_0_bits_decodeResult_orderReduce = _RANDOM[9'h48][19];
        shifterReg_12_0_bits_decodeResult_floatMul = _RANDOM[9'h48][20];
        shifterReg_12_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h48][22:21];
        shifterReg_12_0_bits_decodeResult_float = _RANDOM[9'h48][23];
        shifterReg_12_0_bits_decodeResult_specialSlot = _RANDOM[9'h48][24];
        shifterReg_12_0_bits_decodeResult_topUop = _RANDOM[9'h48][29:25];
        shifterReg_12_0_bits_decodeResult_popCount = _RANDOM[9'h48][30];
        shifterReg_12_0_bits_decodeResult_ffo = _RANDOM[9'h48][31];
        shifterReg_12_0_bits_decodeResult_average = _RANDOM[9'h49][0];
        shifterReg_12_0_bits_decodeResult_reverse = _RANDOM[9'h49][1];
        shifterReg_12_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h49][2];
        shifterReg_12_0_bits_decodeResult_scheduler = _RANDOM[9'h49][3];
        shifterReg_12_0_bits_decodeResult_sReadVD = _RANDOM[9'h49][4];
        shifterReg_12_0_bits_decodeResult_vtype = _RANDOM[9'h49][5];
        shifterReg_12_0_bits_decodeResult_sWrite = _RANDOM[9'h49][6];
        shifterReg_12_0_bits_decodeResult_crossRead = _RANDOM[9'h49][7];
        shifterReg_12_0_bits_decodeResult_crossWrite = _RANDOM[9'h49][8];
        shifterReg_12_0_bits_decodeResult_maskUnit = _RANDOM[9'h49][9];
        shifterReg_12_0_bits_decodeResult_special = _RANDOM[9'h49][10];
        shifterReg_12_0_bits_decodeResult_saturate = _RANDOM[9'h49][11];
        shifterReg_12_0_bits_decodeResult_vwmacc = _RANDOM[9'h49][12];
        shifterReg_12_0_bits_decodeResult_readOnly = _RANDOM[9'h49][13];
        shifterReg_12_0_bits_decodeResult_maskSource = _RANDOM[9'h49][14];
        shifterReg_12_0_bits_decodeResult_maskDestination = _RANDOM[9'h49][15];
        shifterReg_12_0_bits_decodeResult_maskLogic = _RANDOM[9'h49][16];
        shifterReg_12_0_bits_decodeResult_uop = _RANDOM[9'h49][20:17];
        shifterReg_12_0_bits_decodeResult_iota = _RANDOM[9'h49][21];
        shifterReg_12_0_bits_decodeResult_mv = _RANDOM[9'h49][22];
        shifterReg_12_0_bits_decodeResult_extend = _RANDOM[9'h49][23];
        shifterReg_12_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h49][24];
        shifterReg_12_0_bits_decodeResult_compress = _RANDOM[9'h49][25];
        shifterReg_12_0_bits_decodeResult_gather16 = _RANDOM[9'h49][26];
        shifterReg_12_0_bits_decodeResult_gather = _RANDOM[9'h49][27];
        shifterReg_12_0_bits_decodeResult_slid = _RANDOM[9'h49][28];
        shifterReg_12_0_bits_decodeResult_targetRd = _RANDOM[9'h49][29];
        shifterReg_12_0_bits_decodeResult_widenReduce = _RANDOM[9'h49][30];
        shifterReg_12_0_bits_decodeResult_red = _RANDOM[9'h49][31];
        shifterReg_12_0_bits_decodeResult_nr = _RANDOM[9'h4A][0];
        shifterReg_12_0_bits_decodeResult_itype = _RANDOM[9'h4A][1];
        shifterReg_12_0_bits_decodeResult_unsigned1 = _RANDOM[9'h4A][2];
        shifterReg_12_0_bits_decodeResult_unsigned0 = _RANDOM[9'h4A][3];
        shifterReg_12_0_bits_decodeResult_other = _RANDOM[9'h4A][4];
        shifterReg_12_0_bits_decodeResult_multiCycle = _RANDOM[9'h4A][5];
        shifterReg_12_0_bits_decodeResult_divider = _RANDOM[9'h4A][6];
        shifterReg_12_0_bits_decodeResult_multiplier = _RANDOM[9'h4A][7];
        shifterReg_12_0_bits_decodeResult_shift = _RANDOM[9'h4A][8];
        shifterReg_12_0_bits_decodeResult_adder = _RANDOM[9'h4A][9];
        shifterReg_12_0_bits_decodeResult_logic = _RANDOM[9'h4A][10];
        shifterReg_12_0_bits_loadStore = _RANDOM[9'h4A][11];
        shifterReg_12_0_bits_issueInst = _RANDOM[9'h4A][12];
        shifterReg_12_0_bits_store = _RANDOM[9'h4A][13];
        shifterReg_12_0_bits_special = _RANDOM[9'h4A][14];
        shifterReg_12_0_bits_lsWholeReg = _RANDOM[9'h4A][15];
        shifterReg_12_0_bits_vs1 = _RANDOM[9'h4A][20:16];
        shifterReg_12_0_bits_vs2 = _RANDOM[9'h4A][25:21];
        shifterReg_12_0_bits_vd = _RANDOM[9'h4A][30:26];
        shifterReg_12_0_bits_loadStoreEEW = {_RANDOM[9'h4A][31], _RANDOM[9'h4B][0]};
        shifterReg_12_0_bits_mask = _RANDOM[9'h4B][1];
        shifterReg_12_0_bits_segment = _RANDOM[9'h4B][4:2];
        shifterReg_12_0_bits_readFromScalar = {_RANDOM[9'h4B][31:5], _RANDOM[9'h4C][4:0]};
        shifterReg_12_0_bits_csrInterface_vl = _RANDOM[9'h4C][16:5];
        shifterReg_12_0_bits_csrInterface_vStart = _RANDOM[9'h4C][28:17];
        shifterReg_12_0_bits_csrInterface_vlmul = _RANDOM[9'h4C][31:29];
        shifterReg_12_0_bits_csrInterface_vSew = _RANDOM[9'h4D][1:0];
        shifterReg_12_0_bits_csrInterface_vxrm = _RANDOM[9'h4D][3:2];
        shifterReg_12_0_bits_csrInterface_vta = _RANDOM[9'h4D][4];
        shifterReg_12_0_bits_csrInterface_vma = _RANDOM[9'h4D][5];
        releasePipe_pipe_v_13 = _RANDOM[9'h4D][6];
        tokenCheck_counter_13 = _RANDOM[9'h4D][9:7];
        shifterReg_13_0_valid = _RANDOM[9'h4D][10];
        shifterReg_13_0_bits_instructionIndex = _RANDOM[9'h4D][13:11];
        shifterReg_13_0_bits_decodeResult_orderReduce = _RANDOM[9'h4D][14];
        shifterReg_13_0_bits_decodeResult_floatMul = _RANDOM[9'h4D][15];
        shifterReg_13_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h4D][17:16];
        shifterReg_13_0_bits_decodeResult_float = _RANDOM[9'h4D][18];
        shifterReg_13_0_bits_decodeResult_specialSlot = _RANDOM[9'h4D][19];
        shifterReg_13_0_bits_decodeResult_topUop = _RANDOM[9'h4D][24:20];
        shifterReg_13_0_bits_decodeResult_popCount = _RANDOM[9'h4D][25];
        shifterReg_13_0_bits_decodeResult_ffo = _RANDOM[9'h4D][26];
        shifterReg_13_0_bits_decodeResult_average = _RANDOM[9'h4D][27];
        shifterReg_13_0_bits_decodeResult_reverse = _RANDOM[9'h4D][28];
        shifterReg_13_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h4D][29];
        shifterReg_13_0_bits_decodeResult_scheduler = _RANDOM[9'h4D][30];
        shifterReg_13_0_bits_decodeResult_sReadVD = _RANDOM[9'h4D][31];
        shifterReg_13_0_bits_decodeResult_vtype = _RANDOM[9'h4E][0];
        shifterReg_13_0_bits_decodeResult_sWrite = _RANDOM[9'h4E][1];
        shifterReg_13_0_bits_decodeResult_crossRead = _RANDOM[9'h4E][2];
        shifterReg_13_0_bits_decodeResult_crossWrite = _RANDOM[9'h4E][3];
        shifterReg_13_0_bits_decodeResult_maskUnit = _RANDOM[9'h4E][4];
        shifterReg_13_0_bits_decodeResult_special = _RANDOM[9'h4E][5];
        shifterReg_13_0_bits_decodeResult_saturate = _RANDOM[9'h4E][6];
        shifterReg_13_0_bits_decodeResult_vwmacc = _RANDOM[9'h4E][7];
        shifterReg_13_0_bits_decodeResult_readOnly = _RANDOM[9'h4E][8];
        shifterReg_13_0_bits_decodeResult_maskSource = _RANDOM[9'h4E][9];
        shifterReg_13_0_bits_decodeResult_maskDestination = _RANDOM[9'h4E][10];
        shifterReg_13_0_bits_decodeResult_maskLogic = _RANDOM[9'h4E][11];
        shifterReg_13_0_bits_decodeResult_uop = _RANDOM[9'h4E][15:12];
        shifterReg_13_0_bits_decodeResult_iota = _RANDOM[9'h4E][16];
        shifterReg_13_0_bits_decodeResult_mv = _RANDOM[9'h4E][17];
        shifterReg_13_0_bits_decodeResult_extend = _RANDOM[9'h4E][18];
        shifterReg_13_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h4E][19];
        shifterReg_13_0_bits_decodeResult_compress = _RANDOM[9'h4E][20];
        shifterReg_13_0_bits_decodeResult_gather16 = _RANDOM[9'h4E][21];
        shifterReg_13_0_bits_decodeResult_gather = _RANDOM[9'h4E][22];
        shifterReg_13_0_bits_decodeResult_slid = _RANDOM[9'h4E][23];
        shifterReg_13_0_bits_decodeResult_targetRd = _RANDOM[9'h4E][24];
        shifterReg_13_0_bits_decodeResult_widenReduce = _RANDOM[9'h4E][25];
        shifterReg_13_0_bits_decodeResult_red = _RANDOM[9'h4E][26];
        shifterReg_13_0_bits_decodeResult_nr = _RANDOM[9'h4E][27];
        shifterReg_13_0_bits_decodeResult_itype = _RANDOM[9'h4E][28];
        shifterReg_13_0_bits_decodeResult_unsigned1 = _RANDOM[9'h4E][29];
        shifterReg_13_0_bits_decodeResult_unsigned0 = _RANDOM[9'h4E][30];
        shifterReg_13_0_bits_decodeResult_other = _RANDOM[9'h4E][31];
        shifterReg_13_0_bits_decodeResult_multiCycle = _RANDOM[9'h4F][0];
        shifterReg_13_0_bits_decodeResult_divider = _RANDOM[9'h4F][1];
        shifterReg_13_0_bits_decodeResult_multiplier = _RANDOM[9'h4F][2];
        shifterReg_13_0_bits_decodeResult_shift = _RANDOM[9'h4F][3];
        shifterReg_13_0_bits_decodeResult_adder = _RANDOM[9'h4F][4];
        shifterReg_13_0_bits_decodeResult_logic = _RANDOM[9'h4F][5];
        shifterReg_13_0_bits_loadStore = _RANDOM[9'h4F][6];
        shifterReg_13_0_bits_issueInst = _RANDOM[9'h4F][7];
        shifterReg_13_0_bits_store = _RANDOM[9'h4F][8];
        shifterReg_13_0_bits_special = _RANDOM[9'h4F][9];
        shifterReg_13_0_bits_lsWholeReg = _RANDOM[9'h4F][10];
        shifterReg_13_0_bits_vs1 = _RANDOM[9'h4F][15:11];
        shifterReg_13_0_bits_vs2 = _RANDOM[9'h4F][20:16];
        shifterReg_13_0_bits_vd = _RANDOM[9'h4F][25:21];
        shifterReg_13_0_bits_loadStoreEEW = _RANDOM[9'h4F][27:26];
        shifterReg_13_0_bits_mask = _RANDOM[9'h4F][28];
        shifterReg_13_0_bits_segment = _RANDOM[9'h4F][31:29];
        shifterReg_13_0_bits_readFromScalar = _RANDOM[9'h50];
        shifterReg_13_0_bits_csrInterface_vl = _RANDOM[9'h51][11:0];
        shifterReg_13_0_bits_csrInterface_vStart = _RANDOM[9'h51][23:12];
        shifterReg_13_0_bits_csrInterface_vlmul = _RANDOM[9'h51][26:24];
        shifterReg_13_0_bits_csrInterface_vSew = _RANDOM[9'h51][28:27];
        shifterReg_13_0_bits_csrInterface_vxrm = _RANDOM[9'h51][30:29];
        shifterReg_13_0_bits_csrInterface_vta = _RANDOM[9'h51][31];
        shifterReg_13_0_bits_csrInterface_vma = _RANDOM[9'h52][0];
        releasePipe_pipe_v_14 = _RANDOM[9'h52][1];
        tokenCheck_counter_14 = _RANDOM[9'h52][4:2];
        shifterReg_14_0_valid = _RANDOM[9'h52][5];
        shifterReg_14_0_bits_instructionIndex = _RANDOM[9'h52][8:6];
        shifterReg_14_0_bits_decodeResult_orderReduce = _RANDOM[9'h52][9];
        shifterReg_14_0_bits_decodeResult_floatMul = _RANDOM[9'h52][10];
        shifterReg_14_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h52][12:11];
        shifterReg_14_0_bits_decodeResult_float = _RANDOM[9'h52][13];
        shifterReg_14_0_bits_decodeResult_specialSlot = _RANDOM[9'h52][14];
        shifterReg_14_0_bits_decodeResult_topUop = _RANDOM[9'h52][19:15];
        shifterReg_14_0_bits_decodeResult_popCount = _RANDOM[9'h52][20];
        shifterReg_14_0_bits_decodeResult_ffo = _RANDOM[9'h52][21];
        shifterReg_14_0_bits_decodeResult_average = _RANDOM[9'h52][22];
        shifterReg_14_0_bits_decodeResult_reverse = _RANDOM[9'h52][23];
        shifterReg_14_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h52][24];
        shifterReg_14_0_bits_decodeResult_scheduler = _RANDOM[9'h52][25];
        shifterReg_14_0_bits_decodeResult_sReadVD = _RANDOM[9'h52][26];
        shifterReg_14_0_bits_decodeResult_vtype = _RANDOM[9'h52][27];
        shifterReg_14_0_bits_decodeResult_sWrite = _RANDOM[9'h52][28];
        shifterReg_14_0_bits_decodeResult_crossRead = _RANDOM[9'h52][29];
        shifterReg_14_0_bits_decodeResult_crossWrite = _RANDOM[9'h52][30];
        shifterReg_14_0_bits_decodeResult_maskUnit = _RANDOM[9'h52][31];
        shifterReg_14_0_bits_decodeResult_special = _RANDOM[9'h53][0];
        shifterReg_14_0_bits_decodeResult_saturate = _RANDOM[9'h53][1];
        shifterReg_14_0_bits_decodeResult_vwmacc = _RANDOM[9'h53][2];
        shifterReg_14_0_bits_decodeResult_readOnly = _RANDOM[9'h53][3];
        shifterReg_14_0_bits_decodeResult_maskSource = _RANDOM[9'h53][4];
        shifterReg_14_0_bits_decodeResult_maskDestination = _RANDOM[9'h53][5];
        shifterReg_14_0_bits_decodeResult_maskLogic = _RANDOM[9'h53][6];
        shifterReg_14_0_bits_decodeResult_uop = _RANDOM[9'h53][10:7];
        shifterReg_14_0_bits_decodeResult_iota = _RANDOM[9'h53][11];
        shifterReg_14_0_bits_decodeResult_mv = _RANDOM[9'h53][12];
        shifterReg_14_0_bits_decodeResult_extend = _RANDOM[9'h53][13];
        shifterReg_14_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h53][14];
        shifterReg_14_0_bits_decodeResult_compress = _RANDOM[9'h53][15];
        shifterReg_14_0_bits_decodeResult_gather16 = _RANDOM[9'h53][16];
        shifterReg_14_0_bits_decodeResult_gather = _RANDOM[9'h53][17];
        shifterReg_14_0_bits_decodeResult_slid = _RANDOM[9'h53][18];
        shifterReg_14_0_bits_decodeResult_targetRd = _RANDOM[9'h53][19];
        shifterReg_14_0_bits_decodeResult_widenReduce = _RANDOM[9'h53][20];
        shifterReg_14_0_bits_decodeResult_red = _RANDOM[9'h53][21];
        shifterReg_14_0_bits_decodeResult_nr = _RANDOM[9'h53][22];
        shifterReg_14_0_bits_decodeResult_itype = _RANDOM[9'h53][23];
        shifterReg_14_0_bits_decodeResult_unsigned1 = _RANDOM[9'h53][24];
        shifterReg_14_0_bits_decodeResult_unsigned0 = _RANDOM[9'h53][25];
        shifterReg_14_0_bits_decodeResult_other = _RANDOM[9'h53][26];
        shifterReg_14_0_bits_decodeResult_multiCycle = _RANDOM[9'h53][27];
        shifterReg_14_0_bits_decodeResult_divider = _RANDOM[9'h53][28];
        shifterReg_14_0_bits_decodeResult_multiplier = _RANDOM[9'h53][29];
        shifterReg_14_0_bits_decodeResult_shift = _RANDOM[9'h53][30];
        shifterReg_14_0_bits_decodeResult_adder = _RANDOM[9'h53][31];
        shifterReg_14_0_bits_decodeResult_logic = _RANDOM[9'h54][0];
        shifterReg_14_0_bits_loadStore = _RANDOM[9'h54][1];
        shifterReg_14_0_bits_issueInst = _RANDOM[9'h54][2];
        shifterReg_14_0_bits_store = _RANDOM[9'h54][3];
        shifterReg_14_0_bits_special = _RANDOM[9'h54][4];
        shifterReg_14_0_bits_lsWholeReg = _RANDOM[9'h54][5];
        shifterReg_14_0_bits_vs1 = _RANDOM[9'h54][10:6];
        shifterReg_14_0_bits_vs2 = _RANDOM[9'h54][15:11];
        shifterReg_14_0_bits_vd = _RANDOM[9'h54][20:16];
        shifterReg_14_0_bits_loadStoreEEW = _RANDOM[9'h54][22:21];
        shifterReg_14_0_bits_mask = _RANDOM[9'h54][23];
        shifterReg_14_0_bits_segment = _RANDOM[9'h54][26:24];
        shifterReg_14_0_bits_readFromScalar = {_RANDOM[9'h54][31:27], _RANDOM[9'h55][26:0]};
        shifterReg_14_0_bits_csrInterface_vl = {_RANDOM[9'h55][31:27], _RANDOM[9'h56][6:0]};
        shifterReg_14_0_bits_csrInterface_vStart = _RANDOM[9'h56][18:7];
        shifterReg_14_0_bits_csrInterface_vlmul = _RANDOM[9'h56][21:19];
        shifterReg_14_0_bits_csrInterface_vSew = _RANDOM[9'h56][23:22];
        shifterReg_14_0_bits_csrInterface_vxrm = _RANDOM[9'h56][25:24];
        shifterReg_14_0_bits_csrInterface_vta = _RANDOM[9'h56][26];
        shifterReg_14_0_bits_csrInterface_vma = _RANDOM[9'h56][27];
        releasePipe_pipe_v_15 = _RANDOM[9'h56][28];
        tokenCheck_counter_15 = _RANDOM[9'h56][31:29];
        shifterReg_15_0_valid = _RANDOM[9'h57][0];
        shifterReg_15_0_bits_instructionIndex = _RANDOM[9'h57][3:1];
        shifterReg_15_0_bits_decodeResult_orderReduce = _RANDOM[9'h57][4];
        shifterReg_15_0_bits_decodeResult_floatMul = _RANDOM[9'h57][5];
        shifterReg_15_0_bits_decodeResult_fpExecutionType = _RANDOM[9'h57][7:6];
        shifterReg_15_0_bits_decodeResult_float = _RANDOM[9'h57][8];
        shifterReg_15_0_bits_decodeResult_specialSlot = _RANDOM[9'h57][9];
        shifterReg_15_0_bits_decodeResult_topUop = _RANDOM[9'h57][14:10];
        shifterReg_15_0_bits_decodeResult_popCount = _RANDOM[9'h57][15];
        shifterReg_15_0_bits_decodeResult_ffo = _RANDOM[9'h57][16];
        shifterReg_15_0_bits_decodeResult_average = _RANDOM[9'h57][17];
        shifterReg_15_0_bits_decodeResult_reverse = _RANDOM[9'h57][18];
        shifterReg_15_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h57][19];
        shifterReg_15_0_bits_decodeResult_scheduler = _RANDOM[9'h57][20];
        shifterReg_15_0_bits_decodeResult_sReadVD = _RANDOM[9'h57][21];
        shifterReg_15_0_bits_decodeResult_vtype = _RANDOM[9'h57][22];
        shifterReg_15_0_bits_decodeResult_sWrite = _RANDOM[9'h57][23];
        shifterReg_15_0_bits_decodeResult_crossRead = _RANDOM[9'h57][24];
        shifterReg_15_0_bits_decodeResult_crossWrite = _RANDOM[9'h57][25];
        shifterReg_15_0_bits_decodeResult_maskUnit = _RANDOM[9'h57][26];
        shifterReg_15_0_bits_decodeResult_special = _RANDOM[9'h57][27];
        shifterReg_15_0_bits_decodeResult_saturate = _RANDOM[9'h57][28];
        shifterReg_15_0_bits_decodeResult_vwmacc = _RANDOM[9'h57][29];
        shifterReg_15_0_bits_decodeResult_readOnly = _RANDOM[9'h57][30];
        shifterReg_15_0_bits_decodeResult_maskSource = _RANDOM[9'h57][31];
        shifterReg_15_0_bits_decodeResult_maskDestination = _RANDOM[9'h58][0];
        shifterReg_15_0_bits_decodeResult_maskLogic = _RANDOM[9'h58][1];
        shifterReg_15_0_bits_decodeResult_uop = _RANDOM[9'h58][5:2];
        shifterReg_15_0_bits_decodeResult_iota = _RANDOM[9'h58][6];
        shifterReg_15_0_bits_decodeResult_mv = _RANDOM[9'h58][7];
        shifterReg_15_0_bits_decodeResult_extend = _RANDOM[9'h58][8];
        shifterReg_15_0_bits_decodeResult_unOrderWrite = _RANDOM[9'h58][9];
        shifterReg_15_0_bits_decodeResult_compress = _RANDOM[9'h58][10];
        shifterReg_15_0_bits_decodeResult_gather16 = _RANDOM[9'h58][11];
        shifterReg_15_0_bits_decodeResult_gather = _RANDOM[9'h58][12];
        shifterReg_15_0_bits_decodeResult_slid = _RANDOM[9'h58][13];
        shifterReg_15_0_bits_decodeResult_targetRd = _RANDOM[9'h58][14];
        shifterReg_15_0_bits_decodeResult_widenReduce = _RANDOM[9'h58][15];
        shifterReg_15_0_bits_decodeResult_red = _RANDOM[9'h58][16];
        shifterReg_15_0_bits_decodeResult_nr = _RANDOM[9'h58][17];
        shifterReg_15_0_bits_decodeResult_itype = _RANDOM[9'h58][18];
        shifterReg_15_0_bits_decodeResult_unsigned1 = _RANDOM[9'h58][19];
        shifterReg_15_0_bits_decodeResult_unsigned0 = _RANDOM[9'h58][20];
        shifterReg_15_0_bits_decodeResult_other = _RANDOM[9'h58][21];
        shifterReg_15_0_bits_decodeResult_multiCycle = _RANDOM[9'h58][22];
        shifterReg_15_0_bits_decodeResult_divider = _RANDOM[9'h58][23];
        shifterReg_15_0_bits_decodeResult_multiplier = _RANDOM[9'h58][24];
        shifterReg_15_0_bits_decodeResult_shift = _RANDOM[9'h58][25];
        shifterReg_15_0_bits_decodeResult_adder = _RANDOM[9'h58][26];
        shifterReg_15_0_bits_decodeResult_logic = _RANDOM[9'h58][27];
        shifterReg_15_0_bits_loadStore = _RANDOM[9'h58][28];
        shifterReg_15_0_bits_issueInst = _RANDOM[9'h58][29];
        shifterReg_15_0_bits_store = _RANDOM[9'h58][30];
        shifterReg_15_0_bits_special = _RANDOM[9'h58][31];
        shifterReg_15_0_bits_lsWholeReg = _RANDOM[9'h59][0];
        shifterReg_15_0_bits_vs1 = _RANDOM[9'h59][5:1];
        shifterReg_15_0_bits_vs2 = _RANDOM[9'h59][10:6];
        shifterReg_15_0_bits_vd = _RANDOM[9'h59][15:11];
        shifterReg_15_0_bits_loadStoreEEW = _RANDOM[9'h59][17:16];
        shifterReg_15_0_bits_mask = _RANDOM[9'h59][18];
        shifterReg_15_0_bits_segment = _RANDOM[9'h59][21:19];
        shifterReg_15_0_bits_readFromScalar = {_RANDOM[9'h59][31:22], _RANDOM[9'h5A][21:0]};
        shifterReg_15_0_bits_csrInterface_vl = {_RANDOM[9'h5A][31:22], _RANDOM[9'h5B][1:0]};
        shifterReg_15_0_bits_csrInterface_vStart = _RANDOM[9'h5B][13:2];
        shifterReg_15_0_bits_csrInterface_vlmul = _RANDOM[9'h5B][16:14];
        shifterReg_15_0_bits_csrInterface_vSew = _RANDOM[9'h5B][18:17];
        shifterReg_15_0_bits_csrInterface_vxrm = _RANDOM[9'h5B][20:19];
        shifterReg_15_0_bits_csrInterface_vta = _RANDOM[9'h5B][21];
        shifterReg_15_0_bits_csrInterface_vma = _RANDOM[9'h5B][22];
        sinkVec_releasePipe_pipe_v = _RANDOM[9'h5B][23];
        sinkVec_tokenCheck_counter = _RANDOM[9'h5B][26:24];
        sinkVec_shifterReg_0_valid = _RANDOM[9'h5B][27];
        sinkVec_shifterReg_0_bits_vs = {_RANDOM[9'h5B][31:28], _RANDOM[9'h5C][0]};
        sinkVec_shifterReg_0_bits_readSource = _RANDOM[9'h5C][2:1];
        sinkVec_shifterReg_0_bits_offset = _RANDOM[9'h5C][4:3];
        sinkVec_shifterReg_0_bits_instructionIndex = _RANDOM[9'h5C][7:5];
        sinkVec_releasePipe_pipe_v_1 = _RANDOM[9'h5C][8];
        sinkVec_tokenCheck_counter_1 = _RANDOM[9'h5C][11:9];
        sinkVec_shifterReg_1_0_valid = _RANDOM[9'h5C][12];
        sinkVec_shifterReg_1_0_bits_vs = _RANDOM[9'h5C][17:13];
        sinkVec_shifterReg_1_0_bits_readSource = _RANDOM[9'h5C][19:18];
        sinkVec_shifterReg_1_0_bits_offset = _RANDOM[9'h5C][21:20];
        sinkVec_shifterReg_1_0_bits_instructionIndex = _RANDOM[9'h5C][24:22];
        maskUnitFirst = _RANDOM[9'h5C][25];
        accessDataValid_pipe_v = _RANDOM[9'h5C][26];
        accessDataValid_pipe_pipe_v = _RANDOM[9'h5C][27];
        shifterReg_16_0_valid = _RANDOM[9'h5C][28];
        shifterReg_16_0_bits = {_RANDOM[9'h5C][31:29], _RANDOM[9'h5D][28:0]};
        accessDataValid_pipe_v_1 = _RANDOM[9'h5D][29];
        accessDataValid_pipe_pipe_v_1 = _RANDOM[9'h5D][30];
        shifterReg_17_0_valid = _RANDOM[9'h5D][31];
        shifterReg_17_0_bits = _RANDOM[9'h5E];
        sinkVec_releasePipe_pipe_v_2 = _RANDOM[9'h5F][0];
        sinkVec_tokenCheck_counter_2 = _RANDOM[9'h5F][3:1];
        sinkVec_shifterReg_2_0_valid = _RANDOM[9'h5F][4];
        sinkVec_shifterReg_2_0_bits_vd = _RANDOM[9'h5F][9:5];
        sinkVec_shifterReg_2_0_bits_offset = _RANDOM[9'h5F][11:10];
        sinkVec_shifterReg_2_0_bits_mask = _RANDOM[9'h5F][15:12];
        sinkVec_shifterReg_2_0_bits_data = {_RANDOM[9'h5F][31:16], _RANDOM[9'h60][15:0]};
        sinkVec_shifterReg_2_0_bits_instructionIndex = _RANDOM[9'h60][19:17];
        sinkVec_releasePipe_pipe_v_3 = _RANDOM[9'h60][20];
        sinkVec_tokenCheck_counter_3 = _RANDOM[9'h60][23:21];
        sinkVec_shifterReg_3_0_valid = _RANDOM[9'h60][24];
        sinkVec_shifterReg_3_0_bits_vd = _RANDOM[9'h60][29:25];
        sinkVec_shifterReg_3_0_bits_offset = _RANDOM[9'h60][31:30];
        sinkVec_shifterReg_3_0_bits_mask = _RANDOM[9'h61][3:0];
        sinkVec_shifterReg_3_0_bits_data = {_RANDOM[9'h61][31:4], _RANDOM[9'h62][3:0]};
        sinkVec_shifterReg_3_0_bits_last = _RANDOM[9'h62][4];
        sinkVec_shifterReg_3_0_bits_instructionIndex = _RANDOM[9'h62][7:5];
        maskUnitFirst_1 = _RANDOM[9'h62][8];
        view__writeRelease_0_pipe_v = _RANDOM[9'h62][9];
        pipe_v = _RANDOM[9'h62][10];
        instructionFinishedPipe_pipe_v = _RANDOM[9'h62][11];
        instructionFinishedPipe_pipe_b = _RANDOM[9'h62][19:12];
        pipe_v_1 = _RANDOM[9'h62][20];
        pipe_b_1 = {_RANDOM[9'h62][31:21], _RANDOM[9'h63][20:0]};
        pipe_pipe_v = _RANDOM[9'h63][21];
        pipe_pipe_b = {_RANDOM[9'h63][31:22], _RANDOM[9'h64][21:0]};
        view__laneMaskSelect_0_pipe_v = _RANDOM[9'h64][22];
        view__laneMaskSelect_0_pipe_b = _RANDOM[9'h64][28:23];
        view__laneMaskSelect_0_pipe_pipe_v = _RANDOM[9'h64][29];
        view__laneMaskSelect_0_pipe_pipe_b = {_RANDOM[9'h64][31:30], _RANDOM[9'h65][3:0]};
        view__laneMaskSewSelect_0_pipe_v = _RANDOM[9'h65][4];
        view__laneMaskSewSelect_0_pipe_b = _RANDOM[9'h65][6:5];
        view__laneMaskSewSelect_0_pipe_pipe_v = _RANDOM[9'h65][7];
        view__laneMaskSewSelect_0_pipe_pipe_b = _RANDOM[9'h65][9:8];
        lsuLastPipe_pipe_v = _RANDOM[9'h65][10];
        lsuLastPipe_pipe_b = _RANDOM[9'h65][18:11];
        maskLastPipe_pipe_v = _RANDOM[9'h65][19];
        maskLastPipe_pipe_b = _RANDOM[9'h65][27:20];
        pipe_v_2 = _RANDOM[9'h65][28];
        pipe_b_2 = {_RANDOM[9'h65][31:29], _RANDOM[9'h66][2:0]};
        sinkVec_releasePipe_pipe_v_4 = _RANDOM[9'h66][3];
        sinkVec_tokenCheck_counter_4 = _RANDOM[9'h66][6:4];
        sinkVec_shifterReg_4_0_valid = _RANDOM[9'h66][7];
        sinkVec_shifterReg_4_0_bits_vs = _RANDOM[9'h66][12:8];
        sinkVec_shifterReg_4_0_bits_readSource = _RANDOM[9'h66][14:13];
        sinkVec_shifterReg_4_0_bits_offset = _RANDOM[9'h66][16:15];
        sinkVec_shifterReg_4_0_bits_instructionIndex = _RANDOM[9'h66][19:17];
        sinkVec_releasePipe_pipe_v_5 = _RANDOM[9'h66][20];
        sinkVec_tokenCheck_counter_5 = _RANDOM[9'h66][23:21];
        sinkVec_shifterReg_5_0_valid = _RANDOM[9'h66][24];
        sinkVec_shifterReg_5_0_bits_vs = _RANDOM[9'h66][29:25];
        sinkVec_shifterReg_5_0_bits_readSource = _RANDOM[9'h66][31:30];
        sinkVec_shifterReg_5_0_bits_offset = _RANDOM[9'h67][1:0];
        sinkVec_shifterReg_5_0_bits_instructionIndex = _RANDOM[9'h67][4:2];
        maskUnitFirst_2 = _RANDOM[9'h67][5];
        accessDataValid_pipe_v_2 = _RANDOM[9'h67][6];
        accessDataValid_pipe_pipe_v_2 = _RANDOM[9'h67][7];
        shifterReg_18_0_valid = _RANDOM[9'h67][8];
        shifterReg_18_0_bits = {_RANDOM[9'h67][31:9], _RANDOM[9'h68][8:0]};
        accessDataValid_pipe_v_3 = _RANDOM[9'h68][9];
        accessDataValid_pipe_pipe_v_3 = _RANDOM[9'h68][10];
        shifterReg_19_0_valid = _RANDOM[9'h68][11];
        shifterReg_19_0_bits = {_RANDOM[9'h68][31:12], _RANDOM[9'h69][11:0]};
        sinkVec_releasePipe_pipe_v_6 = _RANDOM[9'h69][12];
        sinkVec_tokenCheck_counter_6 = _RANDOM[9'h69][15:13];
        sinkVec_shifterReg_6_0_valid = _RANDOM[9'h69][16];
        sinkVec_shifterReg_6_0_bits_vd = _RANDOM[9'h69][21:17];
        sinkVec_shifterReg_6_0_bits_offset = _RANDOM[9'h69][23:22];
        sinkVec_shifterReg_6_0_bits_mask = _RANDOM[9'h69][27:24];
        sinkVec_shifterReg_6_0_bits_data = {_RANDOM[9'h69][31:28], _RANDOM[9'h6A][27:0]};
        sinkVec_shifterReg_6_0_bits_instructionIndex = _RANDOM[9'h6A][31:29];
        sinkVec_releasePipe_pipe_v_7 = _RANDOM[9'h6B][0];
        sinkVec_tokenCheck_counter_7 = _RANDOM[9'h6B][3:1];
        sinkVec_shifterReg_7_0_valid = _RANDOM[9'h6B][4];
        sinkVec_shifterReg_7_0_bits_vd = _RANDOM[9'h6B][9:5];
        sinkVec_shifterReg_7_0_bits_offset = _RANDOM[9'h6B][11:10];
        sinkVec_shifterReg_7_0_bits_mask = _RANDOM[9'h6B][15:12];
        sinkVec_shifterReg_7_0_bits_data = {_RANDOM[9'h6B][31:16], _RANDOM[9'h6C][15:0]};
        sinkVec_shifterReg_7_0_bits_last = _RANDOM[9'h6C][16];
        sinkVec_shifterReg_7_0_bits_instructionIndex = _RANDOM[9'h6C][19:17];
        maskUnitFirst_3 = _RANDOM[9'h6C][20];
        view__writeRelease_1_pipe_v = _RANDOM[9'h6C][21];
        pipe_v_3 = _RANDOM[9'h6C][22];
        instructionFinishedPipe_pipe_v_1 = _RANDOM[9'h6C][23];
        instructionFinishedPipe_pipe_b_1 = _RANDOM[9'h6C][31:24];
        pipe_v_4 = _RANDOM[9'h6D][0];
        pipe_b_4 = {_RANDOM[9'h6D][31:1], _RANDOM[9'h6E][0]};
        pipe_pipe_v_1 = _RANDOM[9'h6E][1];
        pipe_pipe_b_1 = {_RANDOM[9'h6E][31:2], _RANDOM[9'h6F][1:0]};
        view__laneMaskSelect_1_pipe_v = _RANDOM[9'h6F][2];
        view__laneMaskSelect_1_pipe_b = _RANDOM[9'h6F][8:3];
        view__laneMaskSelect_1_pipe_pipe_v = _RANDOM[9'h6F][9];
        view__laneMaskSelect_1_pipe_pipe_b = _RANDOM[9'h6F][15:10];
        view__laneMaskSewSelect_1_pipe_v = _RANDOM[9'h6F][16];
        view__laneMaskSewSelect_1_pipe_b = _RANDOM[9'h6F][18:17];
        view__laneMaskSewSelect_1_pipe_pipe_v = _RANDOM[9'h6F][19];
        view__laneMaskSewSelect_1_pipe_pipe_b = _RANDOM[9'h6F][21:20];
        lsuLastPipe_pipe_v_1 = _RANDOM[9'h6F][22];
        lsuLastPipe_pipe_b_1 = _RANDOM[9'h6F][30:23];
        maskLastPipe_pipe_v_1 = _RANDOM[9'h6F][31];
        maskLastPipe_pipe_b_1 = _RANDOM[9'h70][7:0];
        pipe_v_5 = _RANDOM[9'h70][8];
        pipe_b_5 = _RANDOM[9'h70][14:9];
        sinkVec_releasePipe_pipe_v_8 = _RANDOM[9'h70][15];
        sinkVec_tokenCheck_counter_8 = _RANDOM[9'h70][18:16];
        sinkVec_shifterReg_8_0_valid = _RANDOM[9'h70][19];
        sinkVec_shifterReg_8_0_bits_vs = _RANDOM[9'h70][24:20];
        sinkVec_shifterReg_8_0_bits_readSource = _RANDOM[9'h70][26:25];
        sinkVec_shifterReg_8_0_bits_offset = _RANDOM[9'h70][28:27];
        sinkVec_shifterReg_8_0_bits_instructionIndex = _RANDOM[9'h70][31:29];
        sinkVec_releasePipe_pipe_v_9 = _RANDOM[9'h71][0];
        sinkVec_tokenCheck_counter_9 = _RANDOM[9'h71][3:1];
        sinkVec_shifterReg_9_0_valid = _RANDOM[9'h71][4];
        sinkVec_shifterReg_9_0_bits_vs = _RANDOM[9'h71][9:5];
        sinkVec_shifterReg_9_0_bits_readSource = _RANDOM[9'h71][11:10];
        sinkVec_shifterReg_9_0_bits_offset = _RANDOM[9'h71][13:12];
        sinkVec_shifterReg_9_0_bits_instructionIndex = _RANDOM[9'h71][16:14];
        maskUnitFirst_4 = _RANDOM[9'h71][17];
        accessDataValid_pipe_v_4 = _RANDOM[9'h71][18];
        accessDataValid_pipe_pipe_v_4 = _RANDOM[9'h71][19];
        shifterReg_20_0_valid = _RANDOM[9'h71][20];
        shifterReg_20_0_bits = {_RANDOM[9'h71][31:21], _RANDOM[9'h72][20:0]};
        accessDataValid_pipe_v_5 = _RANDOM[9'h72][21];
        accessDataValid_pipe_pipe_v_5 = _RANDOM[9'h72][22];
        shifterReg_21_0_valid = _RANDOM[9'h72][23];
        shifterReg_21_0_bits = {_RANDOM[9'h72][31:24], _RANDOM[9'h73][23:0]};
        sinkVec_releasePipe_pipe_v_10 = _RANDOM[9'h73][24];
        sinkVec_tokenCheck_counter_10 = _RANDOM[9'h73][27:25];
        sinkVec_shifterReg_10_0_valid = _RANDOM[9'h73][28];
        sinkVec_shifterReg_10_0_bits_vd = {_RANDOM[9'h73][31:29], _RANDOM[9'h74][1:0]};
        sinkVec_shifterReg_10_0_bits_offset = _RANDOM[9'h74][3:2];
        sinkVec_shifterReg_10_0_bits_mask = _RANDOM[9'h74][7:4];
        sinkVec_shifterReg_10_0_bits_data = {_RANDOM[9'h74][31:8], _RANDOM[9'h75][7:0]};
        sinkVec_shifterReg_10_0_bits_instructionIndex = _RANDOM[9'h75][11:9];
        sinkVec_releasePipe_pipe_v_11 = _RANDOM[9'h75][12];
        sinkVec_tokenCheck_counter_11 = _RANDOM[9'h75][15:13];
        sinkVec_shifterReg_11_0_valid = _RANDOM[9'h75][16];
        sinkVec_shifterReg_11_0_bits_vd = _RANDOM[9'h75][21:17];
        sinkVec_shifterReg_11_0_bits_offset = _RANDOM[9'h75][23:22];
        sinkVec_shifterReg_11_0_bits_mask = _RANDOM[9'h75][27:24];
        sinkVec_shifterReg_11_0_bits_data = {_RANDOM[9'h75][31:28], _RANDOM[9'h76][27:0]};
        sinkVec_shifterReg_11_0_bits_last = _RANDOM[9'h76][28];
        sinkVec_shifterReg_11_0_bits_instructionIndex = _RANDOM[9'h76][31:29];
        maskUnitFirst_5 = _RANDOM[9'h77][0];
        view__writeRelease_2_pipe_v = _RANDOM[9'h77][1];
        pipe_v_6 = _RANDOM[9'h77][2];
        instructionFinishedPipe_pipe_v_2 = _RANDOM[9'h77][3];
        instructionFinishedPipe_pipe_b_2 = _RANDOM[9'h77][11:4];
        pipe_v_7 = _RANDOM[9'h77][12];
        pipe_b_7 = {_RANDOM[9'h77][31:13], _RANDOM[9'h78][12:0]};
        pipe_pipe_v_2 = _RANDOM[9'h78][13];
        pipe_pipe_b_2 = {_RANDOM[9'h78][31:14], _RANDOM[9'h79][13:0]};
        view__laneMaskSelect_2_pipe_v = _RANDOM[9'h79][14];
        view__laneMaskSelect_2_pipe_b = _RANDOM[9'h79][20:15];
        view__laneMaskSelect_2_pipe_pipe_v = _RANDOM[9'h79][21];
        view__laneMaskSelect_2_pipe_pipe_b = _RANDOM[9'h79][27:22];
        view__laneMaskSewSelect_2_pipe_v = _RANDOM[9'h79][28];
        view__laneMaskSewSelect_2_pipe_b = _RANDOM[9'h79][30:29];
        view__laneMaskSewSelect_2_pipe_pipe_v = _RANDOM[9'h79][31];
        view__laneMaskSewSelect_2_pipe_pipe_b = _RANDOM[9'h7A][1:0];
        lsuLastPipe_pipe_v_2 = _RANDOM[9'h7A][2];
        lsuLastPipe_pipe_b_2 = _RANDOM[9'h7A][10:3];
        maskLastPipe_pipe_v_2 = _RANDOM[9'h7A][11];
        maskLastPipe_pipe_b_2 = _RANDOM[9'h7A][19:12];
        pipe_v_8 = _RANDOM[9'h7A][20];
        pipe_b_8 = _RANDOM[9'h7A][26:21];
        sinkVec_releasePipe_pipe_v_12 = _RANDOM[9'h7A][27];
        sinkVec_tokenCheck_counter_12 = _RANDOM[9'h7A][30:28];
        sinkVec_shifterReg_12_0_valid = _RANDOM[9'h7A][31];
        sinkVec_shifterReg_12_0_bits_vs = _RANDOM[9'h7B][4:0];
        sinkVec_shifterReg_12_0_bits_readSource = _RANDOM[9'h7B][6:5];
        sinkVec_shifterReg_12_0_bits_offset = _RANDOM[9'h7B][8:7];
        sinkVec_shifterReg_12_0_bits_instructionIndex = _RANDOM[9'h7B][11:9];
        sinkVec_releasePipe_pipe_v_13 = _RANDOM[9'h7B][12];
        sinkVec_tokenCheck_counter_13 = _RANDOM[9'h7B][15:13];
        sinkVec_shifterReg_13_0_valid = _RANDOM[9'h7B][16];
        sinkVec_shifterReg_13_0_bits_vs = _RANDOM[9'h7B][21:17];
        sinkVec_shifterReg_13_0_bits_readSource = _RANDOM[9'h7B][23:22];
        sinkVec_shifterReg_13_0_bits_offset = _RANDOM[9'h7B][25:24];
        sinkVec_shifterReg_13_0_bits_instructionIndex = _RANDOM[9'h7B][28:26];
        maskUnitFirst_6 = _RANDOM[9'h7B][29];
        accessDataValid_pipe_v_6 = _RANDOM[9'h7B][30];
        accessDataValid_pipe_pipe_v_6 = _RANDOM[9'h7B][31];
        shifterReg_22_0_valid = _RANDOM[9'h7C][0];
        shifterReg_22_0_bits = {_RANDOM[9'h7C][31:1], _RANDOM[9'h7D][0]};
        accessDataValid_pipe_v_7 = _RANDOM[9'h7D][1];
        accessDataValid_pipe_pipe_v_7 = _RANDOM[9'h7D][2];
        shifterReg_23_0_valid = _RANDOM[9'h7D][3];
        shifterReg_23_0_bits = {_RANDOM[9'h7D][31:4], _RANDOM[9'h7E][3:0]};
        sinkVec_releasePipe_pipe_v_14 = _RANDOM[9'h7E][4];
        sinkVec_tokenCheck_counter_14 = _RANDOM[9'h7E][7:5];
        sinkVec_shifterReg_14_0_valid = _RANDOM[9'h7E][8];
        sinkVec_shifterReg_14_0_bits_vd = _RANDOM[9'h7E][13:9];
        sinkVec_shifterReg_14_0_bits_offset = _RANDOM[9'h7E][15:14];
        sinkVec_shifterReg_14_0_bits_mask = _RANDOM[9'h7E][19:16];
        sinkVec_shifterReg_14_0_bits_data = {_RANDOM[9'h7E][31:20], _RANDOM[9'h7F][19:0]};
        sinkVec_shifterReg_14_0_bits_instructionIndex = _RANDOM[9'h7F][23:21];
        sinkVec_releasePipe_pipe_v_15 = _RANDOM[9'h7F][24];
        sinkVec_tokenCheck_counter_15 = _RANDOM[9'h7F][27:25];
        sinkVec_shifterReg_15_0_valid = _RANDOM[9'h7F][28];
        sinkVec_shifterReg_15_0_bits_vd = {_RANDOM[9'h7F][31:29], _RANDOM[9'h80][1:0]};
        sinkVec_shifterReg_15_0_bits_offset = _RANDOM[9'h80][3:2];
        sinkVec_shifterReg_15_0_bits_mask = _RANDOM[9'h80][7:4];
        sinkVec_shifterReg_15_0_bits_data = {_RANDOM[9'h80][31:8], _RANDOM[9'h81][7:0]};
        sinkVec_shifterReg_15_0_bits_last = _RANDOM[9'h81][8];
        sinkVec_shifterReg_15_0_bits_instructionIndex = _RANDOM[9'h81][11:9];
        maskUnitFirst_7 = _RANDOM[9'h81][12];
        view__writeRelease_3_pipe_v = _RANDOM[9'h81][13];
        pipe_v_9 = _RANDOM[9'h81][14];
        instructionFinishedPipe_pipe_v_3 = _RANDOM[9'h81][15];
        instructionFinishedPipe_pipe_b_3 = _RANDOM[9'h81][23:16];
        pipe_v_10 = _RANDOM[9'h81][24];
        pipe_b_10 = {_RANDOM[9'h81][31:25], _RANDOM[9'h82][24:0]};
        pipe_pipe_v_3 = _RANDOM[9'h82][25];
        pipe_pipe_b_3 = {_RANDOM[9'h82][31:26], _RANDOM[9'h83][25:0]};
        view__laneMaskSelect_3_pipe_v = _RANDOM[9'h83][26];
        view__laneMaskSelect_3_pipe_b = {_RANDOM[9'h83][31:27], _RANDOM[9'h84][0]};
        view__laneMaskSelect_3_pipe_pipe_v = _RANDOM[9'h84][1];
        view__laneMaskSelect_3_pipe_pipe_b = _RANDOM[9'h84][7:2];
        view__laneMaskSewSelect_3_pipe_v = _RANDOM[9'h84][8];
        view__laneMaskSewSelect_3_pipe_b = _RANDOM[9'h84][10:9];
        view__laneMaskSewSelect_3_pipe_pipe_v = _RANDOM[9'h84][11];
        view__laneMaskSewSelect_3_pipe_pipe_b = _RANDOM[9'h84][13:12];
        lsuLastPipe_pipe_v_3 = _RANDOM[9'h84][14];
        lsuLastPipe_pipe_b_3 = _RANDOM[9'h84][22:15];
        maskLastPipe_pipe_v_3 = _RANDOM[9'h84][23];
        maskLastPipe_pipe_b_3 = _RANDOM[9'h84][31:24];
        pipe_v_11 = _RANDOM[9'h85][0];
        pipe_b_11 = _RANDOM[9'h85][6:1];
        sinkVec_releasePipe_pipe_v_16 = _RANDOM[9'h85][7];
        sinkVec_tokenCheck_counter_16 = _RANDOM[9'h85][10:8];
        sinkVec_shifterReg_16_0_valid = _RANDOM[9'h85][11];
        sinkVec_shifterReg_16_0_bits_vs = _RANDOM[9'h85][16:12];
        sinkVec_shifterReg_16_0_bits_readSource = _RANDOM[9'h85][18:17];
        sinkVec_shifterReg_16_0_bits_offset = _RANDOM[9'h85][20:19];
        sinkVec_shifterReg_16_0_bits_instructionIndex = _RANDOM[9'h85][23:21];
        sinkVec_releasePipe_pipe_v_17 = _RANDOM[9'h85][24];
        sinkVec_tokenCheck_counter_17 = _RANDOM[9'h85][27:25];
        sinkVec_shifterReg_17_0_valid = _RANDOM[9'h85][28];
        sinkVec_shifterReg_17_0_bits_vs = {_RANDOM[9'h85][31:29], _RANDOM[9'h86][1:0]};
        sinkVec_shifterReg_17_0_bits_readSource = _RANDOM[9'h86][3:2];
        sinkVec_shifterReg_17_0_bits_offset = _RANDOM[9'h86][5:4];
        sinkVec_shifterReg_17_0_bits_instructionIndex = _RANDOM[9'h86][8:6];
        maskUnitFirst_8 = _RANDOM[9'h86][9];
        accessDataValid_pipe_v_8 = _RANDOM[9'h86][10];
        accessDataValid_pipe_pipe_v_8 = _RANDOM[9'h86][11];
        shifterReg_24_0_valid = _RANDOM[9'h86][12];
        shifterReg_24_0_bits = {_RANDOM[9'h86][31:13], _RANDOM[9'h87][12:0]};
        accessDataValid_pipe_v_9 = _RANDOM[9'h87][13];
        accessDataValid_pipe_pipe_v_9 = _RANDOM[9'h87][14];
        shifterReg_25_0_valid = _RANDOM[9'h87][15];
        shifterReg_25_0_bits = {_RANDOM[9'h87][31:16], _RANDOM[9'h88][15:0]};
        sinkVec_releasePipe_pipe_v_18 = _RANDOM[9'h88][16];
        sinkVec_tokenCheck_counter_18 = _RANDOM[9'h88][19:17];
        sinkVec_shifterReg_18_0_valid = _RANDOM[9'h88][20];
        sinkVec_shifterReg_18_0_bits_vd = _RANDOM[9'h88][25:21];
        sinkVec_shifterReg_18_0_bits_offset = _RANDOM[9'h88][27:26];
        sinkVec_shifterReg_18_0_bits_mask = _RANDOM[9'h88][31:28];
        sinkVec_shifterReg_18_0_bits_data = _RANDOM[9'h89];
        sinkVec_shifterReg_18_0_bits_instructionIndex = _RANDOM[9'h8A][3:1];
        sinkVec_releasePipe_pipe_v_19 = _RANDOM[9'h8A][4];
        sinkVec_tokenCheck_counter_19 = _RANDOM[9'h8A][7:5];
        sinkVec_shifterReg_19_0_valid = _RANDOM[9'h8A][8];
        sinkVec_shifterReg_19_0_bits_vd = _RANDOM[9'h8A][13:9];
        sinkVec_shifterReg_19_0_bits_offset = _RANDOM[9'h8A][15:14];
        sinkVec_shifterReg_19_0_bits_mask = _RANDOM[9'h8A][19:16];
        sinkVec_shifterReg_19_0_bits_data = {_RANDOM[9'h8A][31:20], _RANDOM[9'h8B][19:0]};
        sinkVec_shifterReg_19_0_bits_last = _RANDOM[9'h8B][20];
        sinkVec_shifterReg_19_0_bits_instructionIndex = _RANDOM[9'h8B][23:21];
        maskUnitFirst_9 = _RANDOM[9'h8B][24];
        view__writeRelease_4_pipe_v = _RANDOM[9'h8B][25];
        pipe_v_12 = _RANDOM[9'h8B][26];
        instructionFinishedPipe_pipe_v_4 = _RANDOM[9'h8B][27];
        instructionFinishedPipe_pipe_b_4 = {_RANDOM[9'h8B][31:28], _RANDOM[9'h8C][3:0]};
        pipe_v_13 = _RANDOM[9'h8C][4];
        pipe_b_13 = {_RANDOM[9'h8C][31:5], _RANDOM[9'h8D][4:0]};
        pipe_pipe_v_4 = _RANDOM[9'h8D][5];
        pipe_pipe_b_4 = {_RANDOM[9'h8D][31:6], _RANDOM[9'h8E][5:0]};
        view__laneMaskSelect_4_pipe_v = _RANDOM[9'h8E][6];
        view__laneMaskSelect_4_pipe_b = _RANDOM[9'h8E][12:7];
        view__laneMaskSelect_4_pipe_pipe_v = _RANDOM[9'h8E][13];
        view__laneMaskSelect_4_pipe_pipe_b = _RANDOM[9'h8E][19:14];
        view__laneMaskSewSelect_4_pipe_v = _RANDOM[9'h8E][20];
        view__laneMaskSewSelect_4_pipe_b = _RANDOM[9'h8E][22:21];
        view__laneMaskSewSelect_4_pipe_pipe_v = _RANDOM[9'h8E][23];
        view__laneMaskSewSelect_4_pipe_pipe_b = _RANDOM[9'h8E][25:24];
        lsuLastPipe_pipe_v_4 = _RANDOM[9'h8E][26];
        lsuLastPipe_pipe_b_4 = {_RANDOM[9'h8E][31:27], _RANDOM[9'h8F][2:0]};
        maskLastPipe_pipe_v_4 = _RANDOM[9'h8F][3];
        maskLastPipe_pipe_b_4 = _RANDOM[9'h8F][11:4];
        pipe_v_14 = _RANDOM[9'h8F][12];
        pipe_b_14 = _RANDOM[9'h8F][18:13];
        sinkVec_releasePipe_pipe_v_20 = _RANDOM[9'h8F][19];
        sinkVec_tokenCheck_counter_20 = _RANDOM[9'h8F][22:20];
        sinkVec_shifterReg_20_0_valid = _RANDOM[9'h8F][23];
        sinkVec_shifterReg_20_0_bits_vs = _RANDOM[9'h8F][28:24];
        sinkVec_shifterReg_20_0_bits_readSource = _RANDOM[9'h8F][30:29];
        sinkVec_shifterReg_20_0_bits_offset = {_RANDOM[9'h8F][31], _RANDOM[9'h90][0]};
        sinkVec_shifterReg_20_0_bits_instructionIndex = _RANDOM[9'h90][3:1];
        sinkVec_releasePipe_pipe_v_21 = _RANDOM[9'h90][4];
        sinkVec_tokenCheck_counter_21 = _RANDOM[9'h90][7:5];
        sinkVec_shifterReg_21_0_valid = _RANDOM[9'h90][8];
        sinkVec_shifterReg_21_0_bits_vs = _RANDOM[9'h90][13:9];
        sinkVec_shifterReg_21_0_bits_readSource = _RANDOM[9'h90][15:14];
        sinkVec_shifterReg_21_0_bits_offset = _RANDOM[9'h90][17:16];
        sinkVec_shifterReg_21_0_bits_instructionIndex = _RANDOM[9'h90][20:18];
        maskUnitFirst_10 = _RANDOM[9'h90][21];
        accessDataValid_pipe_v_10 = _RANDOM[9'h90][22];
        accessDataValid_pipe_pipe_v_10 = _RANDOM[9'h90][23];
        shifterReg_26_0_valid = _RANDOM[9'h90][24];
        shifterReg_26_0_bits = {_RANDOM[9'h90][31:25], _RANDOM[9'h91][24:0]};
        accessDataValid_pipe_v_11 = _RANDOM[9'h91][25];
        accessDataValid_pipe_pipe_v_11 = _RANDOM[9'h91][26];
        shifterReg_27_0_valid = _RANDOM[9'h91][27];
        shifterReg_27_0_bits = {_RANDOM[9'h91][31:28], _RANDOM[9'h92][27:0]};
        sinkVec_releasePipe_pipe_v_22 = _RANDOM[9'h92][28];
        sinkVec_tokenCheck_counter_22 = _RANDOM[9'h92][31:29];
        sinkVec_shifterReg_22_0_valid = _RANDOM[9'h93][0];
        sinkVec_shifterReg_22_0_bits_vd = _RANDOM[9'h93][5:1];
        sinkVec_shifterReg_22_0_bits_offset = _RANDOM[9'h93][7:6];
        sinkVec_shifterReg_22_0_bits_mask = _RANDOM[9'h93][11:8];
        sinkVec_shifterReg_22_0_bits_data = {_RANDOM[9'h93][31:12], _RANDOM[9'h94][11:0]};
        sinkVec_shifterReg_22_0_bits_instructionIndex = _RANDOM[9'h94][15:13];
        sinkVec_releasePipe_pipe_v_23 = _RANDOM[9'h94][16];
        sinkVec_tokenCheck_counter_23 = _RANDOM[9'h94][19:17];
        sinkVec_shifterReg_23_0_valid = _RANDOM[9'h94][20];
        sinkVec_shifterReg_23_0_bits_vd = _RANDOM[9'h94][25:21];
        sinkVec_shifterReg_23_0_bits_offset = _RANDOM[9'h94][27:26];
        sinkVec_shifterReg_23_0_bits_mask = _RANDOM[9'h94][31:28];
        sinkVec_shifterReg_23_0_bits_data = _RANDOM[9'h95];
        sinkVec_shifterReg_23_0_bits_last = _RANDOM[9'h96][0];
        sinkVec_shifterReg_23_0_bits_instructionIndex = _RANDOM[9'h96][3:1];
        maskUnitFirst_11 = _RANDOM[9'h96][4];
        view__writeRelease_5_pipe_v = _RANDOM[9'h96][5];
        pipe_v_15 = _RANDOM[9'h96][6];
        instructionFinishedPipe_pipe_v_5 = _RANDOM[9'h96][7];
        instructionFinishedPipe_pipe_b_5 = _RANDOM[9'h96][15:8];
        pipe_v_16 = _RANDOM[9'h96][16];
        pipe_b_16 = {_RANDOM[9'h96][31:17], _RANDOM[9'h97][16:0]};
        pipe_pipe_v_5 = _RANDOM[9'h97][17];
        pipe_pipe_b_5 = {_RANDOM[9'h97][31:18], _RANDOM[9'h98][17:0]};
        view__laneMaskSelect_5_pipe_v = _RANDOM[9'h98][18];
        view__laneMaskSelect_5_pipe_b = _RANDOM[9'h98][24:19];
        view__laneMaskSelect_5_pipe_pipe_v = _RANDOM[9'h98][25];
        view__laneMaskSelect_5_pipe_pipe_b = _RANDOM[9'h98][31:26];
        view__laneMaskSewSelect_5_pipe_v = _RANDOM[9'h99][0];
        view__laneMaskSewSelect_5_pipe_b = _RANDOM[9'h99][2:1];
        view__laneMaskSewSelect_5_pipe_pipe_v = _RANDOM[9'h99][3];
        view__laneMaskSewSelect_5_pipe_pipe_b = _RANDOM[9'h99][5:4];
        lsuLastPipe_pipe_v_5 = _RANDOM[9'h99][6];
        lsuLastPipe_pipe_b_5 = _RANDOM[9'h99][14:7];
        maskLastPipe_pipe_v_5 = _RANDOM[9'h99][15];
        maskLastPipe_pipe_b_5 = _RANDOM[9'h99][23:16];
        pipe_v_17 = _RANDOM[9'h99][24];
        pipe_b_17 = _RANDOM[9'h99][30:25];
        sinkVec_releasePipe_pipe_v_24 = _RANDOM[9'h99][31];
        sinkVec_tokenCheck_counter_24 = _RANDOM[9'h9A][2:0];
        sinkVec_shifterReg_24_0_valid = _RANDOM[9'h9A][3];
        sinkVec_shifterReg_24_0_bits_vs = _RANDOM[9'h9A][8:4];
        sinkVec_shifterReg_24_0_bits_readSource = _RANDOM[9'h9A][10:9];
        sinkVec_shifterReg_24_0_bits_offset = _RANDOM[9'h9A][12:11];
        sinkVec_shifterReg_24_0_bits_instructionIndex = _RANDOM[9'h9A][15:13];
        sinkVec_releasePipe_pipe_v_25 = _RANDOM[9'h9A][16];
        sinkVec_tokenCheck_counter_25 = _RANDOM[9'h9A][19:17];
        sinkVec_shifterReg_25_0_valid = _RANDOM[9'h9A][20];
        sinkVec_shifterReg_25_0_bits_vs = _RANDOM[9'h9A][25:21];
        sinkVec_shifterReg_25_0_bits_readSource = _RANDOM[9'h9A][27:26];
        sinkVec_shifterReg_25_0_bits_offset = _RANDOM[9'h9A][29:28];
        sinkVec_shifterReg_25_0_bits_instructionIndex = {_RANDOM[9'h9A][31:30], _RANDOM[9'h9B][0]};
        maskUnitFirst_12 = _RANDOM[9'h9B][1];
        accessDataValid_pipe_v_12 = _RANDOM[9'h9B][2];
        accessDataValid_pipe_pipe_v_12 = _RANDOM[9'h9B][3];
        shifterReg_28_0_valid = _RANDOM[9'h9B][4];
        shifterReg_28_0_bits = {_RANDOM[9'h9B][31:5], _RANDOM[9'h9C][4:0]};
        accessDataValid_pipe_v_13 = _RANDOM[9'h9C][5];
        accessDataValid_pipe_pipe_v_13 = _RANDOM[9'h9C][6];
        shifterReg_29_0_valid = _RANDOM[9'h9C][7];
        shifterReg_29_0_bits = {_RANDOM[9'h9C][31:8], _RANDOM[9'h9D][7:0]};
        sinkVec_releasePipe_pipe_v_26 = _RANDOM[9'h9D][8];
        sinkVec_tokenCheck_counter_26 = _RANDOM[9'h9D][11:9];
        sinkVec_shifterReg_26_0_valid = _RANDOM[9'h9D][12];
        sinkVec_shifterReg_26_0_bits_vd = _RANDOM[9'h9D][17:13];
        sinkVec_shifterReg_26_0_bits_offset = _RANDOM[9'h9D][19:18];
        sinkVec_shifterReg_26_0_bits_mask = _RANDOM[9'h9D][23:20];
        sinkVec_shifterReg_26_0_bits_data = {_RANDOM[9'h9D][31:24], _RANDOM[9'h9E][23:0]};
        sinkVec_shifterReg_26_0_bits_instructionIndex = _RANDOM[9'h9E][27:25];
        sinkVec_releasePipe_pipe_v_27 = _RANDOM[9'h9E][28];
        sinkVec_tokenCheck_counter_27 = _RANDOM[9'h9E][31:29];
        sinkVec_shifterReg_27_0_valid = _RANDOM[9'h9F][0];
        sinkVec_shifterReg_27_0_bits_vd = _RANDOM[9'h9F][5:1];
        sinkVec_shifterReg_27_0_bits_offset = _RANDOM[9'h9F][7:6];
        sinkVec_shifterReg_27_0_bits_mask = _RANDOM[9'h9F][11:8];
        sinkVec_shifterReg_27_0_bits_data = {_RANDOM[9'h9F][31:12], _RANDOM[9'hA0][11:0]};
        sinkVec_shifterReg_27_0_bits_last = _RANDOM[9'hA0][12];
        sinkVec_shifterReg_27_0_bits_instructionIndex = _RANDOM[9'hA0][15:13];
        maskUnitFirst_13 = _RANDOM[9'hA0][16];
        view__writeRelease_6_pipe_v = _RANDOM[9'hA0][17];
        pipe_v_18 = _RANDOM[9'hA0][18];
        instructionFinishedPipe_pipe_v_6 = _RANDOM[9'hA0][19];
        instructionFinishedPipe_pipe_b_6 = _RANDOM[9'hA0][27:20];
        pipe_v_19 = _RANDOM[9'hA0][28];
        pipe_b_19 = {_RANDOM[9'hA0][31:29], _RANDOM[9'hA1][28:0]};
        pipe_pipe_v_6 = _RANDOM[9'hA1][29];
        pipe_pipe_b_6 = {_RANDOM[9'hA1][31:30], _RANDOM[9'hA2][29:0]};
        view__laneMaskSelect_6_pipe_v = _RANDOM[9'hA2][30];
        view__laneMaskSelect_6_pipe_b = {_RANDOM[9'hA2][31], _RANDOM[9'hA3][4:0]};
        view__laneMaskSelect_6_pipe_pipe_v = _RANDOM[9'hA3][5];
        view__laneMaskSelect_6_pipe_pipe_b = _RANDOM[9'hA3][11:6];
        view__laneMaskSewSelect_6_pipe_v = _RANDOM[9'hA3][12];
        view__laneMaskSewSelect_6_pipe_b = _RANDOM[9'hA3][14:13];
        view__laneMaskSewSelect_6_pipe_pipe_v = _RANDOM[9'hA3][15];
        view__laneMaskSewSelect_6_pipe_pipe_b = _RANDOM[9'hA3][17:16];
        lsuLastPipe_pipe_v_6 = _RANDOM[9'hA3][18];
        lsuLastPipe_pipe_b_6 = _RANDOM[9'hA3][26:19];
        maskLastPipe_pipe_v_6 = _RANDOM[9'hA3][27];
        maskLastPipe_pipe_b_6 = {_RANDOM[9'hA3][31:28], _RANDOM[9'hA4][3:0]};
        pipe_v_20 = _RANDOM[9'hA4][4];
        pipe_b_20 = _RANDOM[9'hA4][10:5];
        sinkVec_releasePipe_pipe_v_28 = _RANDOM[9'hA4][11];
        sinkVec_tokenCheck_counter_28 = _RANDOM[9'hA4][14:12];
        sinkVec_shifterReg_28_0_valid = _RANDOM[9'hA4][15];
        sinkVec_shifterReg_28_0_bits_vs = _RANDOM[9'hA4][20:16];
        sinkVec_shifterReg_28_0_bits_readSource = _RANDOM[9'hA4][22:21];
        sinkVec_shifterReg_28_0_bits_offset = _RANDOM[9'hA4][24:23];
        sinkVec_shifterReg_28_0_bits_instructionIndex = _RANDOM[9'hA4][27:25];
        sinkVec_releasePipe_pipe_v_29 = _RANDOM[9'hA4][28];
        sinkVec_tokenCheck_counter_29 = _RANDOM[9'hA4][31:29];
        sinkVec_shifterReg_29_0_valid = _RANDOM[9'hA5][0];
        sinkVec_shifterReg_29_0_bits_vs = _RANDOM[9'hA5][5:1];
        sinkVec_shifterReg_29_0_bits_readSource = _RANDOM[9'hA5][7:6];
        sinkVec_shifterReg_29_0_bits_offset = _RANDOM[9'hA5][9:8];
        sinkVec_shifterReg_29_0_bits_instructionIndex = _RANDOM[9'hA5][12:10];
        maskUnitFirst_14 = _RANDOM[9'hA5][13];
        accessDataValid_pipe_v_14 = _RANDOM[9'hA5][14];
        accessDataValid_pipe_pipe_v_14 = _RANDOM[9'hA5][15];
        shifterReg_30_0_valid = _RANDOM[9'hA5][16];
        shifterReg_30_0_bits = {_RANDOM[9'hA5][31:17], _RANDOM[9'hA6][16:0]};
        accessDataValid_pipe_v_15 = _RANDOM[9'hA6][17];
        accessDataValid_pipe_pipe_v_15 = _RANDOM[9'hA6][18];
        shifterReg_31_0_valid = _RANDOM[9'hA6][19];
        shifterReg_31_0_bits = {_RANDOM[9'hA6][31:20], _RANDOM[9'hA7][19:0]};
        sinkVec_releasePipe_pipe_v_30 = _RANDOM[9'hA7][20];
        sinkVec_tokenCheck_counter_30 = _RANDOM[9'hA7][23:21];
        sinkVec_shifterReg_30_0_valid = _RANDOM[9'hA7][24];
        sinkVec_shifterReg_30_0_bits_vd = _RANDOM[9'hA7][29:25];
        sinkVec_shifterReg_30_0_bits_offset = _RANDOM[9'hA7][31:30];
        sinkVec_shifterReg_30_0_bits_mask = _RANDOM[9'hA8][3:0];
        sinkVec_shifterReg_30_0_bits_data = {_RANDOM[9'hA8][31:4], _RANDOM[9'hA9][3:0]};
        sinkVec_shifterReg_30_0_bits_instructionIndex = _RANDOM[9'hA9][7:5];
        sinkVec_releasePipe_pipe_v_31 = _RANDOM[9'hA9][8];
        sinkVec_tokenCheck_counter_31 = _RANDOM[9'hA9][11:9];
        sinkVec_shifterReg_31_0_valid = _RANDOM[9'hA9][12];
        sinkVec_shifterReg_31_0_bits_vd = _RANDOM[9'hA9][17:13];
        sinkVec_shifterReg_31_0_bits_offset = _RANDOM[9'hA9][19:18];
        sinkVec_shifterReg_31_0_bits_mask = _RANDOM[9'hA9][23:20];
        sinkVec_shifterReg_31_0_bits_data = {_RANDOM[9'hA9][31:24], _RANDOM[9'hAA][23:0]};
        sinkVec_shifterReg_31_0_bits_last = _RANDOM[9'hAA][24];
        sinkVec_shifterReg_31_0_bits_instructionIndex = _RANDOM[9'hAA][27:25];
        maskUnitFirst_15 = _RANDOM[9'hAA][28];
        view__writeRelease_7_pipe_v = _RANDOM[9'hAA][29];
        pipe_v_21 = _RANDOM[9'hAA][30];
        instructionFinishedPipe_pipe_v_7 = _RANDOM[9'hAA][31];
        instructionFinishedPipe_pipe_b_7 = _RANDOM[9'hAB][7:0];
        pipe_v_22 = _RANDOM[9'hAB][8];
        pipe_b_22 = {_RANDOM[9'hAB][31:9], _RANDOM[9'hAC][8:0]};
        pipe_pipe_v_7 = _RANDOM[9'hAC][9];
        pipe_pipe_b_7 = {_RANDOM[9'hAC][31:10], _RANDOM[9'hAD][9:0]};
        view__laneMaskSelect_7_pipe_v = _RANDOM[9'hAD][10];
        view__laneMaskSelect_7_pipe_b = _RANDOM[9'hAD][16:11];
        view__laneMaskSelect_7_pipe_pipe_v = _RANDOM[9'hAD][17];
        view__laneMaskSelect_7_pipe_pipe_b = _RANDOM[9'hAD][23:18];
        view__laneMaskSewSelect_7_pipe_v = _RANDOM[9'hAD][24];
        view__laneMaskSewSelect_7_pipe_b = _RANDOM[9'hAD][26:25];
        view__laneMaskSewSelect_7_pipe_pipe_v = _RANDOM[9'hAD][27];
        view__laneMaskSewSelect_7_pipe_pipe_b = _RANDOM[9'hAD][29:28];
        lsuLastPipe_pipe_v_7 = _RANDOM[9'hAD][30];
        lsuLastPipe_pipe_b_7 = {_RANDOM[9'hAD][31], _RANDOM[9'hAE][6:0]};
        maskLastPipe_pipe_v_7 = _RANDOM[9'hAE][7];
        maskLastPipe_pipe_b_7 = _RANDOM[9'hAE][15:8];
        pipe_v_23 = _RANDOM[9'hAE][16];
        pipe_b_23 = _RANDOM[9'hAE][22:17];
        sinkVec_releasePipe_pipe_v_32 = _RANDOM[9'hAE][23];
        sinkVec_tokenCheck_counter_32 = _RANDOM[9'hAE][26:24];
        sinkVec_shifterReg_32_0_valid = _RANDOM[9'hAE][27];
        sinkVec_shifterReg_32_0_bits_vs = {_RANDOM[9'hAE][31:28], _RANDOM[9'hAF][0]};
        sinkVec_shifterReg_32_0_bits_readSource = _RANDOM[9'hAF][2:1];
        sinkVec_shifterReg_32_0_bits_offset = _RANDOM[9'hAF][4:3];
        sinkVec_shifterReg_32_0_bits_instructionIndex = _RANDOM[9'hAF][7:5];
        sinkVec_releasePipe_pipe_v_33 = _RANDOM[9'hAF][8];
        sinkVec_tokenCheck_counter_33 = _RANDOM[9'hAF][11:9];
        sinkVec_shifterReg_33_0_valid = _RANDOM[9'hAF][12];
        sinkVec_shifterReg_33_0_bits_vs = _RANDOM[9'hAF][17:13];
        sinkVec_shifterReg_33_0_bits_readSource = _RANDOM[9'hAF][19:18];
        sinkVec_shifterReg_33_0_bits_offset = _RANDOM[9'hAF][21:20];
        sinkVec_shifterReg_33_0_bits_instructionIndex = _RANDOM[9'hAF][24:22];
        maskUnitFirst_16 = _RANDOM[9'hAF][25];
        accessDataValid_pipe_v_16 = _RANDOM[9'hAF][26];
        accessDataValid_pipe_pipe_v_16 = _RANDOM[9'hAF][27];
        shifterReg_32_0_valid = _RANDOM[9'hAF][28];
        shifterReg_32_0_bits = {_RANDOM[9'hAF][31:29], _RANDOM[9'hB0][28:0]};
        accessDataValid_pipe_v_17 = _RANDOM[9'hB0][29];
        accessDataValid_pipe_pipe_v_17 = _RANDOM[9'hB0][30];
        shifterReg_33_0_valid = _RANDOM[9'hB0][31];
        shifterReg_33_0_bits = _RANDOM[9'hB1];
        sinkVec_releasePipe_pipe_v_34 = _RANDOM[9'hB2][0];
        sinkVec_tokenCheck_counter_34 = _RANDOM[9'hB2][3:1];
        sinkVec_shifterReg_34_0_valid = _RANDOM[9'hB2][4];
        sinkVec_shifterReg_34_0_bits_vd = _RANDOM[9'hB2][9:5];
        sinkVec_shifterReg_34_0_bits_offset = _RANDOM[9'hB2][11:10];
        sinkVec_shifterReg_34_0_bits_mask = _RANDOM[9'hB2][15:12];
        sinkVec_shifterReg_34_0_bits_data = {_RANDOM[9'hB2][31:16], _RANDOM[9'hB3][15:0]};
        sinkVec_shifterReg_34_0_bits_instructionIndex = _RANDOM[9'hB3][19:17];
        sinkVec_releasePipe_pipe_v_35 = _RANDOM[9'hB3][20];
        sinkVec_tokenCheck_counter_35 = _RANDOM[9'hB3][23:21];
        sinkVec_shifterReg_35_0_valid = _RANDOM[9'hB3][24];
        sinkVec_shifterReg_35_0_bits_vd = _RANDOM[9'hB3][29:25];
        sinkVec_shifterReg_35_0_bits_offset = _RANDOM[9'hB3][31:30];
        sinkVec_shifterReg_35_0_bits_mask = _RANDOM[9'hB4][3:0];
        sinkVec_shifterReg_35_0_bits_data = {_RANDOM[9'hB4][31:4], _RANDOM[9'hB5][3:0]};
        sinkVec_shifterReg_35_0_bits_last = _RANDOM[9'hB5][4];
        sinkVec_shifterReg_35_0_bits_instructionIndex = _RANDOM[9'hB5][7:5];
        maskUnitFirst_17 = _RANDOM[9'hB5][8];
        view__writeRelease_8_pipe_v = _RANDOM[9'hB5][9];
        pipe_v_24 = _RANDOM[9'hB5][10];
        instructionFinishedPipe_pipe_v_8 = _RANDOM[9'hB5][11];
        instructionFinishedPipe_pipe_b_8 = _RANDOM[9'hB5][19:12];
        pipe_v_25 = _RANDOM[9'hB5][20];
        pipe_b_25 = {_RANDOM[9'hB5][31:21], _RANDOM[9'hB6][20:0]};
        pipe_pipe_v_8 = _RANDOM[9'hB6][21];
        pipe_pipe_b_8 = {_RANDOM[9'hB6][31:22], _RANDOM[9'hB7][21:0]};
        view__laneMaskSelect_8_pipe_v = _RANDOM[9'hB7][22];
        view__laneMaskSelect_8_pipe_b = _RANDOM[9'hB7][28:23];
        view__laneMaskSelect_8_pipe_pipe_v = _RANDOM[9'hB7][29];
        view__laneMaskSelect_8_pipe_pipe_b = {_RANDOM[9'hB7][31:30], _RANDOM[9'hB8][3:0]};
        view__laneMaskSewSelect_8_pipe_v = _RANDOM[9'hB8][4];
        view__laneMaskSewSelect_8_pipe_b = _RANDOM[9'hB8][6:5];
        view__laneMaskSewSelect_8_pipe_pipe_v = _RANDOM[9'hB8][7];
        view__laneMaskSewSelect_8_pipe_pipe_b = _RANDOM[9'hB8][9:8];
        lsuLastPipe_pipe_v_8 = _RANDOM[9'hB8][10];
        lsuLastPipe_pipe_b_8 = _RANDOM[9'hB8][18:11];
        maskLastPipe_pipe_v_8 = _RANDOM[9'hB8][19];
        maskLastPipe_pipe_b_8 = _RANDOM[9'hB8][27:20];
        pipe_v_26 = _RANDOM[9'hB8][28];
        pipe_b_26 = {_RANDOM[9'hB8][31:29], _RANDOM[9'hB9][2:0]};
        sinkVec_releasePipe_pipe_v_36 = _RANDOM[9'hB9][3];
        sinkVec_tokenCheck_counter_36 = _RANDOM[9'hB9][6:4];
        sinkVec_shifterReg_36_0_valid = _RANDOM[9'hB9][7];
        sinkVec_shifterReg_36_0_bits_vs = _RANDOM[9'hB9][12:8];
        sinkVec_shifterReg_36_0_bits_readSource = _RANDOM[9'hB9][14:13];
        sinkVec_shifterReg_36_0_bits_offset = _RANDOM[9'hB9][16:15];
        sinkVec_shifterReg_36_0_bits_instructionIndex = _RANDOM[9'hB9][19:17];
        sinkVec_releasePipe_pipe_v_37 = _RANDOM[9'hB9][20];
        sinkVec_tokenCheck_counter_37 = _RANDOM[9'hB9][23:21];
        sinkVec_shifterReg_37_0_valid = _RANDOM[9'hB9][24];
        sinkVec_shifterReg_37_0_bits_vs = _RANDOM[9'hB9][29:25];
        sinkVec_shifterReg_37_0_bits_readSource = _RANDOM[9'hB9][31:30];
        sinkVec_shifterReg_37_0_bits_offset = _RANDOM[9'hBA][1:0];
        sinkVec_shifterReg_37_0_bits_instructionIndex = _RANDOM[9'hBA][4:2];
        maskUnitFirst_18 = _RANDOM[9'hBA][5];
        accessDataValid_pipe_v_18 = _RANDOM[9'hBA][6];
        accessDataValid_pipe_pipe_v_18 = _RANDOM[9'hBA][7];
        shifterReg_34_0_valid = _RANDOM[9'hBA][8];
        shifterReg_34_0_bits = {_RANDOM[9'hBA][31:9], _RANDOM[9'hBB][8:0]};
        accessDataValid_pipe_v_19 = _RANDOM[9'hBB][9];
        accessDataValid_pipe_pipe_v_19 = _RANDOM[9'hBB][10];
        shifterReg_35_0_valid = _RANDOM[9'hBB][11];
        shifterReg_35_0_bits = {_RANDOM[9'hBB][31:12], _RANDOM[9'hBC][11:0]};
        sinkVec_releasePipe_pipe_v_38 = _RANDOM[9'hBC][12];
        sinkVec_tokenCheck_counter_38 = _RANDOM[9'hBC][15:13];
        sinkVec_shifterReg_38_0_valid = _RANDOM[9'hBC][16];
        sinkVec_shifterReg_38_0_bits_vd = _RANDOM[9'hBC][21:17];
        sinkVec_shifterReg_38_0_bits_offset = _RANDOM[9'hBC][23:22];
        sinkVec_shifterReg_38_0_bits_mask = _RANDOM[9'hBC][27:24];
        sinkVec_shifterReg_38_0_bits_data = {_RANDOM[9'hBC][31:28], _RANDOM[9'hBD][27:0]};
        sinkVec_shifterReg_38_0_bits_instructionIndex = _RANDOM[9'hBD][31:29];
        sinkVec_releasePipe_pipe_v_39 = _RANDOM[9'hBE][0];
        sinkVec_tokenCheck_counter_39 = _RANDOM[9'hBE][3:1];
        sinkVec_shifterReg_39_0_valid = _RANDOM[9'hBE][4];
        sinkVec_shifterReg_39_0_bits_vd = _RANDOM[9'hBE][9:5];
        sinkVec_shifterReg_39_0_bits_offset = _RANDOM[9'hBE][11:10];
        sinkVec_shifterReg_39_0_bits_mask = _RANDOM[9'hBE][15:12];
        sinkVec_shifterReg_39_0_bits_data = {_RANDOM[9'hBE][31:16], _RANDOM[9'hBF][15:0]};
        sinkVec_shifterReg_39_0_bits_last = _RANDOM[9'hBF][16];
        sinkVec_shifterReg_39_0_bits_instructionIndex = _RANDOM[9'hBF][19:17];
        maskUnitFirst_19 = _RANDOM[9'hBF][20];
        view__writeRelease_9_pipe_v = _RANDOM[9'hBF][21];
        pipe_v_27 = _RANDOM[9'hBF][22];
        instructionFinishedPipe_pipe_v_9 = _RANDOM[9'hBF][23];
        instructionFinishedPipe_pipe_b_9 = _RANDOM[9'hBF][31:24];
        pipe_v_28 = _RANDOM[9'hC0][0];
        pipe_b_28 = {_RANDOM[9'hC0][31:1], _RANDOM[9'hC1][0]};
        pipe_pipe_v_9 = _RANDOM[9'hC1][1];
        pipe_pipe_b_9 = {_RANDOM[9'hC1][31:2], _RANDOM[9'hC2][1:0]};
        view__laneMaskSelect_9_pipe_v = _RANDOM[9'hC2][2];
        view__laneMaskSelect_9_pipe_b = _RANDOM[9'hC2][8:3];
        view__laneMaskSelect_9_pipe_pipe_v = _RANDOM[9'hC2][9];
        view__laneMaskSelect_9_pipe_pipe_b = _RANDOM[9'hC2][15:10];
        view__laneMaskSewSelect_9_pipe_v = _RANDOM[9'hC2][16];
        view__laneMaskSewSelect_9_pipe_b = _RANDOM[9'hC2][18:17];
        view__laneMaskSewSelect_9_pipe_pipe_v = _RANDOM[9'hC2][19];
        view__laneMaskSewSelect_9_pipe_pipe_b = _RANDOM[9'hC2][21:20];
        lsuLastPipe_pipe_v_9 = _RANDOM[9'hC2][22];
        lsuLastPipe_pipe_b_9 = _RANDOM[9'hC2][30:23];
        maskLastPipe_pipe_v_9 = _RANDOM[9'hC2][31];
        maskLastPipe_pipe_b_9 = _RANDOM[9'hC3][7:0];
        pipe_v_29 = _RANDOM[9'hC3][8];
        pipe_b_29 = _RANDOM[9'hC3][14:9];
        sinkVec_releasePipe_pipe_v_40 = _RANDOM[9'hC3][15];
        sinkVec_tokenCheck_counter_40 = _RANDOM[9'hC3][18:16];
        sinkVec_shifterReg_40_0_valid = _RANDOM[9'hC3][19];
        sinkVec_shifterReg_40_0_bits_vs = _RANDOM[9'hC3][24:20];
        sinkVec_shifterReg_40_0_bits_readSource = _RANDOM[9'hC3][26:25];
        sinkVec_shifterReg_40_0_bits_offset = _RANDOM[9'hC3][28:27];
        sinkVec_shifterReg_40_0_bits_instructionIndex = _RANDOM[9'hC3][31:29];
        sinkVec_releasePipe_pipe_v_41 = _RANDOM[9'hC4][0];
        sinkVec_tokenCheck_counter_41 = _RANDOM[9'hC4][3:1];
        sinkVec_shifterReg_41_0_valid = _RANDOM[9'hC4][4];
        sinkVec_shifterReg_41_0_bits_vs = _RANDOM[9'hC4][9:5];
        sinkVec_shifterReg_41_0_bits_readSource = _RANDOM[9'hC4][11:10];
        sinkVec_shifterReg_41_0_bits_offset = _RANDOM[9'hC4][13:12];
        sinkVec_shifterReg_41_0_bits_instructionIndex = _RANDOM[9'hC4][16:14];
        maskUnitFirst_20 = _RANDOM[9'hC4][17];
        accessDataValid_pipe_v_20 = _RANDOM[9'hC4][18];
        accessDataValid_pipe_pipe_v_20 = _RANDOM[9'hC4][19];
        shifterReg_36_0_valid = _RANDOM[9'hC4][20];
        shifterReg_36_0_bits = {_RANDOM[9'hC4][31:21], _RANDOM[9'hC5][20:0]};
        accessDataValid_pipe_v_21 = _RANDOM[9'hC5][21];
        accessDataValid_pipe_pipe_v_21 = _RANDOM[9'hC5][22];
        shifterReg_37_0_valid = _RANDOM[9'hC5][23];
        shifterReg_37_0_bits = {_RANDOM[9'hC5][31:24], _RANDOM[9'hC6][23:0]};
        sinkVec_releasePipe_pipe_v_42 = _RANDOM[9'hC6][24];
        sinkVec_tokenCheck_counter_42 = _RANDOM[9'hC6][27:25];
        sinkVec_shifterReg_42_0_valid = _RANDOM[9'hC6][28];
        sinkVec_shifterReg_42_0_bits_vd = {_RANDOM[9'hC6][31:29], _RANDOM[9'hC7][1:0]};
        sinkVec_shifterReg_42_0_bits_offset = _RANDOM[9'hC7][3:2];
        sinkVec_shifterReg_42_0_bits_mask = _RANDOM[9'hC7][7:4];
        sinkVec_shifterReg_42_0_bits_data = {_RANDOM[9'hC7][31:8], _RANDOM[9'hC8][7:0]};
        sinkVec_shifterReg_42_0_bits_instructionIndex = _RANDOM[9'hC8][11:9];
        sinkVec_releasePipe_pipe_v_43 = _RANDOM[9'hC8][12];
        sinkVec_tokenCheck_counter_43 = _RANDOM[9'hC8][15:13];
        sinkVec_shifterReg_43_0_valid = _RANDOM[9'hC8][16];
        sinkVec_shifterReg_43_0_bits_vd = _RANDOM[9'hC8][21:17];
        sinkVec_shifterReg_43_0_bits_offset = _RANDOM[9'hC8][23:22];
        sinkVec_shifterReg_43_0_bits_mask = _RANDOM[9'hC8][27:24];
        sinkVec_shifterReg_43_0_bits_data = {_RANDOM[9'hC8][31:28], _RANDOM[9'hC9][27:0]};
        sinkVec_shifterReg_43_0_bits_last = _RANDOM[9'hC9][28];
        sinkVec_shifterReg_43_0_bits_instructionIndex = _RANDOM[9'hC9][31:29];
        maskUnitFirst_21 = _RANDOM[9'hCA][0];
        view__writeRelease_10_pipe_v = _RANDOM[9'hCA][1];
        pipe_v_30 = _RANDOM[9'hCA][2];
        instructionFinishedPipe_pipe_v_10 = _RANDOM[9'hCA][3];
        instructionFinishedPipe_pipe_b_10 = _RANDOM[9'hCA][11:4];
        pipe_v_31 = _RANDOM[9'hCA][12];
        pipe_b_31 = {_RANDOM[9'hCA][31:13], _RANDOM[9'hCB][12:0]};
        pipe_pipe_v_10 = _RANDOM[9'hCB][13];
        pipe_pipe_b_10 = {_RANDOM[9'hCB][31:14], _RANDOM[9'hCC][13:0]};
        view__laneMaskSelect_10_pipe_v = _RANDOM[9'hCC][14];
        view__laneMaskSelect_10_pipe_b = _RANDOM[9'hCC][20:15];
        view__laneMaskSelect_10_pipe_pipe_v = _RANDOM[9'hCC][21];
        view__laneMaskSelect_10_pipe_pipe_b = _RANDOM[9'hCC][27:22];
        view__laneMaskSewSelect_10_pipe_v = _RANDOM[9'hCC][28];
        view__laneMaskSewSelect_10_pipe_b = _RANDOM[9'hCC][30:29];
        view__laneMaskSewSelect_10_pipe_pipe_v = _RANDOM[9'hCC][31];
        view__laneMaskSewSelect_10_pipe_pipe_b = _RANDOM[9'hCD][1:0];
        lsuLastPipe_pipe_v_10 = _RANDOM[9'hCD][2];
        lsuLastPipe_pipe_b_10 = _RANDOM[9'hCD][10:3];
        maskLastPipe_pipe_v_10 = _RANDOM[9'hCD][11];
        maskLastPipe_pipe_b_10 = _RANDOM[9'hCD][19:12];
        pipe_v_32 = _RANDOM[9'hCD][20];
        pipe_b_32 = _RANDOM[9'hCD][26:21];
        sinkVec_releasePipe_pipe_v_44 = _RANDOM[9'hCD][27];
        sinkVec_tokenCheck_counter_44 = _RANDOM[9'hCD][30:28];
        sinkVec_shifterReg_44_0_valid = _RANDOM[9'hCD][31];
        sinkVec_shifterReg_44_0_bits_vs = _RANDOM[9'hCE][4:0];
        sinkVec_shifterReg_44_0_bits_readSource = _RANDOM[9'hCE][6:5];
        sinkVec_shifterReg_44_0_bits_offset = _RANDOM[9'hCE][8:7];
        sinkVec_shifterReg_44_0_bits_instructionIndex = _RANDOM[9'hCE][11:9];
        sinkVec_releasePipe_pipe_v_45 = _RANDOM[9'hCE][12];
        sinkVec_tokenCheck_counter_45 = _RANDOM[9'hCE][15:13];
        sinkVec_shifterReg_45_0_valid = _RANDOM[9'hCE][16];
        sinkVec_shifterReg_45_0_bits_vs = _RANDOM[9'hCE][21:17];
        sinkVec_shifterReg_45_0_bits_readSource = _RANDOM[9'hCE][23:22];
        sinkVec_shifterReg_45_0_bits_offset = _RANDOM[9'hCE][25:24];
        sinkVec_shifterReg_45_0_bits_instructionIndex = _RANDOM[9'hCE][28:26];
        maskUnitFirst_22 = _RANDOM[9'hCE][29];
        accessDataValid_pipe_v_22 = _RANDOM[9'hCE][30];
        accessDataValid_pipe_pipe_v_22 = _RANDOM[9'hCE][31];
        shifterReg_38_0_valid = _RANDOM[9'hCF][0];
        shifterReg_38_0_bits = {_RANDOM[9'hCF][31:1], _RANDOM[9'hD0][0]};
        accessDataValid_pipe_v_23 = _RANDOM[9'hD0][1];
        accessDataValid_pipe_pipe_v_23 = _RANDOM[9'hD0][2];
        shifterReg_39_0_valid = _RANDOM[9'hD0][3];
        shifterReg_39_0_bits = {_RANDOM[9'hD0][31:4], _RANDOM[9'hD1][3:0]};
        sinkVec_releasePipe_pipe_v_46 = _RANDOM[9'hD1][4];
        sinkVec_tokenCheck_counter_46 = _RANDOM[9'hD1][7:5];
        sinkVec_shifterReg_46_0_valid = _RANDOM[9'hD1][8];
        sinkVec_shifterReg_46_0_bits_vd = _RANDOM[9'hD1][13:9];
        sinkVec_shifterReg_46_0_bits_offset = _RANDOM[9'hD1][15:14];
        sinkVec_shifterReg_46_0_bits_mask = _RANDOM[9'hD1][19:16];
        sinkVec_shifterReg_46_0_bits_data = {_RANDOM[9'hD1][31:20], _RANDOM[9'hD2][19:0]};
        sinkVec_shifterReg_46_0_bits_instructionIndex = _RANDOM[9'hD2][23:21];
        sinkVec_releasePipe_pipe_v_47 = _RANDOM[9'hD2][24];
        sinkVec_tokenCheck_counter_47 = _RANDOM[9'hD2][27:25];
        sinkVec_shifterReg_47_0_valid = _RANDOM[9'hD2][28];
        sinkVec_shifterReg_47_0_bits_vd = {_RANDOM[9'hD2][31:29], _RANDOM[9'hD3][1:0]};
        sinkVec_shifterReg_47_0_bits_offset = _RANDOM[9'hD3][3:2];
        sinkVec_shifterReg_47_0_bits_mask = _RANDOM[9'hD3][7:4];
        sinkVec_shifterReg_47_0_bits_data = {_RANDOM[9'hD3][31:8], _RANDOM[9'hD4][7:0]};
        sinkVec_shifterReg_47_0_bits_last = _RANDOM[9'hD4][8];
        sinkVec_shifterReg_47_0_bits_instructionIndex = _RANDOM[9'hD4][11:9];
        maskUnitFirst_23 = _RANDOM[9'hD4][12];
        view__writeRelease_11_pipe_v = _RANDOM[9'hD4][13];
        pipe_v_33 = _RANDOM[9'hD4][14];
        instructionFinishedPipe_pipe_v_11 = _RANDOM[9'hD4][15];
        instructionFinishedPipe_pipe_b_11 = _RANDOM[9'hD4][23:16];
        pipe_v_34 = _RANDOM[9'hD4][24];
        pipe_b_34 = {_RANDOM[9'hD4][31:25], _RANDOM[9'hD5][24:0]};
        pipe_pipe_v_11 = _RANDOM[9'hD5][25];
        pipe_pipe_b_11 = {_RANDOM[9'hD5][31:26], _RANDOM[9'hD6][25:0]};
        view__laneMaskSelect_11_pipe_v = _RANDOM[9'hD6][26];
        view__laneMaskSelect_11_pipe_b = {_RANDOM[9'hD6][31:27], _RANDOM[9'hD7][0]};
        view__laneMaskSelect_11_pipe_pipe_v = _RANDOM[9'hD7][1];
        view__laneMaskSelect_11_pipe_pipe_b = _RANDOM[9'hD7][7:2];
        view__laneMaskSewSelect_11_pipe_v = _RANDOM[9'hD7][8];
        view__laneMaskSewSelect_11_pipe_b = _RANDOM[9'hD7][10:9];
        view__laneMaskSewSelect_11_pipe_pipe_v = _RANDOM[9'hD7][11];
        view__laneMaskSewSelect_11_pipe_pipe_b = _RANDOM[9'hD7][13:12];
        lsuLastPipe_pipe_v_11 = _RANDOM[9'hD7][14];
        lsuLastPipe_pipe_b_11 = _RANDOM[9'hD7][22:15];
        maskLastPipe_pipe_v_11 = _RANDOM[9'hD7][23];
        maskLastPipe_pipe_b_11 = _RANDOM[9'hD7][31:24];
        pipe_v_35 = _RANDOM[9'hD8][0];
        pipe_b_35 = _RANDOM[9'hD8][6:1];
        sinkVec_releasePipe_pipe_v_48 = _RANDOM[9'hD8][7];
        sinkVec_tokenCheck_counter_48 = _RANDOM[9'hD8][10:8];
        sinkVec_shifterReg_48_0_valid = _RANDOM[9'hD8][11];
        sinkVec_shifterReg_48_0_bits_vs = _RANDOM[9'hD8][16:12];
        sinkVec_shifterReg_48_0_bits_readSource = _RANDOM[9'hD8][18:17];
        sinkVec_shifterReg_48_0_bits_offset = _RANDOM[9'hD8][20:19];
        sinkVec_shifterReg_48_0_bits_instructionIndex = _RANDOM[9'hD8][23:21];
        sinkVec_releasePipe_pipe_v_49 = _RANDOM[9'hD8][24];
        sinkVec_tokenCheck_counter_49 = _RANDOM[9'hD8][27:25];
        sinkVec_shifterReg_49_0_valid = _RANDOM[9'hD8][28];
        sinkVec_shifterReg_49_0_bits_vs = {_RANDOM[9'hD8][31:29], _RANDOM[9'hD9][1:0]};
        sinkVec_shifterReg_49_0_bits_readSource = _RANDOM[9'hD9][3:2];
        sinkVec_shifterReg_49_0_bits_offset = _RANDOM[9'hD9][5:4];
        sinkVec_shifterReg_49_0_bits_instructionIndex = _RANDOM[9'hD9][8:6];
        maskUnitFirst_24 = _RANDOM[9'hD9][9];
        accessDataValid_pipe_v_24 = _RANDOM[9'hD9][10];
        accessDataValid_pipe_pipe_v_24 = _RANDOM[9'hD9][11];
        shifterReg_40_0_valid = _RANDOM[9'hD9][12];
        shifterReg_40_0_bits = {_RANDOM[9'hD9][31:13], _RANDOM[9'hDA][12:0]};
        accessDataValid_pipe_v_25 = _RANDOM[9'hDA][13];
        accessDataValid_pipe_pipe_v_25 = _RANDOM[9'hDA][14];
        shifterReg_41_0_valid = _RANDOM[9'hDA][15];
        shifterReg_41_0_bits = {_RANDOM[9'hDA][31:16], _RANDOM[9'hDB][15:0]};
        sinkVec_releasePipe_pipe_v_50 = _RANDOM[9'hDB][16];
        sinkVec_tokenCheck_counter_50 = _RANDOM[9'hDB][19:17];
        sinkVec_shifterReg_50_0_valid = _RANDOM[9'hDB][20];
        sinkVec_shifterReg_50_0_bits_vd = _RANDOM[9'hDB][25:21];
        sinkVec_shifterReg_50_0_bits_offset = _RANDOM[9'hDB][27:26];
        sinkVec_shifterReg_50_0_bits_mask = _RANDOM[9'hDB][31:28];
        sinkVec_shifterReg_50_0_bits_data = _RANDOM[9'hDC];
        sinkVec_shifterReg_50_0_bits_instructionIndex = _RANDOM[9'hDD][3:1];
        sinkVec_releasePipe_pipe_v_51 = _RANDOM[9'hDD][4];
        sinkVec_tokenCheck_counter_51 = _RANDOM[9'hDD][7:5];
        sinkVec_shifterReg_51_0_valid = _RANDOM[9'hDD][8];
        sinkVec_shifterReg_51_0_bits_vd = _RANDOM[9'hDD][13:9];
        sinkVec_shifterReg_51_0_bits_offset = _RANDOM[9'hDD][15:14];
        sinkVec_shifterReg_51_0_bits_mask = _RANDOM[9'hDD][19:16];
        sinkVec_shifterReg_51_0_bits_data = {_RANDOM[9'hDD][31:20], _RANDOM[9'hDE][19:0]};
        sinkVec_shifterReg_51_0_bits_last = _RANDOM[9'hDE][20];
        sinkVec_shifterReg_51_0_bits_instructionIndex = _RANDOM[9'hDE][23:21];
        maskUnitFirst_25 = _RANDOM[9'hDE][24];
        view__writeRelease_12_pipe_v = _RANDOM[9'hDE][25];
        pipe_v_36 = _RANDOM[9'hDE][26];
        instructionFinishedPipe_pipe_v_12 = _RANDOM[9'hDE][27];
        instructionFinishedPipe_pipe_b_12 = {_RANDOM[9'hDE][31:28], _RANDOM[9'hDF][3:0]};
        pipe_v_37 = _RANDOM[9'hDF][4];
        pipe_b_37 = {_RANDOM[9'hDF][31:5], _RANDOM[9'hE0][4:0]};
        pipe_pipe_v_12 = _RANDOM[9'hE0][5];
        pipe_pipe_b_12 = {_RANDOM[9'hE0][31:6], _RANDOM[9'hE1][5:0]};
        view__laneMaskSelect_12_pipe_v = _RANDOM[9'hE1][6];
        view__laneMaskSelect_12_pipe_b = _RANDOM[9'hE1][12:7];
        view__laneMaskSelect_12_pipe_pipe_v = _RANDOM[9'hE1][13];
        view__laneMaskSelect_12_pipe_pipe_b = _RANDOM[9'hE1][19:14];
        view__laneMaskSewSelect_12_pipe_v = _RANDOM[9'hE1][20];
        view__laneMaskSewSelect_12_pipe_b = _RANDOM[9'hE1][22:21];
        view__laneMaskSewSelect_12_pipe_pipe_v = _RANDOM[9'hE1][23];
        view__laneMaskSewSelect_12_pipe_pipe_b = _RANDOM[9'hE1][25:24];
        lsuLastPipe_pipe_v_12 = _RANDOM[9'hE1][26];
        lsuLastPipe_pipe_b_12 = {_RANDOM[9'hE1][31:27], _RANDOM[9'hE2][2:0]};
        maskLastPipe_pipe_v_12 = _RANDOM[9'hE2][3];
        maskLastPipe_pipe_b_12 = _RANDOM[9'hE2][11:4];
        pipe_v_38 = _RANDOM[9'hE2][12];
        pipe_b_38 = _RANDOM[9'hE2][18:13];
        sinkVec_releasePipe_pipe_v_52 = _RANDOM[9'hE2][19];
        sinkVec_tokenCheck_counter_52 = _RANDOM[9'hE2][22:20];
        sinkVec_shifterReg_52_0_valid = _RANDOM[9'hE2][23];
        sinkVec_shifterReg_52_0_bits_vs = _RANDOM[9'hE2][28:24];
        sinkVec_shifterReg_52_0_bits_readSource = _RANDOM[9'hE2][30:29];
        sinkVec_shifterReg_52_0_bits_offset = {_RANDOM[9'hE2][31], _RANDOM[9'hE3][0]};
        sinkVec_shifterReg_52_0_bits_instructionIndex = _RANDOM[9'hE3][3:1];
        sinkVec_releasePipe_pipe_v_53 = _RANDOM[9'hE3][4];
        sinkVec_tokenCheck_counter_53 = _RANDOM[9'hE3][7:5];
        sinkVec_shifterReg_53_0_valid = _RANDOM[9'hE3][8];
        sinkVec_shifterReg_53_0_bits_vs = _RANDOM[9'hE3][13:9];
        sinkVec_shifterReg_53_0_bits_readSource = _RANDOM[9'hE3][15:14];
        sinkVec_shifterReg_53_0_bits_offset = _RANDOM[9'hE3][17:16];
        sinkVec_shifterReg_53_0_bits_instructionIndex = _RANDOM[9'hE3][20:18];
        maskUnitFirst_26 = _RANDOM[9'hE3][21];
        accessDataValid_pipe_v_26 = _RANDOM[9'hE3][22];
        accessDataValid_pipe_pipe_v_26 = _RANDOM[9'hE3][23];
        shifterReg_42_0_valid = _RANDOM[9'hE3][24];
        shifterReg_42_0_bits = {_RANDOM[9'hE3][31:25], _RANDOM[9'hE4][24:0]};
        accessDataValid_pipe_v_27 = _RANDOM[9'hE4][25];
        accessDataValid_pipe_pipe_v_27 = _RANDOM[9'hE4][26];
        shifterReg_43_0_valid = _RANDOM[9'hE4][27];
        shifterReg_43_0_bits = {_RANDOM[9'hE4][31:28], _RANDOM[9'hE5][27:0]};
        sinkVec_releasePipe_pipe_v_54 = _RANDOM[9'hE5][28];
        sinkVec_tokenCheck_counter_54 = _RANDOM[9'hE5][31:29];
        sinkVec_shifterReg_54_0_valid = _RANDOM[9'hE6][0];
        sinkVec_shifterReg_54_0_bits_vd = _RANDOM[9'hE6][5:1];
        sinkVec_shifterReg_54_0_bits_offset = _RANDOM[9'hE6][7:6];
        sinkVec_shifterReg_54_0_bits_mask = _RANDOM[9'hE6][11:8];
        sinkVec_shifterReg_54_0_bits_data = {_RANDOM[9'hE6][31:12], _RANDOM[9'hE7][11:0]};
        sinkVec_shifterReg_54_0_bits_instructionIndex = _RANDOM[9'hE7][15:13];
        sinkVec_releasePipe_pipe_v_55 = _RANDOM[9'hE7][16];
        sinkVec_tokenCheck_counter_55 = _RANDOM[9'hE7][19:17];
        sinkVec_shifterReg_55_0_valid = _RANDOM[9'hE7][20];
        sinkVec_shifterReg_55_0_bits_vd = _RANDOM[9'hE7][25:21];
        sinkVec_shifterReg_55_0_bits_offset = _RANDOM[9'hE7][27:26];
        sinkVec_shifterReg_55_0_bits_mask = _RANDOM[9'hE7][31:28];
        sinkVec_shifterReg_55_0_bits_data = _RANDOM[9'hE8];
        sinkVec_shifterReg_55_0_bits_last = _RANDOM[9'hE9][0];
        sinkVec_shifterReg_55_0_bits_instructionIndex = _RANDOM[9'hE9][3:1];
        maskUnitFirst_27 = _RANDOM[9'hE9][4];
        view__writeRelease_13_pipe_v = _RANDOM[9'hE9][5];
        pipe_v_39 = _RANDOM[9'hE9][6];
        instructionFinishedPipe_pipe_v_13 = _RANDOM[9'hE9][7];
        instructionFinishedPipe_pipe_b_13 = _RANDOM[9'hE9][15:8];
        pipe_v_40 = _RANDOM[9'hE9][16];
        pipe_b_40 = {_RANDOM[9'hE9][31:17], _RANDOM[9'hEA][16:0]};
        pipe_pipe_v_13 = _RANDOM[9'hEA][17];
        pipe_pipe_b_13 = {_RANDOM[9'hEA][31:18], _RANDOM[9'hEB][17:0]};
        view__laneMaskSelect_13_pipe_v = _RANDOM[9'hEB][18];
        view__laneMaskSelect_13_pipe_b = _RANDOM[9'hEB][24:19];
        view__laneMaskSelect_13_pipe_pipe_v = _RANDOM[9'hEB][25];
        view__laneMaskSelect_13_pipe_pipe_b = _RANDOM[9'hEB][31:26];
        view__laneMaskSewSelect_13_pipe_v = _RANDOM[9'hEC][0];
        view__laneMaskSewSelect_13_pipe_b = _RANDOM[9'hEC][2:1];
        view__laneMaskSewSelect_13_pipe_pipe_v = _RANDOM[9'hEC][3];
        view__laneMaskSewSelect_13_pipe_pipe_b = _RANDOM[9'hEC][5:4];
        lsuLastPipe_pipe_v_13 = _RANDOM[9'hEC][6];
        lsuLastPipe_pipe_b_13 = _RANDOM[9'hEC][14:7];
        maskLastPipe_pipe_v_13 = _RANDOM[9'hEC][15];
        maskLastPipe_pipe_b_13 = _RANDOM[9'hEC][23:16];
        pipe_v_41 = _RANDOM[9'hEC][24];
        pipe_b_41 = _RANDOM[9'hEC][30:25];
        sinkVec_releasePipe_pipe_v_56 = _RANDOM[9'hEC][31];
        sinkVec_tokenCheck_counter_56 = _RANDOM[9'hED][2:0];
        sinkVec_shifterReg_56_0_valid = _RANDOM[9'hED][3];
        sinkVec_shifterReg_56_0_bits_vs = _RANDOM[9'hED][8:4];
        sinkVec_shifterReg_56_0_bits_readSource = _RANDOM[9'hED][10:9];
        sinkVec_shifterReg_56_0_bits_offset = _RANDOM[9'hED][12:11];
        sinkVec_shifterReg_56_0_bits_instructionIndex = _RANDOM[9'hED][15:13];
        sinkVec_releasePipe_pipe_v_57 = _RANDOM[9'hED][16];
        sinkVec_tokenCheck_counter_57 = _RANDOM[9'hED][19:17];
        sinkVec_shifterReg_57_0_valid = _RANDOM[9'hED][20];
        sinkVec_shifterReg_57_0_bits_vs = _RANDOM[9'hED][25:21];
        sinkVec_shifterReg_57_0_bits_readSource = _RANDOM[9'hED][27:26];
        sinkVec_shifterReg_57_0_bits_offset = _RANDOM[9'hED][29:28];
        sinkVec_shifterReg_57_0_bits_instructionIndex = {_RANDOM[9'hED][31:30], _RANDOM[9'hEE][0]};
        maskUnitFirst_28 = _RANDOM[9'hEE][1];
        accessDataValid_pipe_v_28 = _RANDOM[9'hEE][2];
        accessDataValid_pipe_pipe_v_28 = _RANDOM[9'hEE][3];
        shifterReg_44_0_valid = _RANDOM[9'hEE][4];
        shifterReg_44_0_bits = {_RANDOM[9'hEE][31:5], _RANDOM[9'hEF][4:0]};
        accessDataValid_pipe_v_29 = _RANDOM[9'hEF][5];
        accessDataValid_pipe_pipe_v_29 = _RANDOM[9'hEF][6];
        shifterReg_45_0_valid = _RANDOM[9'hEF][7];
        shifterReg_45_0_bits = {_RANDOM[9'hEF][31:8], _RANDOM[9'hF0][7:0]};
        sinkVec_releasePipe_pipe_v_58 = _RANDOM[9'hF0][8];
        sinkVec_tokenCheck_counter_58 = _RANDOM[9'hF0][11:9];
        sinkVec_shifterReg_58_0_valid = _RANDOM[9'hF0][12];
        sinkVec_shifterReg_58_0_bits_vd = _RANDOM[9'hF0][17:13];
        sinkVec_shifterReg_58_0_bits_offset = _RANDOM[9'hF0][19:18];
        sinkVec_shifterReg_58_0_bits_mask = _RANDOM[9'hF0][23:20];
        sinkVec_shifterReg_58_0_bits_data = {_RANDOM[9'hF0][31:24], _RANDOM[9'hF1][23:0]};
        sinkVec_shifterReg_58_0_bits_instructionIndex = _RANDOM[9'hF1][27:25];
        sinkVec_releasePipe_pipe_v_59 = _RANDOM[9'hF1][28];
        sinkVec_tokenCheck_counter_59 = _RANDOM[9'hF1][31:29];
        sinkVec_shifterReg_59_0_valid = _RANDOM[9'hF2][0];
        sinkVec_shifterReg_59_0_bits_vd = _RANDOM[9'hF2][5:1];
        sinkVec_shifterReg_59_0_bits_offset = _RANDOM[9'hF2][7:6];
        sinkVec_shifterReg_59_0_bits_mask = _RANDOM[9'hF2][11:8];
        sinkVec_shifterReg_59_0_bits_data = {_RANDOM[9'hF2][31:12], _RANDOM[9'hF3][11:0]};
        sinkVec_shifterReg_59_0_bits_last = _RANDOM[9'hF3][12];
        sinkVec_shifterReg_59_0_bits_instructionIndex = _RANDOM[9'hF3][15:13];
        maskUnitFirst_29 = _RANDOM[9'hF3][16];
        view__writeRelease_14_pipe_v = _RANDOM[9'hF3][17];
        pipe_v_42 = _RANDOM[9'hF3][18];
        instructionFinishedPipe_pipe_v_14 = _RANDOM[9'hF3][19];
        instructionFinishedPipe_pipe_b_14 = _RANDOM[9'hF3][27:20];
        pipe_v_43 = _RANDOM[9'hF3][28];
        pipe_b_43 = {_RANDOM[9'hF3][31:29], _RANDOM[9'hF4][28:0]};
        pipe_pipe_v_14 = _RANDOM[9'hF4][29];
        pipe_pipe_b_14 = {_RANDOM[9'hF4][31:30], _RANDOM[9'hF5][29:0]};
        view__laneMaskSelect_14_pipe_v = _RANDOM[9'hF5][30];
        view__laneMaskSelect_14_pipe_b = {_RANDOM[9'hF5][31], _RANDOM[9'hF6][4:0]};
        view__laneMaskSelect_14_pipe_pipe_v = _RANDOM[9'hF6][5];
        view__laneMaskSelect_14_pipe_pipe_b = _RANDOM[9'hF6][11:6];
        view__laneMaskSewSelect_14_pipe_v = _RANDOM[9'hF6][12];
        view__laneMaskSewSelect_14_pipe_b = _RANDOM[9'hF6][14:13];
        view__laneMaskSewSelect_14_pipe_pipe_v = _RANDOM[9'hF6][15];
        view__laneMaskSewSelect_14_pipe_pipe_b = _RANDOM[9'hF6][17:16];
        lsuLastPipe_pipe_v_14 = _RANDOM[9'hF6][18];
        lsuLastPipe_pipe_b_14 = _RANDOM[9'hF6][26:19];
        maskLastPipe_pipe_v_14 = _RANDOM[9'hF6][27];
        maskLastPipe_pipe_b_14 = {_RANDOM[9'hF6][31:28], _RANDOM[9'hF7][3:0]};
        pipe_v_44 = _RANDOM[9'hF7][4];
        pipe_b_44 = _RANDOM[9'hF7][10:5];
        sinkVec_releasePipe_pipe_v_60 = _RANDOM[9'hF7][11];
        sinkVec_tokenCheck_counter_60 = _RANDOM[9'hF7][14:12];
        sinkVec_shifterReg_60_0_valid = _RANDOM[9'hF7][15];
        sinkVec_shifterReg_60_0_bits_vs = _RANDOM[9'hF7][20:16];
        sinkVec_shifterReg_60_0_bits_readSource = _RANDOM[9'hF7][22:21];
        sinkVec_shifterReg_60_0_bits_offset = _RANDOM[9'hF7][24:23];
        sinkVec_shifterReg_60_0_bits_instructionIndex = _RANDOM[9'hF7][27:25];
        sinkVec_releasePipe_pipe_v_61 = _RANDOM[9'hF7][28];
        sinkVec_tokenCheck_counter_61 = _RANDOM[9'hF7][31:29];
        sinkVec_shifterReg_61_0_valid = _RANDOM[9'hF8][0];
        sinkVec_shifterReg_61_0_bits_vs = _RANDOM[9'hF8][5:1];
        sinkVec_shifterReg_61_0_bits_readSource = _RANDOM[9'hF8][7:6];
        sinkVec_shifterReg_61_0_bits_offset = _RANDOM[9'hF8][9:8];
        sinkVec_shifterReg_61_0_bits_instructionIndex = _RANDOM[9'hF8][12:10];
        maskUnitFirst_30 = _RANDOM[9'hF8][13];
        accessDataValid_pipe_v_30 = _RANDOM[9'hF8][14];
        accessDataValid_pipe_pipe_v_30 = _RANDOM[9'hF8][15];
        shifterReg_46_0_valid = _RANDOM[9'hF8][16];
        shifterReg_46_0_bits = {_RANDOM[9'hF8][31:17], _RANDOM[9'hF9][16:0]};
        accessDataValid_pipe_v_31 = _RANDOM[9'hF9][17];
        accessDataValid_pipe_pipe_v_31 = _RANDOM[9'hF9][18];
        shifterReg_47_0_valid = _RANDOM[9'hF9][19];
        shifterReg_47_0_bits = {_RANDOM[9'hF9][31:20], _RANDOM[9'hFA][19:0]};
        sinkVec_releasePipe_pipe_v_62 = _RANDOM[9'hFA][20];
        sinkVec_tokenCheck_counter_62 = _RANDOM[9'hFA][23:21];
        sinkVec_shifterReg_62_0_valid = _RANDOM[9'hFA][24];
        sinkVec_shifterReg_62_0_bits_vd = _RANDOM[9'hFA][29:25];
        sinkVec_shifterReg_62_0_bits_offset = _RANDOM[9'hFA][31:30];
        sinkVec_shifterReg_62_0_bits_mask = _RANDOM[9'hFB][3:0];
        sinkVec_shifterReg_62_0_bits_data = {_RANDOM[9'hFB][31:4], _RANDOM[9'hFC][3:0]};
        sinkVec_shifterReg_62_0_bits_instructionIndex = _RANDOM[9'hFC][7:5];
        sinkVec_releasePipe_pipe_v_63 = _RANDOM[9'hFC][8];
        sinkVec_tokenCheck_counter_63 = _RANDOM[9'hFC][11:9];
        sinkVec_shifterReg_63_0_valid = _RANDOM[9'hFC][12];
        sinkVec_shifterReg_63_0_bits_vd = _RANDOM[9'hFC][17:13];
        sinkVec_shifterReg_63_0_bits_offset = _RANDOM[9'hFC][19:18];
        sinkVec_shifterReg_63_0_bits_mask = _RANDOM[9'hFC][23:20];
        sinkVec_shifterReg_63_0_bits_data = {_RANDOM[9'hFC][31:24], _RANDOM[9'hFD][23:0]};
        sinkVec_shifterReg_63_0_bits_last = _RANDOM[9'hFD][24];
        sinkVec_shifterReg_63_0_bits_instructionIndex = _RANDOM[9'hFD][27:25];
        maskUnitFirst_31 = _RANDOM[9'hFD][28];
        view__writeRelease_15_pipe_v = _RANDOM[9'hFD][29];
        pipe_v_45 = _RANDOM[9'hFD][30];
        instructionFinishedPipe_pipe_v_15 = _RANDOM[9'hFD][31];
        instructionFinishedPipe_pipe_b_15 = _RANDOM[9'hFE][7:0];
        pipe_v_46 = _RANDOM[9'hFE][8];
        pipe_b_46 = {_RANDOM[9'hFE][31:9], _RANDOM[9'hFF][8:0]};
        pipe_pipe_v_15 = _RANDOM[9'hFF][9];
        pipe_pipe_b_15 = {_RANDOM[9'hFF][31:10], _RANDOM[9'h100][9:0]};
        view__laneMaskSelect_15_pipe_v = _RANDOM[9'h100][10];
        view__laneMaskSelect_15_pipe_b = _RANDOM[9'h100][16:11];
        view__laneMaskSelect_15_pipe_pipe_v = _RANDOM[9'h100][17];
        view__laneMaskSelect_15_pipe_pipe_b = _RANDOM[9'h100][23:18];
        view__laneMaskSewSelect_15_pipe_v = _RANDOM[9'h100][24];
        view__laneMaskSewSelect_15_pipe_b = _RANDOM[9'h100][26:25];
        view__laneMaskSewSelect_15_pipe_pipe_v = _RANDOM[9'h100][27];
        view__laneMaskSewSelect_15_pipe_pipe_b = _RANDOM[9'h100][29:28];
        lsuLastPipe_pipe_v_15 = _RANDOM[9'h100][30];
        lsuLastPipe_pipe_b_15 = {_RANDOM[9'h100][31], _RANDOM[9'h101][6:0]};
        maskLastPipe_pipe_v_15 = _RANDOM[9'h101][7];
        maskLastPipe_pipe_b_15 = _RANDOM[9'h101][15:8];
        pipe_v_47 = _RANDOM[9'h101][16];
        pipe_b_47 = _RANDOM[9'h101][22:17];
        pipe_v_48 = _RANDOM[9'h101][23];
        shifterReg_48_0_valid = _RANDOM[9'h101][24];
        shifterReg_48_0_bits_data = {_RANDOM[9'h101][31:25], _RANDOM[9'h102][24:0]};
        pipe_v_49 = _RANDOM[9'h102][25];
        shifterReg_49_0_valid = _RANDOM[9'h102][26];
        shifterReg_49_0_bits_data = {_RANDOM[9'h102][31:27], _RANDOM[9'h103][26:0]};
        shifterReg_49_0_bits_mask = _RANDOM[9'h103][28:27];
        shifterReg_49_0_bits_instructionIndex = _RANDOM[9'h103][31:29];
        shifterReg_49_0_bits_counter = _RANDOM[9'h104][5:0];
        pipe_v_50 = _RANDOM[9'h104][6];
        shifterReg_50_0_valid = _RANDOM[9'h104][7];
        shifterReg_50_0_bits_data = {_RANDOM[9'h104][31:8], _RANDOM[9'h105][7:0]};
        pipe_v_51 = _RANDOM[9'h105][8];
        shifterReg_51_0_valid = _RANDOM[9'h105][9];
        shifterReg_51_0_bits_data = {_RANDOM[9'h105][31:10], _RANDOM[9'h106][9:0]};
        shifterReg_51_0_bits_mask = _RANDOM[9'h106][11:10];
        shifterReg_51_0_bits_instructionIndex = _RANDOM[9'h106][14:12];
        shifterReg_51_0_bits_counter = _RANDOM[9'h106][20:15];
        pipe_v_52 = _RANDOM[9'h106][21];
        shifterReg_52_0_valid = _RANDOM[9'h106][22];
        shifterReg_52_0_bits_data = {_RANDOM[9'h106][31:23], _RANDOM[9'h107][22:0]};
        pipe_v_53 = _RANDOM[9'h107][23];
        shifterReg_53_0_valid = _RANDOM[9'h107][24];
        shifterReg_53_0_bits_data = {_RANDOM[9'h107][31:25], _RANDOM[9'h108][24:0]};
        shifterReg_53_0_bits_mask = _RANDOM[9'h108][26:25];
        shifterReg_53_0_bits_instructionIndex = _RANDOM[9'h108][29:27];
        shifterReg_53_0_bits_counter = {_RANDOM[9'h108][31:30], _RANDOM[9'h109][3:0]};
        pipe_v_54 = _RANDOM[9'h109][4];
        shifterReg_54_0_valid = _RANDOM[9'h109][5];
        shifterReg_54_0_bits_data = {_RANDOM[9'h109][31:6], _RANDOM[9'h10A][5:0]};
        pipe_v_55 = _RANDOM[9'h10A][6];
        shifterReg_55_0_valid = _RANDOM[9'h10A][7];
        shifterReg_55_0_bits_data = {_RANDOM[9'h10A][31:8], _RANDOM[9'h10B][7:0]};
        shifterReg_55_0_bits_mask = _RANDOM[9'h10B][9:8];
        shifterReg_55_0_bits_instructionIndex = _RANDOM[9'h10B][12:10];
        shifterReg_55_0_bits_counter = _RANDOM[9'h10B][18:13];
        pipe_v_56 = _RANDOM[9'h10B][19];
        shifterReg_56_0_valid = _RANDOM[9'h10B][20];
        shifterReg_56_0_bits_data = {_RANDOM[9'h10B][31:21], _RANDOM[9'h10C][20:0]};
        pipe_v_57 = _RANDOM[9'h10C][21];
        shifterReg_57_0_valid = _RANDOM[9'h10C][22];
        shifterReg_57_0_bits_data = {_RANDOM[9'h10C][31:23], _RANDOM[9'h10D][22:0]};
        shifterReg_57_0_bits_mask = _RANDOM[9'h10D][24:23];
        shifterReg_57_0_bits_instructionIndex = _RANDOM[9'h10D][27:25];
        shifterReg_57_0_bits_counter = {_RANDOM[9'h10D][31:28], _RANDOM[9'h10E][1:0]};
        pipe_v_58 = _RANDOM[9'h10E][2];
        shifterReg_58_0_valid = _RANDOM[9'h10E][3];
        shifterReg_58_0_bits_data = {_RANDOM[9'h10E][31:4], _RANDOM[9'h10F][3:0]};
        pipe_v_59 = _RANDOM[9'h10F][4];
        shifterReg_59_0_valid = _RANDOM[9'h10F][5];
        shifterReg_59_0_bits_data = {_RANDOM[9'h10F][31:6], _RANDOM[9'h110][5:0]};
        shifterReg_59_0_bits_mask = _RANDOM[9'h110][7:6];
        shifterReg_59_0_bits_instructionIndex = _RANDOM[9'h110][10:8];
        shifterReg_59_0_bits_counter = _RANDOM[9'h110][16:11];
        pipe_v_60 = _RANDOM[9'h110][17];
        shifterReg_60_0_valid = _RANDOM[9'h110][18];
        shifterReg_60_0_bits_data = {_RANDOM[9'h110][31:19], _RANDOM[9'h111][18:0]};
        pipe_v_61 = _RANDOM[9'h111][19];
        shifterReg_61_0_valid = _RANDOM[9'h111][20];
        shifterReg_61_0_bits_data = {_RANDOM[9'h111][31:21], _RANDOM[9'h112][20:0]};
        shifterReg_61_0_bits_mask = _RANDOM[9'h112][22:21];
        shifterReg_61_0_bits_instructionIndex = _RANDOM[9'h112][25:23];
        shifterReg_61_0_bits_counter = _RANDOM[9'h112][31:26];
        pipe_v_62 = _RANDOM[9'h113][0];
        shifterReg_62_0_valid = _RANDOM[9'h113][1];
        shifterReg_62_0_bits_data = {_RANDOM[9'h113][31:2], _RANDOM[9'h114][1:0]};
        pipe_v_63 = _RANDOM[9'h114][2];
        shifterReg_63_0_valid = _RANDOM[9'h114][3];
        shifterReg_63_0_bits_data = {_RANDOM[9'h114][31:4], _RANDOM[9'h115][3:0]};
        shifterReg_63_0_bits_mask = _RANDOM[9'h115][5:4];
        shifterReg_63_0_bits_instructionIndex = _RANDOM[9'h115][8:6];
        shifterReg_63_0_bits_counter = _RANDOM[9'h115][14:9];
        pipe_v_64 = _RANDOM[9'h115][15];
        shifterReg_64_0_valid = _RANDOM[9'h115][16];
        shifterReg_64_0_bits_data = {_RANDOM[9'h115][31:17], _RANDOM[9'h116][16:0]};
        pipe_v_65 = _RANDOM[9'h116][17];
        shifterReg_65_0_valid = _RANDOM[9'h116][18];
        shifterReg_65_0_bits_data = {_RANDOM[9'h116][31:19], _RANDOM[9'h117][18:0]};
        shifterReg_65_0_bits_mask = _RANDOM[9'h117][20:19];
        shifterReg_65_0_bits_instructionIndex = _RANDOM[9'h117][23:21];
        shifterReg_65_0_bits_counter = _RANDOM[9'h117][29:24];
        pipe_v_66 = _RANDOM[9'h117][30];
        shifterReg_66_0_valid = _RANDOM[9'h117][31];
        shifterReg_66_0_bits_data = _RANDOM[9'h118];
        pipe_v_67 = _RANDOM[9'h119][0];
        shifterReg_67_0_valid = _RANDOM[9'h119][1];
        shifterReg_67_0_bits_data = {_RANDOM[9'h119][31:2], _RANDOM[9'h11A][1:0]};
        shifterReg_67_0_bits_mask = _RANDOM[9'h11A][3:2];
        shifterReg_67_0_bits_instructionIndex = _RANDOM[9'h11A][6:4];
        shifterReg_67_0_bits_counter = _RANDOM[9'h11A][12:7];
        pipe_v_68 = _RANDOM[9'h11A][13];
        shifterReg_68_0_valid = _RANDOM[9'h11A][14];
        shifterReg_68_0_bits_data = {_RANDOM[9'h11A][31:15], _RANDOM[9'h11B][14:0]};
        pipe_v_69 = _RANDOM[9'h11B][15];
        shifterReg_69_0_valid = _RANDOM[9'h11B][16];
        shifterReg_69_0_bits_data = {_RANDOM[9'h11B][31:17], _RANDOM[9'h11C][16:0]};
        shifterReg_69_0_bits_mask = _RANDOM[9'h11C][18:17];
        shifterReg_69_0_bits_instructionIndex = _RANDOM[9'h11C][21:19];
        shifterReg_69_0_bits_counter = _RANDOM[9'h11C][27:22];
        pipe_v_70 = _RANDOM[9'h11C][28];
        shifterReg_70_0_valid = _RANDOM[9'h11C][29];
        shifterReg_70_0_bits_data = {_RANDOM[9'h11C][31:30], _RANDOM[9'h11D][29:0]};
        pipe_v_71 = _RANDOM[9'h11D][30];
        shifterReg_71_0_valid = _RANDOM[9'h11D][31];
        shifterReg_71_0_bits_data = _RANDOM[9'h11E];
        shifterReg_71_0_bits_mask = _RANDOM[9'h11F][1:0];
        shifterReg_71_0_bits_instructionIndex = _RANDOM[9'h11F][4:2];
        shifterReg_71_0_bits_counter = _RANDOM[9'h11F][10:5];
        pipe_v_72 = _RANDOM[9'h11F][11];
        shifterReg_72_0_valid = _RANDOM[9'h11F][12];
        shifterReg_72_0_bits_data = {_RANDOM[9'h11F][31:13], _RANDOM[9'h120][12:0]};
        pipe_v_73 = _RANDOM[9'h120][13];
        shifterReg_73_0_valid = _RANDOM[9'h120][14];
        shifterReg_73_0_bits_data = {_RANDOM[9'h120][31:15], _RANDOM[9'h121][14:0]};
        shifterReg_73_0_bits_mask = _RANDOM[9'h121][16:15];
        shifterReg_73_0_bits_instructionIndex = _RANDOM[9'h121][19:17];
        shifterReg_73_0_bits_counter = _RANDOM[9'h121][25:20];
        pipe_v_74 = _RANDOM[9'h121][26];
        shifterReg_74_0_valid = _RANDOM[9'h121][27];
        shifterReg_74_0_bits_data = {_RANDOM[9'h121][31:28], _RANDOM[9'h122][27:0]};
        pipe_v_75 = _RANDOM[9'h122][28];
        shifterReg_75_0_valid = _RANDOM[9'h122][29];
        shifterReg_75_0_bits_data = {_RANDOM[9'h122][31:30], _RANDOM[9'h123][29:0]};
        shifterReg_75_0_bits_mask = _RANDOM[9'h123][31:30];
        shifterReg_75_0_bits_instructionIndex = _RANDOM[9'h124][2:0];
        shifterReg_75_0_bits_counter = _RANDOM[9'h124][8:3];
        pipe_v_76 = _RANDOM[9'h124][9];
        shifterReg_76_0_valid = _RANDOM[9'h124][10];
        shifterReg_76_0_bits_data = {_RANDOM[9'h124][31:11], _RANDOM[9'h125][10:0]};
        pipe_v_77 = _RANDOM[9'h125][11];
        shifterReg_77_0_valid = _RANDOM[9'h125][12];
        shifterReg_77_0_bits_data = {_RANDOM[9'h125][31:13], _RANDOM[9'h126][12:0]};
        shifterReg_77_0_bits_mask = _RANDOM[9'h126][14:13];
        shifterReg_77_0_bits_instructionIndex = _RANDOM[9'h126][17:15];
        shifterReg_77_0_bits_counter = _RANDOM[9'h126][23:18];
        pipe_v_78 = _RANDOM[9'h126][24];
        shifterReg_78_0_valid = _RANDOM[9'h126][25];
        shifterReg_78_0_bits_data = {_RANDOM[9'h126][31:26], _RANDOM[9'h127][25:0]};
        pipe_v_79 = _RANDOM[9'h127][26];
        shifterReg_79_0_valid = _RANDOM[9'h127][27];
        shifterReg_79_0_bits_data = {_RANDOM[9'h127][31:28], _RANDOM[9'h128][27:0]};
        shifterReg_79_0_bits_mask = _RANDOM[9'h128][29:28];
        shifterReg_79_0_bits_instructionIndex = {_RANDOM[9'h128][31:30], _RANDOM[9'h129][0]};
        shifterReg_79_0_bits_counter = _RANDOM[9'h129][6:1];
        pipe_v_80 = _RANDOM[9'h129][7];
        shifterReg_80_0_valid = _RANDOM[9'h129][8];
        shifterReg_80_0_bits_data = {_RANDOM[9'h129][31:9], _RANDOM[9'h12A][8:0]};
        pipe_v_81 = _RANDOM[9'h12A][9];
        shifterReg_81_0_valid = _RANDOM[9'h12A][10];
        shifterReg_81_0_bits_data = {_RANDOM[9'h12A][31:11], _RANDOM[9'h12B][10:0]};
        shifterReg_81_0_bits_mask = _RANDOM[9'h12B][12:11];
        shifterReg_81_0_bits_instructionIndex = _RANDOM[9'h12B][15:13];
        shifterReg_81_0_bits_counter = _RANDOM[9'h12B][21:16];
        pipe_v_82 = _RANDOM[9'h12B][22];
        shifterReg_82_0_valid = _RANDOM[9'h12B][23];
        shifterReg_82_0_bits_data = {_RANDOM[9'h12B][31:24], _RANDOM[9'h12C][23:0]};
        pipe_v_83 = _RANDOM[9'h12C][24];
        shifterReg_83_0_valid = _RANDOM[9'h12C][25];
        shifterReg_83_0_bits_data = {_RANDOM[9'h12C][31:26], _RANDOM[9'h12D][25:0]};
        shifterReg_83_0_bits_mask = _RANDOM[9'h12D][27:26];
        shifterReg_83_0_bits_instructionIndex = _RANDOM[9'h12D][30:28];
        shifterReg_83_0_bits_counter = {_RANDOM[9'h12D][31], _RANDOM[9'h12E][4:0]};
        pipe_v_84 = _RANDOM[9'h12E][5];
        shifterReg_84_0_valid = _RANDOM[9'h12E][6];
        shifterReg_84_0_bits_data = {_RANDOM[9'h12E][31:7], _RANDOM[9'h12F][6:0]};
        pipe_v_85 = _RANDOM[9'h12F][7];
        shifterReg_85_0_valid = _RANDOM[9'h12F][8];
        shifterReg_85_0_bits_data = {_RANDOM[9'h12F][31:9], _RANDOM[9'h130][8:0]};
        shifterReg_85_0_bits_mask = _RANDOM[9'h130][10:9];
        shifterReg_85_0_bits_instructionIndex = _RANDOM[9'h130][13:11];
        shifterReg_85_0_bits_counter = _RANDOM[9'h130][19:14];
        pipe_v_86 = _RANDOM[9'h130][20];
        shifterReg_86_0_valid = _RANDOM[9'h130][21];
        shifterReg_86_0_bits_data = {_RANDOM[9'h130][31:22], _RANDOM[9'h131][21:0]};
        pipe_v_87 = _RANDOM[9'h131][22];
        shifterReg_87_0_valid = _RANDOM[9'h131][23];
        shifterReg_87_0_bits_data = {_RANDOM[9'h131][31:24], _RANDOM[9'h132][23:0]};
        shifterReg_87_0_bits_mask = _RANDOM[9'h132][25:24];
        shifterReg_87_0_bits_instructionIndex = _RANDOM[9'h132][28:26];
        shifterReg_87_0_bits_counter = {_RANDOM[9'h132][31:29], _RANDOM[9'h133][2:0]};
        pipe_v_88 = _RANDOM[9'h133][3];
        shifterReg_88_0_valid = _RANDOM[9'h133][4];
        shifterReg_88_0_bits_data = {_RANDOM[9'h133][31:5], _RANDOM[9'h134][4:0]};
        pipe_v_89 = _RANDOM[9'h134][5];
        shifterReg_89_0_valid = _RANDOM[9'h134][6];
        shifterReg_89_0_bits_data = {_RANDOM[9'h134][31:7], _RANDOM[9'h135][6:0]};
        shifterReg_89_0_bits_mask = _RANDOM[9'h135][8:7];
        shifterReg_89_0_bits_instructionIndex = _RANDOM[9'h135][11:9];
        shifterReg_89_0_bits_counter = _RANDOM[9'h135][17:12];
        pipe_v_90 = _RANDOM[9'h135][18];
        shifterReg_90_0_valid = _RANDOM[9'h135][19];
        shifterReg_90_0_bits_data = {_RANDOM[9'h135][31:20], _RANDOM[9'h136][19:0]};
        pipe_v_91 = _RANDOM[9'h136][20];
        shifterReg_91_0_valid = _RANDOM[9'h136][21];
        shifterReg_91_0_bits_data = {_RANDOM[9'h136][31:22], _RANDOM[9'h137][21:0]};
        shifterReg_91_0_bits_mask = _RANDOM[9'h137][23:22];
        shifterReg_91_0_bits_instructionIndex = _RANDOM[9'h137][26:24];
        shifterReg_91_0_bits_counter = {_RANDOM[9'h137][31:27], _RANDOM[9'h138][0]};
        pipe_v_92 = _RANDOM[9'h138][1];
        shifterReg_92_0_valid = _RANDOM[9'h138][2];
        shifterReg_92_0_bits_data = {_RANDOM[9'h138][31:3], _RANDOM[9'h139][2:0]};
        pipe_v_93 = _RANDOM[9'h139][3];
        shifterReg_93_0_valid = _RANDOM[9'h139][4];
        shifterReg_93_0_bits_data = {_RANDOM[9'h139][31:5], _RANDOM[9'h13A][4:0]};
        shifterReg_93_0_bits_mask = _RANDOM[9'h13A][6:5];
        shifterReg_93_0_bits_instructionIndex = _RANDOM[9'h13A][9:7];
        shifterReg_93_0_bits_counter = _RANDOM[9'h13A][15:10];
        pipe_v_94 = _RANDOM[9'h13A][16];
        shifterReg_94_0_valid = _RANDOM[9'h13A][17];
        shifterReg_94_0_bits_data = {_RANDOM[9'h13A][31:18], _RANDOM[9'h13B][17:0]};
        pipe_v_95 = _RANDOM[9'h13B][18];
        shifterReg_95_0_valid = _RANDOM[9'h13B][19];
        shifterReg_95_0_bits_data = {_RANDOM[9'h13B][31:20], _RANDOM[9'h13C][19:0]};
        shifterReg_95_0_bits_mask = _RANDOM[9'h13C][21:20];
        shifterReg_95_0_bits_instructionIndex = _RANDOM[9'h13C][24:22];
        shifterReg_95_0_bits_counter = _RANDOM[9'h13C][30:25];
        pipe_v_96 = _RANDOM[9'h13C][31];
        shifterReg_96_0_valid = _RANDOM[9'h13D][0];
        shifterReg_96_0_bits_data = {_RANDOM[9'h13D][31:1], _RANDOM[9'h13E][0]};
        pipe_v_97 = _RANDOM[9'h13E][1];
        shifterReg_97_0_valid = _RANDOM[9'h13E][2];
        shifterReg_97_0_bits_data = {_RANDOM[9'h13E][31:3], _RANDOM[9'h13F][2:0]};
        shifterReg_97_0_bits_mask = _RANDOM[9'h13F][4:3];
        shifterReg_97_0_bits_instructionIndex = _RANDOM[9'h13F][7:5];
        shifterReg_97_0_bits_counter = _RANDOM[9'h13F][13:8];
        pipe_v_98 = _RANDOM[9'h13F][14];
        shifterReg_98_0_valid = _RANDOM[9'h13F][15];
        shifterReg_98_0_bits_data = {_RANDOM[9'h13F][31:16], _RANDOM[9'h140][15:0]};
        pipe_v_99 = _RANDOM[9'h140][16];
        shifterReg_99_0_valid = _RANDOM[9'h140][17];
        shifterReg_99_0_bits_data = {_RANDOM[9'h140][31:18], _RANDOM[9'h141][17:0]};
        shifterReg_99_0_bits_mask = _RANDOM[9'h141][19:18];
        shifterReg_99_0_bits_instructionIndex = _RANDOM[9'h141][22:20];
        shifterReg_99_0_bits_counter = _RANDOM[9'h141][28:23];
        pipe_v_100 = _RANDOM[9'h141][29];
        shifterReg_100_0_valid = _RANDOM[9'h141][30];
        shifterReg_100_0_bits_data = {_RANDOM[9'h141][31], _RANDOM[9'h142][30:0]};
        pipe_v_101 = _RANDOM[9'h142][31];
        shifterReg_101_0_valid = _RANDOM[9'h143][0];
        shifterReg_101_0_bits_data = {_RANDOM[9'h143][31:1], _RANDOM[9'h144][0]};
        shifterReg_101_0_bits_mask = _RANDOM[9'h144][2:1];
        shifterReg_101_0_bits_instructionIndex = _RANDOM[9'h144][5:3];
        shifterReg_101_0_bits_counter = _RANDOM[9'h144][11:6];
        pipe_v_102 = _RANDOM[9'h144][12];
        shifterReg_102_0_valid = _RANDOM[9'h144][13];
        shifterReg_102_0_bits_data = {_RANDOM[9'h144][31:14], _RANDOM[9'h145][13:0]};
        pipe_v_103 = _RANDOM[9'h145][14];
        shifterReg_103_0_valid = _RANDOM[9'h145][15];
        shifterReg_103_0_bits_data = {_RANDOM[9'h145][31:16], _RANDOM[9'h146][15:0]};
        shifterReg_103_0_bits_mask = _RANDOM[9'h146][17:16];
        shifterReg_103_0_bits_instructionIndex = _RANDOM[9'h146][20:18];
        shifterReg_103_0_bits_counter = _RANDOM[9'h146][26:21];
        pipe_v_104 = _RANDOM[9'h146][27];
        shifterReg_104_0_valid = _RANDOM[9'h146][28];
        shifterReg_104_0_bits_data = {_RANDOM[9'h146][31:29], _RANDOM[9'h147][28:0]};
        pipe_v_105 = _RANDOM[9'h147][29];
        shifterReg_105_0_valid = _RANDOM[9'h147][30];
        shifterReg_105_0_bits_data = {_RANDOM[9'h147][31], _RANDOM[9'h148][30:0]};
        shifterReg_105_0_bits_mask = {_RANDOM[9'h148][31], _RANDOM[9'h149][0]};
        shifterReg_105_0_bits_instructionIndex = _RANDOM[9'h149][3:1];
        shifterReg_105_0_bits_counter = _RANDOM[9'h149][9:4];
        pipe_v_106 = _RANDOM[9'h149][10];
        shifterReg_106_0_valid = _RANDOM[9'h149][11];
        shifterReg_106_0_bits_data = {_RANDOM[9'h149][31:12], _RANDOM[9'h14A][11:0]};
        pipe_v_107 = _RANDOM[9'h14A][12];
        shifterReg_107_0_valid = _RANDOM[9'h14A][13];
        shifterReg_107_0_bits_data = {_RANDOM[9'h14A][31:14], _RANDOM[9'h14B][13:0]};
        shifterReg_107_0_bits_mask = _RANDOM[9'h14B][15:14];
        shifterReg_107_0_bits_instructionIndex = _RANDOM[9'h14B][18:16];
        shifterReg_107_0_bits_counter = _RANDOM[9'h14B][24:19];
        pipe_v_108 = _RANDOM[9'h14B][25];
        shifterReg_108_0_valid = _RANDOM[9'h14B][26];
        shifterReg_108_0_bits_data = {_RANDOM[9'h14B][31:27], _RANDOM[9'h14C][26:0]};
        pipe_v_109 = _RANDOM[9'h14C][27];
        shifterReg_109_0_valid = _RANDOM[9'h14C][28];
        shifterReg_109_0_bits_data = {_RANDOM[9'h14C][31:29], _RANDOM[9'h14D][28:0]};
        shifterReg_109_0_bits_mask = _RANDOM[9'h14D][30:29];
        shifterReg_109_0_bits_instructionIndex = {_RANDOM[9'h14D][31], _RANDOM[9'h14E][1:0]};
        shifterReg_109_0_bits_counter = _RANDOM[9'h14E][7:2];
        pipe_v_110 = _RANDOM[9'h14E][8];
        shifterReg_110_0_valid = _RANDOM[9'h14E][9];
        shifterReg_110_0_bits_data = {_RANDOM[9'h14E][31:10], _RANDOM[9'h14F][9:0]};
        pipe_v_111 = _RANDOM[9'h14F][10];
        shifterReg_111_0_valid = _RANDOM[9'h14F][11];
        shifterReg_111_0_bits_data = {_RANDOM[9'h14F][31:12], _RANDOM[9'h150][11:0]};
        shifterReg_111_0_bits_mask = _RANDOM[9'h150][13:12];
        shifterReg_111_0_bits_instructionIndex = _RANDOM[9'h150][16:14];
        shifterReg_111_0_bits_counter = _RANDOM[9'h150][22:17];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign x22_1_valid = _lsu_vrfWritePort_0_valid;
  assign x22_1_bits_vd = _lsu_vrfWritePort_0_bits_vd;
  assign x22_1_bits_mask = _lsu_vrfWritePort_0_bits_mask;
  assign x22_1_bits_instructionIndex = _lsu_vrfWritePort_0_bits_instructionIndex;
  assign x22_1_1_valid = _lsu_vrfWritePort_1_valid;
  assign x22_1_1_bits_vd = _lsu_vrfWritePort_1_bits_vd;
  assign x22_1_1_bits_mask = _lsu_vrfWritePort_1_bits_mask;
  assign x22_1_1_bits_instructionIndex = _lsu_vrfWritePort_1_bits_instructionIndex;
  assign x22_2_1_valid = _lsu_vrfWritePort_2_valid;
  assign x22_2_1_bits_vd = _lsu_vrfWritePort_2_bits_vd;
  assign x22_2_1_bits_mask = _lsu_vrfWritePort_2_bits_mask;
  assign x22_2_1_bits_instructionIndex = _lsu_vrfWritePort_2_bits_instructionIndex;
  assign x22_3_1_valid = _lsu_vrfWritePort_3_valid;
  assign x22_3_1_bits_vd = _lsu_vrfWritePort_3_bits_vd;
  assign x22_3_1_bits_mask = _lsu_vrfWritePort_3_bits_mask;
  assign x22_3_1_bits_instructionIndex = _lsu_vrfWritePort_3_bits_instructionIndex;
  assign x22_4_1_valid = _lsu_vrfWritePort_4_valid;
  assign x22_4_1_bits_vd = _lsu_vrfWritePort_4_bits_vd;
  assign x22_4_1_bits_mask = _lsu_vrfWritePort_4_bits_mask;
  assign x22_4_1_bits_instructionIndex = _lsu_vrfWritePort_4_bits_instructionIndex;
  assign x22_5_1_valid = _lsu_vrfWritePort_5_valid;
  assign x22_5_1_bits_vd = _lsu_vrfWritePort_5_bits_vd;
  assign x22_5_1_bits_mask = _lsu_vrfWritePort_5_bits_mask;
  assign x22_5_1_bits_instructionIndex = _lsu_vrfWritePort_5_bits_instructionIndex;
  assign x22_6_1_valid = _lsu_vrfWritePort_6_valid;
  assign x22_6_1_bits_vd = _lsu_vrfWritePort_6_bits_vd;
  assign x22_6_1_bits_mask = _lsu_vrfWritePort_6_bits_mask;
  assign x22_6_1_bits_instructionIndex = _lsu_vrfWritePort_6_bits_instructionIndex;
  assign x22_7_1_valid = _lsu_vrfWritePort_7_valid;
  assign x22_7_1_bits_vd = _lsu_vrfWritePort_7_bits_vd;
  assign x22_7_1_bits_mask = _lsu_vrfWritePort_7_bits_mask;
  assign x22_7_1_bits_instructionIndex = _lsu_vrfWritePort_7_bits_instructionIndex;
  assign x22_8_1_valid = _lsu_vrfWritePort_8_valid;
  assign x22_8_1_bits_vd = _lsu_vrfWritePort_8_bits_vd;
  assign x22_8_1_bits_mask = _lsu_vrfWritePort_8_bits_mask;
  assign x22_8_1_bits_instructionIndex = _lsu_vrfWritePort_8_bits_instructionIndex;
  assign x22_9_1_valid = _lsu_vrfWritePort_9_valid;
  assign x22_9_1_bits_vd = _lsu_vrfWritePort_9_bits_vd;
  assign x22_9_1_bits_mask = _lsu_vrfWritePort_9_bits_mask;
  assign x22_9_1_bits_instructionIndex = _lsu_vrfWritePort_9_bits_instructionIndex;
  assign x22_10_1_valid = _lsu_vrfWritePort_10_valid;
  assign x22_10_1_bits_vd = _lsu_vrfWritePort_10_bits_vd;
  assign x22_10_1_bits_mask = _lsu_vrfWritePort_10_bits_mask;
  assign x22_10_1_bits_instructionIndex = _lsu_vrfWritePort_10_bits_instructionIndex;
  assign x22_11_1_valid = _lsu_vrfWritePort_11_valid;
  assign x22_11_1_bits_vd = _lsu_vrfWritePort_11_bits_vd;
  assign x22_11_1_bits_mask = _lsu_vrfWritePort_11_bits_mask;
  assign x22_11_1_bits_instructionIndex = _lsu_vrfWritePort_11_bits_instructionIndex;
  assign x22_12_1_valid = _lsu_vrfWritePort_12_valid;
  assign x22_12_1_bits_vd = _lsu_vrfWritePort_12_bits_vd;
  assign x22_12_1_bits_mask = _lsu_vrfWritePort_12_bits_mask;
  assign x22_12_1_bits_instructionIndex = _lsu_vrfWritePort_12_bits_instructionIndex;
  assign x22_13_1_valid = _lsu_vrfWritePort_13_valid;
  assign x22_13_1_bits_vd = _lsu_vrfWritePort_13_bits_vd;
  assign x22_13_1_bits_mask = _lsu_vrfWritePort_13_bits_mask;
  assign x22_13_1_bits_instructionIndex = _lsu_vrfWritePort_13_bits_instructionIndex;
  assign x22_14_1_valid = _lsu_vrfWritePort_14_valid;
  assign x22_14_1_bits_vd = _lsu_vrfWritePort_14_bits_vd;
  assign x22_14_1_bits_mask = _lsu_vrfWritePort_14_bits_mask;
  assign x22_14_1_bits_instructionIndex = _lsu_vrfWritePort_14_bits_instructionIndex;
  assign x22_15_1_valid = _lsu_vrfWritePort_15_valid;
  assign x22_15_1_bits_vd = _lsu_vrfWritePort_15_bits_vd;
  assign x22_15_1_bits_mask = _lsu_vrfWritePort_15_bits_mask;
  assign x22_15_1_bits_instructionIndex = _lsu_vrfWritePort_15_bits_instructionIndex;
  assign x22_0_valid = _maskUnit_exeResp_0_valid;
  assign x22_0_bits_mask = _maskUnit_exeResp_0_bits_mask;
  assign x22_0_bits_instructionIndex = _maskUnit_exeResp_0_bits_instructionIndex;
  assign x22_1_0_valid = _maskUnit_exeResp_1_valid;
  assign x22_1_0_bits_mask = _maskUnit_exeResp_1_bits_mask;
  assign x22_1_0_bits_instructionIndex = _maskUnit_exeResp_1_bits_instructionIndex;
  assign x22_2_0_valid = _maskUnit_exeResp_2_valid;
  assign x22_2_0_bits_mask = _maskUnit_exeResp_2_bits_mask;
  assign x22_2_0_bits_instructionIndex = _maskUnit_exeResp_2_bits_instructionIndex;
  assign x22_3_0_valid = _maskUnit_exeResp_3_valid;
  assign x22_3_0_bits_mask = _maskUnit_exeResp_3_bits_mask;
  assign x22_3_0_bits_instructionIndex = _maskUnit_exeResp_3_bits_instructionIndex;
  assign x22_4_0_valid = _maskUnit_exeResp_4_valid;
  assign x22_4_0_bits_mask = _maskUnit_exeResp_4_bits_mask;
  assign x22_4_0_bits_instructionIndex = _maskUnit_exeResp_4_bits_instructionIndex;
  assign x22_5_0_valid = _maskUnit_exeResp_5_valid;
  assign x22_5_0_bits_mask = _maskUnit_exeResp_5_bits_mask;
  assign x22_5_0_bits_instructionIndex = _maskUnit_exeResp_5_bits_instructionIndex;
  assign x22_6_0_valid = _maskUnit_exeResp_6_valid;
  assign x22_6_0_bits_mask = _maskUnit_exeResp_6_bits_mask;
  assign x22_6_0_bits_instructionIndex = _maskUnit_exeResp_6_bits_instructionIndex;
  assign x22_7_0_valid = _maskUnit_exeResp_7_valid;
  assign x22_7_0_bits_mask = _maskUnit_exeResp_7_bits_mask;
  assign x22_7_0_bits_instructionIndex = _maskUnit_exeResp_7_bits_instructionIndex;
  assign x22_8_0_valid = _maskUnit_exeResp_8_valid;
  assign x22_8_0_bits_mask = _maskUnit_exeResp_8_bits_mask;
  assign x22_8_0_bits_instructionIndex = _maskUnit_exeResp_8_bits_instructionIndex;
  assign x22_9_0_valid = _maskUnit_exeResp_9_valid;
  assign x22_9_0_bits_mask = _maskUnit_exeResp_9_bits_mask;
  assign x22_9_0_bits_instructionIndex = _maskUnit_exeResp_9_bits_instructionIndex;
  assign x22_10_0_valid = _maskUnit_exeResp_10_valid;
  assign x22_10_0_bits_mask = _maskUnit_exeResp_10_bits_mask;
  assign x22_10_0_bits_instructionIndex = _maskUnit_exeResp_10_bits_instructionIndex;
  assign x22_11_0_valid = _maskUnit_exeResp_11_valid;
  assign x22_11_0_bits_mask = _maskUnit_exeResp_11_bits_mask;
  assign x22_11_0_bits_instructionIndex = _maskUnit_exeResp_11_bits_instructionIndex;
  assign x22_12_0_valid = _maskUnit_exeResp_12_valid;
  assign x22_12_0_bits_mask = _maskUnit_exeResp_12_bits_mask;
  assign x22_12_0_bits_instructionIndex = _maskUnit_exeResp_12_bits_instructionIndex;
  assign x22_13_0_valid = _maskUnit_exeResp_13_valid;
  assign x22_13_0_bits_mask = _maskUnit_exeResp_13_bits_mask;
  assign x22_13_0_bits_instructionIndex = _maskUnit_exeResp_13_bits_instructionIndex;
  assign x22_14_0_valid = _maskUnit_exeResp_14_valid;
  assign x22_14_0_bits_mask = _maskUnit_exeResp_14_bits_mask;
  assign x22_14_0_bits_instructionIndex = _maskUnit_exeResp_14_bits_instructionIndex;
  assign x22_15_0_valid = _maskUnit_exeResp_15_valid;
  assign x22_15_0_bits_mask = _maskUnit_exeResp_15_bits_mask;
  assign x22_15_0_bits_instructionIndex = _maskUnit_exeResp_15_bits_instructionIndex;
  wire         queue_empty;
  assign queue_empty = _queue_fifo_empty;
  wire         queue_full;
  assign queue_full = _queue_fifo_full;
  wire         queue_1_empty;
  assign queue_1_empty = _queue_fifo_1_empty;
  wire         queue_1_full;
  assign queue_1_full = _queue_fifo_1_full;
  wire         queue_2_empty;
  assign queue_2_empty = _queue_fifo_2_empty;
  wire         queue_2_full;
  assign queue_2_full = _queue_fifo_2_full;
  wire         queue_3_empty;
  assign queue_3_empty = _queue_fifo_3_empty;
  wire         queue_3_full;
  assign queue_3_full = _queue_fifo_3_full;
  wire         queue_4_empty;
  assign queue_4_empty = _queue_fifo_4_empty;
  wire         queue_4_full;
  assign queue_4_full = _queue_fifo_4_full;
  wire         queue_5_empty;
  assign queue_5_empty = _queue_fifo_5_empty;
  wire         queue_5_full;
  assign queue_5_full = _queue_fifo_5_full;
  wire         queue_6_empty;
  assign queue_6_empty = _queue_fifo_6_empty;
  wire         queue_6_full;
  assign queue_6_full = _queue_fifo_6_full;
  wire         queue_7_empty;
  assign queue_7_empty = _queue_fifo_7_empty;
  wire         queue_7_full;
  assign queue_7_full = _queue_fifo_7_full;
  wire         queue_8_empty;
  assign queue_8_empty = _queue_fifo_8_empty;
  wire         queue_8_full;
  assign queue_8_full = _queue_fifo_8_full;
  wire         queue_9_empty;
  assign queue_9_empty = _queue_fifo_9_empty;
  wire         queue_9_full;
  assign queue_9_full = _queue_fifo_9_full;
  wire         queue_10_empty;
  assign queue_10_empty = _queue_fifo_10_empty;
  wire         queue_10_full;
  assign queue_10_full = _queue_fifo_10_full;
  wire         queue_11_empty;
  assign queue_11_empty = _queue_fifo_11_empty;
  wire         queue_11_full;
  assign queue_11_full = _queue_fifo_11_full;
  wire         queue_12_empty;
  assign queue_12_empty = _queue_fifo_12_empty;
  wire         queue_12_full;
  assign queue_12_full = _queue_fifo_12_full;
  wire         queue_13_empty;
  assign queue_13_empty = _queue_fifo_13_empty;
  wire         queue_13_full;
  assign queue_13_full = _queue_fifo_13_full;
  wire         queue_14_empty;
  assign queue_14_empty = _queue_fifo_14_empty;
  wire         queue_14_full;
  assign queue_14_full = _queue_fifo_14_full;
  wire         queue_15_empty;
  assign queue_15_empty = _queue_fifo_15_empty;
  wire         queue_15_full;
  assign queue_15_full = _queue_fifo_15_full;
  assign accessDataSource_bits = _laneVec_0_vrfReadDataChannel;
  assign accessDataSource_1_bits = _laneVec_0_vrfReadDataChannel;
  wire         sinkVec_queue_empty;
  assign sinkVec_queue_empty = _sinkVec_queue_fifo_empty;
  wire         sinkVec_queue_full;
  assign sinkVec_queue_full = _sinkVec_queue_fifo_full;
  wire         sinkVec_queue_1_empty;
  assign sinkVec_queue_1_empty = _sinkVec_queue_fifo_1_empty;
  wire         sinkVec_queue_1_full;
  assign sinkVec_queue_1_full = _sinkVec_queue_fifo_1_full;
  wire         sinkVec_queue_2_empty;
  assign sinkVec_queue_2_empty = _sinkVec_queue_fifo_2_empty;
  wire         sinkVec_queue_2_full;
  assign sinkVec_queue_2_full = _sinkVec_queue_fifo_2_full;
  wire         sinkVec_queue_3_empty;
  assign sinkVec_queue_3_empty = _sinkVec_queue_fifo_3_empty;
  wire         sinkVec_queue_3_full;
  assign sinkVec_queue_3_full = _sinkVec_queue_fifo_3_full;
  assign accessDataSource_2_bits = _laneVec_1_vrfReadDataChannel;
  assign accessDataSource_3_bits = _laneVec_1_vrfReadDataChannel;
  wire         sinkVec_queue_4_empty;
  assign sinkVec_queue_4_empty = _sinkVec_queue_fifo_4_empty;
  wire         sinkVec_queue_4_full;
  assign sinkVec_queue_4_full = _sinkVec_queue_fifo_4_full;
  wire         sinkVec_queue_5_empty;
  assign sinkVec_queue_5_empty = _sinkVec_queue_fifo_5_empty;
  wire         sinkVec_queue_5_full;
  assign sinkVec_queue_5_full = _sinkVec_queue_fifo_5_full;
  wire         sinkVec_queue_6_empty;
  assign sinkVec_queue_6_empty = _sinkVec_queue_fifo_6_empty;
  wire         sinkVec_queue_6_full;
  assign sinkVec_queue_6_full = _sinkVec_queue_fifo_6_full;
  wire         sinkVec_queue_7_empty;
  assign sinkVec_queue_7_empty = _sinkVec_queue_fifo_7_empty;
  wire         sinkVec_queue_7_full;
  assign sinkVec_queue_7_full = _sinkVec_queue_fifo_7_full;
  assign accessDataSource_4_bits = _laneVec_2_vrfReadDataChannel;
  assign accessDataSource_5_bits = _laneVec_2_vrfReadDataChannel;
  wire         sinkVec_queue_8_empty;
  assign sinkVec_queue_8_empty = _sinkVec_queue_fifo_8_empty;
  wire         sinkVec_queue_8_full;
  assign sinkVec_queue_8_full = _sinkVec_queue_fifo_8_full;
  wire         sinkVec_queue_9_empty;
  assign sinkVec_queue_9_empty = _sinkVec_queue_fifo_9_empty;
  wire         sinkVec_queue_9_full;
  assign sinkVec_queue_9_full = _sinkVec_queue_fifo_9_full;
  wire         sinkVec_queue_10_empty;
  assign sinkVec_queue_10_empty = _sinkVec_queue_fifo_10_empty;
  wire         sinkVec_queue_10_full;
  assign sinkVec_queue_10_full = _sinkVec_queue_fifo_10_full;
  wire         sinkVec_queue_11_empty;
  assign sinkVec_queue_11_empty = _sinkVec_queue_fifo_11_empty;
  wire         sinkVec_queue_11_full;
  assign sinkVec_queue_11_full = _sinkVec_queue_fifo_11_full;
  assign accessDataSource_6_bits = _laneVec_3_vrfReadDataChannel;
  assign accessDataSource_7_bits = _laneVec_3_vrfReadDataChannel;
  wire         sinkVec_queue_12_empty;
  assign sinkVec_queue_12_empty = _sinkVec_queue_fifo_12_empty;
  wire         sinkVec_queue_12_full;
  assign sinkVec_queue_12_full = _sinkVec_queue_fifo_12_full;
  wire         sinkVec_queue_13_empty;
  assign sinkVec_queue_13_empty = _sinkVec_queue_fifo_13_empty;
  wire         sinkVec_queue_13_full;
  assign sinkVec_queue_13_full = _sinkVec_queue_fifo_13_full;
  wire         sinkVec_queue_14_empty;
  assign sinkVec_queue_14_empty = _sinkVec_queue_fifo_14_empty;
  wire         sinkVec_queue_14_full;
  assign sinkVec_queue_14_full = _sinkVec_queue_fifo_14_full;
  wire         sinkVec_queue_15_empty;
  assign sinkVec_queue_15_empty = _sinkVec_queue_fifo_15_empty;
  wire         sinkVec_queue_15_full;
  assign sinkVec_queue_15_full = _sinkVec_queue_fifo_15_full;
  assign accessDataSource_8_bits = _laneVec_4_vrfReadDataChannel;
  assign accessDataSource_9_bits = _laneVec_4_vrfReadDataChannel;
  wire         sinkVec_queue_16_empty;
  assign sinkVec_queue_16_empty = _sinkVec_queue_fifo_16_empty;
  wire         sinkVec_queue_16_full;
  assign sinkVec_queue_16_full = _sinkVec_queue_fifo_16_full;
  wire         sinkVec_queue_17_empty;
  assign sinkVec_queue_17_empty = _sinkVec_queue_fifo_17_empty;
  wire         sinkVec_queue_17_full;
  assign sinkVec_queue_17_full = _sinkVec_queue_fifo_17_full;
  wire         sinkVec_queue_18_empty;
  assign sinkVec_queue_18_empty = _sinkVec_queue_fifo_18_empty;
  wire         sinkVec_queue_18_full;
  assign sinkVec_queue_18_full = _sinkVec_queue_fifo_18_full;
  wire         sinkVec_queue_19_empty;
  assign sinkVec_queue_19_empty = _sinkVec_queue_fifo_19_empty;
  wire         sinkVec_queue_19_full;
  assign sinkVec_queue_19_full = _sinkVec_queue_fifo_19_full;
  assign accessDataSource_10_bits = _laneVec_5_vrfReadDataChannel;
  assign accessDataSource_11_bits = _laneVec_5_vrfReadDataChannel;
  wire         sinkVec_queue_20_empty;
  assign sinkVec_queue_20_empty = _sinkVec_queue_fifo_20_empty;
  wire         sinkVec_queue_20_full;
  assign sinkVec_queue_20_full = _sinkVec_queue_fifo_20_full;
  wire         sinkVec_queue_21_empty;
  assign sinkVec_queue_21_empty = _sinkVec_queue_fifo_21_empty;
  wire         sinkVec_queue_21_full;
  assign sinkVec_queue_21_full = _sinkVec_queue_fifo_21_full;
  wire         sinkVec_queue_22_empty;
  assign sinkVec_queue_22_empty = _sinkVec_queue_fifo_22_empty;
  wire         sinkVec_queue_22_full;
  assign sinkVec_queue_22_full = _sinkVec_queue_fifo_22_full;
  wire         sinkVec_queue_23_empty;
  assign sinkVec_queue_23_empty = _sinkVec_queue_fifo_23_empty;
  wire         sinkVec_queue_23_full;
  assign sinkVec_queue_23_full = _sinkVec_queue_fifo_23_full;
  assign accessDataSource_12_bits = _laneVec_6_vrfReadDataChannel;
  assign accessDataSource_13_bits = _laneVec_6_vrfReadDataChannel;
  wire         sinkVec_queue_24_empty;
  assign sinkVec_queue_24_empty = _sinkVec_queue_fifo_24_empty;
  wire         sinkVec_queue_24_full;
  assign sinkVec_queue_24_full = _sinkVec_queue_fifo_24_full;
  wire         sinkVec_queue_25_empty;
  assign sinkVec_queue_25_empty = _sinkVec_queue_fifo_25_empty;
  wire         sinkVec_queue_25_full;
  assign sinkVec_queue_25_full = _sinkVec_queue_fifo_25_full;
  wire         sinkVec_queue_26_empty;
  assign sinkVec_queue_26_empty = _sinkVec_queue_fifo_26_empty;
  wire         sinkVec_queue_26_full;
  assign sinkVec_queue_26_full = _sinkVec_queue_fifo_26_full;
  wire         sinkVec_queue_27_empty;
  assign sinkVec_queue_27_empty = _sinkVec_queue_fifo_27_empty;
  wire         sinkVec_queue_27_full;
  assign sinkVec_queue_27_full = _sinkVec_queue_fifo_27_full;
  assign accessDataSource_14_bits = _laneVec_7_vrfReadDataChannel;
  assign accessDataSource_15_bits = _laneVec_7_vrfReadDataChannel;
  wire         sinkVec_queue_28_empty;
  assign sinkVec_queue_28_empty = _sinkVec_queue_fifo_28_empty;
  wire         sinkVec_queue_28_full;
  assign sinkVec_queue_28_full = _sinkVec_queue_fifo_28_full;
  wire         sinkVec_queue_29_empty;
  assign sinkVec_queue_29_empty = _sinkVec_queue_fifo_29_empty;
  wire         sinkVec_queue_29_full;
  assign sinkVec_queue_29_full = _sinkVec_queue_fifo_29_full;
  wire         sinkVec_queue_30_empty;
  assign sinkVec_queue_30_empty = _sinkVec_queue_fifo_30_empty;
  wire         sinkVec_queue_30_full;
  assign sinkVec_queue_30_full = _sinkVec_queue_fifo_30_full;
  wire         sinkVec_queue_31_empty;
  assign sinkVec_queue_31_empty = _sinkVec_queue_fifo_31_empty;
  wire         sinkVec_queue_31_full;
  assign sinkVec_queue_31_full = _sinkVec_queue_fifo_31_full;
  assign accessDataSource_16_bits = _laneVec_8_vrfReadDataChannel;
  assign accessDataSource_17_bits = _laneVec_8_vrfReadDataChannel;
  wire         sinkVec_queue_32_empty;
  assign sinkVec_queue_32_empty = _sinkVec_queue_fifo_32_empty;
  wire         sinkVec_queue_32_full;
  assign sinkVec_queue_32_full = _sinkVec_queue_fifo_32_full;
  wire         sinkVec_queue_33_empty;
  assign sinkVec_queue_33_empty = _sinkVec_queue_fifo_33_empty;
  wire         sinkVec_queue_33_full;
  assign sinkVec_queue_33_full = _sinkVec_queue_fifo_33_full;
  wire         sinkVec_queue_34_empty;
  assign sinkVec_queue_34_empty = _sinkVec_queue_fifo_34_empty;
  wire         sinkVec_queue_34_full;
  assign sinkVec_queue_34_full = _sinkVec_queue_fifo_34_full;
  wire         sinkVec_queue_35_empty;
  assign sinkVec_queue_35_empty = _sinkVec_queue_fifo_35_empty;
  wire         sinkVec_queue_35_full;
  assign sinkVec_queue_35_full = _sinkVec_queue_fifo_35_full;
  assign accessDataSource_18_bits = _laneVec_9_vrfReadDataChannel;
  assign accessDataSource_19_bits = _laneVec_9_vrfReadDataChannel;
  wire         sinkVec_queue_36_empty;
  assign sinkVec_queue_36_empty = _sinkVec_queue_fifo_36_empty;
  wire         sinkVec_queue_36_full;
  assign sinkVec_queue_36_full = _sinkVec_queue_fifo_36_full;
  wire         sinkVec_queue_37_empty;
  assign sinkVec_queue_37_empty = _sinkVec_queue_fifo_37_empty;
  wire         sinkVec_queue_37_full;
  assign sinkVec_queue_37_full = _sinkVec_queue_fifo_37_full;
  wire         sinkVec_queue_38_empty;
  assign sinkVec_queue_38_empty = _sinkVec_queue_fifo_38_empty;
  wire         sinkVec_queue_38_full;
  assign sinkVec_queue_38_full = _sinkVec_queue_fifo_38_full;
  wire         sinkVec_queue_39_empty;
  assign sinkVec_queue_39_empty = _sinkVec_queue_fifo_39_empty;
  wire         sinkVec_queue_39_full;
  assign sinkVec_queue_39_full = _sinkVec_queue_fifo_39_full;
  assign accessDataSource_20_bits = _laneVec_10_vrfReadDataChannel;
  assign accessDataSource_21_bits = _laneVec_10_vrfReadDataChannel;
  wire         sinkVec_queue_40_empty;
  assign sinkVec_queue_40_empty = _sinkVec_queue_fifo_40_empty;
  wire         sinkVec_queue_40_full;
  assign sinkVec_queue_40_full = _sinkVec_queue_fifo_40_full;
  wire         sinkVec_queue_41_empty;
  assign sinkVec_queue_41_empty = _sinkVec_queue_fifo_41_empty;
  wire         sinkVec_queue_41_full;
  assign sinkVec_queue_41_full = _sinkVec_queue_fifo_41_full;
  wire         sinkVec_queue_42_empty;
  assign sinkVec_queue_42_empty = _sinkVec_queue_fifo_42_empty;
  wire         sinkVec_queue_42_full;
  assign sinkVec_queue_42_full = _sinkVec_queue_fifo_42_full;
  wire         sinkVec_queue_43_empty;
  assign sinkVec_queue_43_empty = _sinkVec_queue_fifo_43_empty;
  wire         sinkVec_queue_43_full;
  assign sinkVec_queue_43_full = _sinkVec_queue_fifo_43_full;
  assign accessDataSource_22_bits = _laneVec_11_vrfReadDataChannel;
  assign accessDataSource_23_bits = _laneVec_11_vrfReadDataChannel;
  wire         sinkVec_queue_44_empty;
  assign sinkVec_queue_44_empty = _sinkVec_queue_fifo_44_empty;
  wire         sinkVec_queue_44_full;
  assign sinkVec_queue_44_full = _sinkVec_queue_fifo_44_full;
  wire         sinkVec_queue_45_empty;
  assign sinkVec_queue_45_empty = _sinkVec_queue_fifo_45_empty;
  wire         sinkVec_queue_45_full;
  assign sinkVec_queue_45_full = _sinkVec_queue_fifo_45_full;
  wire         sinkVec_queue_46_empty;
  assign sinkVec_queue_46_empty = _sinkVec_queue_fifo_46_empty;
  wire         sinkVec_queue_46_full;
  assign sinkVec_queue_46_full = _sinkVec_queue_fifo_46_full;
  wire         sinkVec_queue_47_empty;
  assign sinkVec_queue_47_empty = _sinkVec_queue_fifo_47_empty;
  wire         sinkVec_queue_47_full;
  assign sinkVec_queue_47_full = _sinkVec_queue_fifo_47_full;
  assign accessDataSource_24_bits = _laneVec_12_vrfReadDataChannel;
  assign accessDataSource_25_bits = _laneVec_12_vrfReadDataChannel;
  wire         sinkVec_queue_48_empty;
  assign sinkVec_queue_48_empty = _sinkVec_queue_fifo_48_empty;
  wire         sinkVec_queue_48_full;
  assign sinkVec_queue_48_full = _sinkVec_queue_fifo_48_full;
  wire         sinkVec_queue_49_empty;
  assign sinkVec_queue_49_empty = _sinkVec_queue_fifo_49_empty;
  wire         sinkVec_queue_49_full;
  assign sinkVec_queue_49_full = _sinkVec_queue_fifo_49_full;
  wire         sinkVec_queue_50_empty;
  assign sinkVec_queue_50_empty = _sinkVec_queue_fifo_50_empty;
  wire         sinkVec_queue_50_full;
  assign sinkVec_queue_50_full = _sinkVec_queue_fifo_50_full;
  wire         sinkVec_queue_51_empty;
  assign sinkVec_queue_51_empty = _sinkVec_queue_fifo_51_empty;
  wire         sinkVec_queue_51_full;
  assign sinkVec_queue_51_full = _sinkVec_queue_fifo_51_full;
  assign accessDataSource_26_bits = _laneVec_13_vrfReadDataChannel;
  assign accessDataSource_27_bits = _laneVec_13_vrfReadDataChannel;
  wire         sinkVec_queue_52_empty;
  assign sinkVec_queue_52_empty = _sinkVec_queue_fifo_52_empty;
  wire         sinkVec_queue_52_full;
  assign sinkVec_queue_52_full = _sinkVec_queue_fifo_52_full;
  wire         sinkVec_queue_53_empty;
  assign sinkVec_queue_53_empty = _sinkVec_queue_fifo_53_empty;
  wire         sinkVec_queue_53_full;
  assign sinkVec_queue_53_full = _sinkVec_queue_fifo_53_full;
  wire         sinkVec_queue_54_empty;
  assign sinkVec_queue_54_empty = _sinkVec_queue_fifo_54_empty;
  wire         sinkVec_queue_54_full;
  assign sinkVec_queue_54_full = _sinkVec_queue_fifo_54_full;
  wire         sinkVec_queue_55_empty;
  assign sinkVec_queue_55_empty = _sinkVec_queue_fifo_55_empty;
  wire         sinkVec_queue_55_full;
  assign sinkVec_queue_55_full = _sinkVec_queue_fifo_55_full;
  assign accessDataSource_28_bits = _laneVec_14_vrfReadDataChannel;
  assign accessDataSource_29_bits = _laneVec_14_vrfReadDataChannel;
  wire         sinkVec_queue_56_empty;
  assign sinkVec_queue_56_empty = _sinkVec_queue_fifo_56_empty;
  wire         sinkVec_queue_56_full;
  assign sinkVec_queue_56_full = _sinkVec_queue_fifo_56_full;
  wire         sinkVec_queue_57_empty;
  assign sinkVec_queue_57_empty = _sinkVec_queue_fifo_57_empty;
  wire         sinkVec_queue_57_full;
  assign sinkVec_queue_57_full = _sinkVec_queue_fifo_57_full;
  wire         sinkVec_queue_58_empty;
  assign sinkVec_queue_58_empty = _sinkVec_queue_fifo_58_empty;
  wire         sinkVec_queue_58_full;
  assign sinkVec_queue_58_full = _sinkVec_queue_fifo_58_full;
  wire         sinkVec_queue_59_empty;
  assign sinkVec_queue_59_empty = _sinkVec_queue_fifo_59_empty;
  wire         sinkVec_queue_59_full;
  assign sinkVec_queue_59_full = _sinkVec_queue_fifo_59_full;
  assign accessDataSource_30_bits = _laneVec_15_vrfReadDataChannel;
  assign accessDataSource_31_bits = _laneVec_15_vrfReadDataChannel;
  wire         sinkVec_queue_60_empty;
  assign sinkVec_queue_60_empty = _sinkVec_queue_fifo_60_empty;
  wire         sinkVec_queue_60_full;
  assign sinkVec_queue_60_full = _sinkVec_queue_fifo_60_full;
  wire         sinkVec_queue_61_empty;
  assign sinkVec_queue_61_empty = _sinkVec_queue_fifo_61_empty;
  wire         sinkVec_queue_61_full;
  assign sinkVec_queue_61_full = _sinkVec_queue_fifo_61_full;
  wire         sinkVec_queue_62_empty;
  assign sinkVec_queue_62_empty = _sinkVec_queue_fifo_62_empty;
  wire         sinkVec_queue_62_full;
  assign sinkVec_queue_62_full = _sinkVec_queue_fifo_62_full;
  wire         sinkVec_queue_63_empty;
  assign sinkVec_queue_63_empty = _sinkVec_queue_fifo_63_empty;
  wire         sinkVec_queue_63_full;
  assign sinkVec_queue_63_full = _sinkVec_queue_fifo_63_full;
  LSU lsu (
    .clock                                               (clock),
    .reset                                               (reset),
    .request_ready                                       (_lsu_request_ready),
    .request_valid                                       (maskUnit_gatherData_ready & isLoadStoreType),
    .request_bits_instructionInformation_nf              (requestRegDequeue_bits_instruction[31:29]),
    .request_bits_instructionInformation_mew             (requestRegDequeue_bits_instruction[28]),
    .request_bits_instructionInformation_mop             (requestRegDequeue_bits_instruction[27:26]),
    .request_bits_instructionInformation_lumop           (requestRegDequeue_bits_instruction[24:20]),
    .request_bits_instructionInformation_eew             (vSewForLsu),
    .request_bits_instructionInformation_vs3             (requestRegDequeue_bits_instruction[11:7]),
    .request_bits_instructionInformation_isStore         (isStoreType),
    .request_bits_instructionInformation_maskedLoadStore (maskType),
    .request_bits_rs1Data                                (requestRegDequeue_bits_rs1Data),
    .request_bits_rs2Data                                (requestRegDequeue_bits_rs2Data),
    .request_bits_instructionIndex                       (requestReg_bits_instructionIndex),
    .v0UpdateVec_0_valid                                 (_laneVec_0_v0Update_valid),
    .v0UpdateVec_0_bits_data                             (_laneVec_0_v0Update_bits_data),
    .v0UpdateVec_0_bits_offset                           (_laneVec_0_v0Update_bits_offset),
    .v0UpdateVec_0_bits_mask                             (_laneVec_0_v0Update_bits_mask),
    .v0UpdateVec_1_valid                                 (_laneVec_1_v0Update_valid),
    .v0UpdateVec_1_bits_data                             (_laneVec_1_v0Update_bits_data),
    .v0UpdateVec_1_bits_offset                           (_laneVec_1_v0Update_bits_offset),
    .v0UpdateVec_1_bits_mask                             (_laneVec_1_v0Update_bits_mask),
    .v0UpdateVec_2_valid                                 (_laneVec_2_v0Update_valid),
    .v0UpdateVec_2_bits_data                             (_laneVec_2_v0Update_bits_data),
    .v0UpdateVec_2_bits_offset                           (_laneVec_2_v0Update_bits_offset),
    .v0UpdateVec_2_bits_mask                             (_laneVec_2_v0Update_bits_mask),
    .v0UpdateVec_3_valid                                 (_laneVec_3_v0Update_valid),
    .v0UpdateVec_3_bits_data                             (_laneVec_3_v0Update_bits_data),
    .v0UpdateVec_3_bits_offset                           (_laneVec_3_v0Update_bits_offset),
    .v0UpdateVec_3_bits_mask                             (_laneVec_3_v0Update_bits_mask),
    .v0UpdateVec_4_valid                                 (_laneVec_4_v0Update_valid),
    .v0UpdateVec_4_bits_data                             (_laneVec_4_v0Update_bits_data),
    .v0UpdateVec_4_bits_offset                           (_laneVec_4_v0Update_bits_offset),
    .v0UpdateVec_4_bits_mask                             (_laneVec_4_v0Update_bits_mask),
    .v0UpdateVec_5_valid                                 (_laneVec_5_v0Update_valid),
    .v0UpdateVec_5_bits_data                             (_laneVec_5_v0Update_bits_data),
    .v0UpdateVec_5_bits_offset                           (_laneVec_5_v0Update_bits_offset),
    .v0UpdateVec_5_bits_mask                             (_laneVec_5_v0Update_bits_mask),
    .v0UpdateVec_6_valid                                 (_laneVec_6_v0Update_valid),
    .v0UpdateVec_6_bits_data                             (_laneVec_6_v0Update_bits_data),
    .v0UpdateVec_6_bits_offset                           (_laneVec_6_v0Update_bits_offset),
    .v0UpdateVec_6_bits_mask                             (_laneVec_6_v0Update_bits_mask),
    .v0UpdateVec_7_valid                                 (_laneVec_7_v0Update_valid),
    .v0UpdateVec_7_bits_data                             (_laneVec_7_v0Update_bits_data),
    .v0UpdateVec_7_bits_offset                           (_laneVec_7_v0Update_bits_offset),
    .v0UpdateVec_7_bits_mask                             (_laneVec_7_v0Update_bits_mask),
    .v0UpdateVec_8_valid                                 (_laneVec_8_v0Update_valid),
    .v0UpdateVec_8_bits_data                             (_laneVec_8_v0Update_bits_data),
    .v0UpdateVec_8_bits_offset                           (_laneVec_8_v0Update_bits_offset),
    .v0UpdateVec_8_bits_mask                             (_laneVec_8_v0Update_bits_mask),
    .v0UpdateVec_9_valid                                 (_laneVec_9_v0Update_valid),
    .v0UpdateVec_9_bits_data                             (_laneVec_9_v0Update_bits_data),
    .v0UpdateVec_9_bits_offset                           (_laneVec_9_v0Update_bits_offset),
    .v0UpdateVec_9_bits_mask                             (_laneVec_9_v0Update_bits_mask),
    .v0UpdateVec_10_valid                                (_laneVec_10_v0Update_valid),
    .v0UpdateVec_10_bits_data                            (_laneVec_10_v0Update_bits_data),
    .v0UpdateVec_10_bits_offset                          (_laneVec_10_v0Update_bits_offset),
    .v0UpdateVec_10_bits_mask                            (_laneVec_10_v0Update_bits_mask),
    .v0UpdateVec_11_valid                                (_laneVec_11_v0Update_valid),
    .v0UpdateVec_11_bits_data                            (_laneVec_11_v0Update_bits_data),
    .v0UpdateVec_11_bits_offset                          (_laneVec_11_v0Update_bits_offset),
    .v0UpdateVec_11_bits_mask                            (_laneVec_11_v0Update_bits_mask),
    .v0UpdateVec_12_valid                                (_laneVec_12_v0Update_valid),
    .v0UpdateVec_12_bits_data                            (_laneVec_12_v0Update_bits_data),
    .v0UpdateVec_12_bits_offset                          (_laneVec_12_v0Update_bits_offset),
    .v0UpdateVec_12_bits_mask                            (_laneVec_12_v0Update_bits_mask),
    .v0UpdateVec_13_valid                                (_laneVec_13_v0Update_valid),
    .v0UpdateVec_13_bits_data                            (_laneVec_13_v0Update_bits_data),
    .v0UpdateVec_13_bits_offset                          (_laneVec_13_v0Update_bits_offset),
    .v0UpdateVec_13_bits_mask                            (_laneVec_13_v0Update_bits_mask),
    .v0UpdateVec_14_valid                                (_laneVec_14_v0Update_valid),
    .v0UpdateVec_14_bits_data                            (_laneVec_14_v0Update_bits_data),
    .v0UpdateVec_14_bits_offset                          (_laneVec_14_v0Update_bits_offset),
    .v0UpdateVec_14_bits_mask                            (_laneVec_14_v0Update_bits_mask),
    .v0UpdateVec_15_valid                                (_laneVec_15_v0Update_valid),
    .v0UpdateVec_15_bits_data                            (_laneVec_15_v0Update_bits_data),
    .v0UpdateVec_15_bits_offset                          (_laneVec_15_v0Update_bits_offset),
    .v0UpdateVec_15_bits_mask                            (_laneVec_15_v0Update_bits_mask),
    .axi4Port_aw_ready                                   (highBandwidthLoadStorePort_aw_ready_0),
    .axi4Port_aw_valid                                   (highBandwidthLoadStorePort_aw_valid_0),
    .axi4Port_aw_bits_id                                 (highBandwidthLoadStorePort_aw_bits_id_0),
    .axi4Port_aw_bits_addr                               (highBandwidthLoadStorePort_aw_bits_addr_0),
    .axi4Port_w_ready                                    (highBandwidthLoadStorePort_w_ready_0),
    .axi4Port_w_valid                                    (highBandwidthLoadStorePort_w_valid_0),
    .axi4Port_w_bits_data                                (highBandwidthLoadStorePort_w_bits_data_0),
    .axi4Port_w_bits_strb                                (highBandwidthLoadStorePort_w_bits_strb_0),
    .axi4Port_b_valid                                    (highBandwidthLoadStorePort_b_valid_0),
    .axi4Port_b_bits_id                                  (highBandwidthLoadStorePort_b_bits_id_0),
    .axi4Port_b_bits_resp                                (highBandwidthLoadStorePort_b_bits_resp_0),
    .axi4Port_ar_ready                                   (highBandwidthLoadStorePort_ar_ready_0),
    .axi4Port_ar_valid                                   (highBandwidthLoadStorePort_ar_valid_0),
    .axi4Port_ar_bits_addr                               (highBandwidthLoadStorePort_ar_bits_addr_0),
    .axi4Port_r_ready                                    (highBandwidthLoadStorePort_r_ready_0),
    .axi4Port_r_valid                                    (highBandwidthLoadStorePort_r_valid_0),
    .axi4Port_r_bits_id                                  (highBandwidthLoadStorePort_r_bits_id_0),
    .axi4Port_r_bits_data                                (highBandwidthLoadStorePort_r_bits_data_0),
    .axi4Port_r_bits_resp                                (highBandwidthLoadStorePort_r_bits_resp_0),
    .axi4Port_r_bits_last                                (highBandwidthLoadStorePort_r_bits_last_0),
    .simpleAccessPorts_aw_ready                          (indexedLoadStorePort_aw_ready_0),
    .simpleAccessPorts_aw_valid                          (indexedLoadStorePort_aw_valid_0),
    .simpleAccessPorts_aw_bits_id                        (indexedLoadStorePort_aw_bits_id_0),
    .simpleAccessPorts_aw_bits_addr                      (indexedLoadStorePort_aw_bits_addr_0),
    .simpleAccessPorts_aw_bits_size                      (indexedLoadStorePort_aw_bits_size_0),
    .simpleAccessPorts_w_ready                           (indexedLoadStorePort_w_ready_0),
    .simpleAccessPorts_w_valid                           (indexedLoadStorePort_w_valid_0),
    .simpleAccessPorts_w_bits_data                       (indexedLoadStorePort_w_bits_data_0),
    .simpleAccessPorts_w_bits_strb                       (indexedLoadStorePort_w_bits_strb_0),
    .simpleAccessPorts_b_valid                           (indexedLoadStorePort_b_valid_0),
    .simpleAccessPorts_b_bits_id                         (indexedLoadStorePort_b_bits_id_0),
    .simpleAccessPorts_b_bits_resp                       (indexedLoadStorePort_b_bits_resp_0),
    .simpleAccessPorts_ar_ready                          (indexedLoadStorePort_ar_ready_0),
    .simpleAccessPorts_ar_valid                          (indexedLoadStorePort_ar_valid_0),
    .simpleAccessPorts_ar_bits_addr                      (indexedLoadStorePort_ar_bits_addr_0),
    .simpleAccessPorts_r_ready                           (indexedLoadStorePort_r_ready_0),
    .simpleAccessPorts_r_valid                           (indexedLoadStorePort_r_valid_0),
    .simpleAccessPorts_r_bits_id                         (indexedLoadStorePort_r_bits_id_0),
    .simpleAccessPorts_r_bits_data                       (indexedLoadStorePort_r_bits_data_0),
    .simpleAccessPorts_r_bits_resp                       (indexedLoadStorePort_r_bits_resp_0),
    .simpleAccessPorts_r_bits_last                       (indexedLoadStorePort_r_bits_last_0),
    .vrfReadDataPorts_0_ready                            (x13_1_ready),
    .vrfReadDataPorts_0_valid                            (x13_1_valid),
    .vrfReadDataPorts_0_bits_vs                          (x13_1_bits_vs),
    .vrfReadDataPorts_0_bits_offset                      (x13_1_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex            (x13_1_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                            (x13_1_1_ready),
    .vrfReadDataPorts_1_valid                            (x13_1_1_valid),
    .vrfReadDataPorts_1_bits_vs                          (x13_1_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                      (x13_1_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex            (x13_1_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                            (x13_2_1_ready),
    .vrfReadDataPorts_2_valid                            (x13_2_1_valid),
    .vrfReadDataPorts_2_bits_vs                          (x13_2_1_bits_vs),
    .vrfReadDataPorts_2_bits_offset                      (x13_2_1_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex            (x13_2_1_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                            (x13_3_1_ready),
    .vrfReadDataPorts_3_valid                            (x13_3_1_valid),
    .vrfReadDataPorts_3_bits_vs                          (x13_3_1_bits_vs),
    .vrfReadDataPorts_3_bits_offset                      (x13_3_1_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex            (x13_3_1_bits_instructionIndex),
    .vrfReadDataPorts_4_ready                            (x13_4_1_ready),
    .vrfReadDataPorts_4_valid                            (x13_4_1_valid),
    .vrfReadDataPorts_4_bits_vs                          (x13_4_1_bits_vs),
    .vrfReadDataPorts_4_bits_offset                      (x13_4_1_bits_offset),
    .vrfReadDataPorts_4_bits_instructionIndex            (x13_4_1_bits_instructionIndex),
    .vrfReadDataPorts_5_ready                            (x13_5_1_ready),
    .vrfReadDataPorts_5_valid                            (x13_5_1_valid),
    .vrfReadDataPorts_5_bits_vs                          (x13_5_1_bits_vs),
    .vrfReadDataPorts_5_bits_offset                      (x13_5_1_bits_offset),
    .vrfReadDataPorts_5_bits_instructionIndex            (x13_5_1_bits_instructionIndex),
    .vrfReadDataPorts_6_ready                            (x13_6_1_ready),
    .vrfReadDataPorts_6_valid                            (x13_6_1_valid),
    .vrfReadDataPorts_6_bits_vs                          (x13_6_1_bits_vs),
    .vrfReadDataPorts_6_bits_offset                      (x13_6_1_bits_offset),
    .vrfReadDataPorts_6_bits_instructionIndex            (x13_6_1_bits_instructionIndex),
    .vrfReadDataPorts_7_ready                            (x13_7_1_ready),
    .vrfReadDataPorts_7_valid                            (x13_7_1_valid),
    .vrfReadDataPorts_7_bits_vs                          (x13_7_1_bits_vs),
    .vrfReadDataPorts_7_bits_offset                      (x13_7_1_bits_offset),
    .vrfReadDataPorts_7_bits_instructionIndex            (x13_7_1_bits_instructionIndex),
    .vrfReadDataPorts_8_ready                            (x13_8_1_ready),
    .vrfReadDataPorts_8_valid                            (x13_8_1_valid),
    .vrfReadDataPorts_8_bits_vs                          (x13_8_1_bits_vs),
    .vrfReadDataPorts_8_bits_offset                      (x13_8_1_bits_offset),
    .vrfReadDataPorts_8_bits_instructionIndex            (x13_8_1_bits_instructionIndex),
    .vrfReadDataPorts_9_ready                            (x13_9_1_ready),
    .vrfReadDataPorts_9_valid                            (x13_9_1_valid),
    .vrfReadDataPorts_9_bits_vs                          (x13_9_1_bits_vs),
    .vrfReadDataPorts_9_bits_offset                      (x13_9_1_bits_offset),
    .vrfReadDataPorts_9_bits_instructionIndex            (x13_9_1_bits_instructionIndex),
    .vrfReadDataPorts_10_ready                           (x13_10_1_ready),
    .vrfReadDataPorts_10_valid                           (x13_10_1_valid),
    .vrfReadDataPorts_10_bits_vs                         (x13_10_1_bits_vs),
    .vrfReadDataPorts_10_bits_offset                     (x13_10_1_bits_offset),
    .vrfReadDataPorts_10_bits_instructionIndex           (x13_10_1_bits_instructionIndex),
    .vrfReadDataPorts_11_ready                           (x13_11_1_ready),
    .vrfReadDataPorts_11_valid                           (x13_11_1_valid),
    .vrfReadDataPorts_11_bits_vs                         (x13_11_1_bits_vs),
    .vrfReadDataPorts_11_bits_offset                     (x13_11_1_bits_offset),
    .vrfReadDataPorts_11_bits_instructionIndex           (x13_11_1_bits_instructionIndex),
    .vrfReadDataPorts_12_ready                           (x13_12_1_ready),
    .vrfReadDataPorts_12_valid                           (x13_12_1_valid),
    .vrfReadDataPorts_12_bits_vs                         (x13_12_1_bits_vs),
    .vrfReadDataPorts_12_bits_offset                     (x13_12_1_bits_offset),
    .vrfReadDataPorts_12_bits_instructionIndex           (x13_12_1_bits_instructionIndex),
    .vrfReadDataPorts_13_ready                           (x13_13_1_ready),
    .vrfReadDataPorts_13_valid                           (x13_13_1_valid),
    .vrfReadDataPorts_13_bits_vs                         (x13_13_1_bits_vs),
    .vrfReadDataPorts_13_bits_offset                     (x13_13_1_bits_offset),
    .vrfReadDataPorts_13_bits_instructionIndex           (x13_13_1_bits_instructionIndex),
    .vrfReadDataPorts_14_ready                           (x13_14_1_ready),
    .vrfReadDataPorts_14_valid                           (x13_14_1_valid),
    .vrfReadDataPorts_14_bits_vs                         (x13_14_1_bits_vs),
    .vrfReadDataPorts_14_bits_offset                     (x13_14_1_bits_offset),
    .vrfReadDataPorts_14_bits_instructionIndex           (x13_14_1_bits_instructionIndex),
    .vrfReadDataPorts_15_ready                           (x13_15_1_ready),
    .vrfReadDataPorts_15_valid                           (x13_15_1_valid),
    .vrfReadDataPorts_15_bits_vs                         (x13_15_1_bits_vs),
    .vrfReadDataPorts_15_bits_offset                     (x13_15_1_bits_offset),
    .vrfReadDataPorts_15_bits_instructionIndex           (x13_15_1_bits_instructionIndex),
    .vrfReadResults_0_valid                              (shifterReg_17_0_valid),
    .vrfReadResults_0_bits                               (shifterReg_17_0_bits),
    .vrfReadResults_1_valid                              (shifterReg_19_0_valid),
    .vrfReadResults_1_bits                               (shifterReg_19_0_bits),
    .vrfReadResults_2_valid                              (shifterReg_21_0_valid),
    .vrfReadResults_2_bits                               (shifterReg_21_0_bits),
    .vrfReadResults_3_valid                              (shifterReg_23_0_valid),
    .vrfReadResults_3_bits                               (shifterReg_23_0_bits),
    .vrfReadResults_4_valid                              (shifterReg_25_0_valid),
    .vrfReadResults_4_bits                               (shifterReg_25_0_bits),
    .vrfReadResults_5_valid                              (shifterReg_27_0_valid),
    .vrfReadResults_5_bits                               (shifterReg_27_0_bits),
    .vrfReadResults_6_valid                              (shifterReg_29_0_valid),
    .vrfReadResults_6_bits                               (shifterReg_29_0_bits),
    .vrfReadResults_7_valid                              (shifterReg_31_0_valid),
    .vrfReadResults_7_bits                               (shifterReg_31_0_bits),
    .vrfReadResults_8_valid                              (shifterReg_33_0_valid),
    .vrfReadResults_8_bits                               (shifterReg_33_0_bits),
    .vrfReadResults_9_valid                              (shifterReg_35_0_valid),
    .vrfReadResults_9_bits                               (shifterReg_35_0_bits),
    .vrfReadResults_10_valid                             (shifterReg_37_0_valid),
    .vrfReadResults_10_bits                              (shifterReg_37_0_bits),
    .vrfReadResults_11_valid                             (shifterReg_39_0_valid),
    .vrfReadResults_11_bits                              (shifterReg_39_0_bits),
    .vrfReadResults_12_valid                             (shifterReg_41_0_valid),
    .vrfReadResults_12_bits                              (shifterReg_41_0_bits),
    .vrfReadResults_13_valid                             (shifterReg_43_0_valid),
    .vrfReadResults_13_bits                              (shifterReg_43_0_bits),
    .vrfReadResults_14_valid                             (shifterReg_45_0_valid),
    .vrfReadResults_14_bits                              (shifterReg_45_0_bits),
    .vrfReadResults_15_valid                             (shifterReg_47_0_valid),
    .vrfReadResults_15_bits                              (shifterReg_47_0_bits),
    .vrfWritePort_0_ready                                (x22_1_ready),
    .vrfWritePort_0_valid                                (_lsu_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                              (_lsu_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                          (x22_1_bits_offset),
    .vrfWritePort_0_bits_mask                            (_lsu_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                            (x22_1_bits_data),
    .vrfWritePort_0_bits_last                            (x22_1_bits_last),
    .vrfWritePort_0_bits_instructionIndex                (_lsu_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                (x22_1_1_ready),
    .vrfWritePort_1_valid                                (_lsu_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                              (_lsu_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                          (x22_1_1_bits_offset),
    .vrfWritePort_1_bits_mask                            (_lsu_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                            (x22_1_1_bits_data),
    .vrfWritePort_1_bits_last                            (x22_1_1_bits_last),
    .vrfWritePort_1_bits_instructionIndex                (_lsu_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                (x22_2_1_ready),
    .vrfWritePort_2_valid                                (_lsu_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                              (_lsu_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                          (x22_2_1_bits_offset),
    .vrfWritePort_2_bits_mask                            (_lsu_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                            (x22_2_1_bits_data),
    .vrfWritePort_2_bits_last                            (x22_2_1_bits_last),
    .vrfWritePort_2_bits_instructionIndex                (_lsu_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                (x22_3_1_ready),
    .vrfWritePort_3_valid                                (_lsu_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                              (_lsu_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                          (x22_3_1_bits_offset),
    .vrfWritePort_3_bits_mask                            (_lsu_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                            (x22_3_1_bits_data),
    .vrfWritePort_3_bits_last                            (x22_3_1_bits_last),
    .vrfWritePort_3_bits_instructionIndex                (_lsu_vrfWritePort_3_bits_instructionIndex),
    .vrfWritePort_4_ready                                (x22_4_1_ready),
    .vrfWritePort_4_valid                                (_lsu_vrfWritePort_4_valid),
    .vrfWritePort_4_bits_vd                              (_lsu_vrfWritePort_4_bits_vd),
    .vrfWritePort_4_bits_offset                          (x22_4_1_bits_offset),
    .vrfWritePort_4_bits_mask                            (_lsu_vrfWritePort_4_bits_mask),
    .vrfWritePort_4_bits_data                            (x22_4_1_bits_data),
    .vrfWritePort_4_bits_last                            (x22_4_1_bits_last),
    .vrfWritePort_4_bits_instructionIndex                (_lsu_vrfWritePort_4_bits_instructionIndex),
    .vrfWritePort_5_ready                                (x22_5_1_ready),
    .vrfWritePort_5_valid                                (_lsu_vrfWritePort_5_valid),
    .vrfWritePort_5_bits_vd                              (_lsu_vrfWritePort_5_bits_vd),
    .vrfWritePort_5_bits_offset                          (x22_5_1_bits_offset),
    .vrfWritePort_5_bits_mask                            (_lsu_vrfWritePort_5_bits_mask),
    .vrfWritePort_5_bits_data                            (x22_5_1_bits_data),
    .vrfWritePort_5_bits_last                            (x22_5_1_bits_last),
    .vrfWritePort_5_bits_instructionIndex                (_lsu_vrfWritePort_5_bits_instructionIndex),
    .vrfWritePort_6_ready                                (x22_6_1_ready),
    .vrfWritePort_6_valid                                (_lsu_vrfWritePort_6_valid),
    .vrfWritePort_6_bits_vd                              (_lsu_vrfWritePort_6_bits_vd),
    .vrfWritePort_6_bits_offset                          (x22_6_1_bits_offset),
    .vrfWritePort_6_bits_mask                            (_lsu_vrfWritePort_6_bits_mask),
    .vrfWritePort_6_bits_data                            (x22_6_1_bits_data),
    .vrfWritePort_6_bits_last                            (x22_6_1_bits_last),
    .vrfWritePort_6_bits_instructionIndex                (_lsu_vrfWritePort_6_bits_instructionIndex),
    .vrfWritePort_7_ready                                (x22_7_1_ready),
    .vrfWritePort_7_valid                                (_lsu_vrfWritePort_7_valid),
    .vrfWritePort_7_bits_vd                              (_lsu_vrfWritePort_7_bits_vd),
    .vrfWritePort_7_bits_offset                          (x22_7_1_bits_offset),
    .vrfWritePort_7_bits_mask                            (_lsu_vrfWritePort_7_bits_mask),
    .vrfWritePort_7_bits_data                            (x22_7_1_bits_data),
    .vrfWritePort_7_bits_last                            (x22_7_1_bits_last),
    .vrfWritePort_7_bits_instructionIndex                (_lsu_vrfWritePort_7_bits_instructionIndex),
    .vrfWritePort_8_ready                                (x22_8_1_ready),
    .vrfWritePort_8_valid                                (_lsu_vrfWritePort_8_valid),
    .vrfWritePort_8_bits_vd                              (_lsu_vrfWritePort_8_bits_vd),
    .vrfWritePort_8_bits_offset                          (x22_8_1_bits_offset),
    .vrfWritePort_8_bits_mask                            (_lsu_vrfWritePort_8_bits_mask),
    .vrfWritePort_8_bits_data                            (x22_8_1_bits_data),
    .vrfWritePort_8_bits_last                            (x22_8_1_bits_last),
    .vrfWritePort_8_bits_instructionIndex                (_lsu_vrfWritePort_8_bits_instructionIndex),
    .vrfWritePort_9_ready                                (x22_9_1_ready),
    .vrfWritePort_9_valid                                (_lsu_vrfWritePort_9_valid),
    .vrfWritePort_9_bits_vd                              (_lsu_vrfWritePort_9_bits_vd),
    .vrfWritePort_9_bits_offset                          (x22_9_1_bits_offset),
    .vrfWritePort_9_bits_mask                            (_lsu_vrfWritePort_9_bits_mask),
    .vrfWritePort_9_bits_data                            (x22_9_1_bits_data),
    .vrfWritePort_9_bits_last                            (x22_9_1_bits_last),
    .vrfWritePort_9_bits_instructionIndex                (_lsu_vrfWritePort_9_bits_instructionIndex),
    .vrfWritePort_10_ready                               (x22_10_1_ready),
    .vrfWritePort_10_valid                               (_lsu_vrfWritePort_10_valid),
    .vrfWritePort_10_bits_vd                             (_lsu_vrfWritePort_10_bits_vd),
    .vrfWritePort_10_bits_offset                         (x22_10_1_bits_offset),
    .vrfWritePort_10_bits_mask                           (_lsu_vrfWritePort_10_bits_mask),
    .vrfWritePort_10_bits_data                           (x22_10_1_bits_data),
    .vrfWritePort_10_bits_last                           (x22_10_1_bits_last),
    .vrfWritePort_10_bits_instructionIndex               (_lsu_vrfWritePort_10_bits_instructionIndex),
    .vrfWritePort_11_ready                               (x22_11_1_ready),
    .vrfWritePort_11_valid                               (_lsu_vrfWritePort_11_valid),
    .vrfWritePort_11_bits_vd                             (_lsu_vrfWritePort_11_bits_vd),
    .vrfWritePort_11_bits_offset                         (x22_11_1_bits_offset),
    .vrfWritePort_11_bits_mask                           (_lsu_vrfWritePort_11_bits_mask),
    .vrfWritePort_11_bits_data                           (x22_11_1_bits_data),
    .vrfWritePort_11_bits_last                           (x22_11_1_bits_last),
    .vrfWritePort_11_bits_instructionIndex               (_lsu_vrfWritePort_11_bits_instructionIndex),
    .vrfWritePort_12_ready                               (x22_12_1_ready),
    .vrfWritePort_12_valid                               (_lsu_vrfWritePort_12_valid),
    .vrfWritePort_12_bits_vd                             (_lsu_vrfWritePort_12_bits_vd),
    .vrfWritePort_12_bits_offset                         (x22_12_1_bits_offset),
    .vrfWritePort_12_bits_mask                           (_lsu_vrfWritePort_12_bits_mask),
    .vrfWritePort_12_bits_data                           (x22_12_1_bits_data),
    .vrfWritePort_12_bits_last                           (x22_12_1_bits_last),
    .vrfWritePort_12_bits_instructionIndex               (_lsu_vrfWritePort_12_bits_instructionIndex),
    .vrfWritePort_13_ready                               (x22_13_1_ready),
    .vrfWritePort_13_valid                               (_lsu_vrfWritePort_13_valid),
    .vrfWritePort_13_bits_vd                             (_lsu_vrfWritePort_13_bits_vd),
    .vrfWritePort_13_bits_offset                         (x22_13_1_bits_offset),
    .vrfWritePort_13_bits_mask                           (_lsu_vrfWritePort_13_bits_mask),
    .vrfWritePort_13_bits_data                           (x22_13_1_bits_data),
    .vrfWritePort_13_bits_last                           (x22_13_1_bits_last),
    .vrfWritePort_13_bits_instructionIndex               (_lsu_vrfWritePort_13_bits_instructionIndex),
    .vrfWritePort_14_ready                               (x22_14_1_ready),
    .vrfWritePort_14_valid                               (_lsu_vrfWritePort_14_valid),
    .vrfWritePort_14_bits_vd                             (_lsu_vrfWritePort_14_bits_vd),
    .vrfWritePort_14_bits_offset                         (x22_14_1_bits_offset),
    .vrfWritePort_14_bits_mask                           (_lsu_vrfWritePort_14_bits_mask),
    .vrfWritePort_14_bits_data                           (x22_14_1_bits_data),
    .vrfWritePort_14_bits_last                           (x22_14_1_bits_last),
    .vrfWritePort_14_bits_instructionIndex               (_lsu_vrfWritePort_14_bits_instructionIndex),
    .vrfWritePort_15_ready                               (x22_15_1_ready),
    .vrfWritePort_15_valid                               (_lsu_vrfWritePort_15_valid),
    .vrfWritePort_15_bits_vd                             (_lsu_vrfWritePort_15_bits_vd),
    .vrfWritePort_15_bits_offset                         (x22_15_1_bits_offset),
    .vrfWritePort_15_bits_mask                           (_lsu_vrfWritePort_15_bits_mask),
    .vrfWritePort_15_bits_data                           (x22_15_1_bits_data),
    .vrfWritePort_15_bits_last                           (x22_15_1_bits_last),
    .vrfWritePort_15_bits_instructionIndex               (_lsu_vrfWritePort_15_bits_instructionIndex),
    .writeRelease_0                                      (pipe_out_valid),
    .writeRelease_1                                      (pipe_out_2_valid),
    .writeRelease_2                                      (pipe_out_4_valid),
    .writeRelease_3                                      (pipe_out_6_valid),
    .writeRelease_4                                      (pipe_out_8_valid),
    .writeRelease_5                                      (pipe_out_10_valid),
    .writeRelease_6                                      (pipe_out_12_valid),
    .writeRelease_7                                      (pipe_out_14_valid),
    .writeRelease_8                                      (pipe_out_16_valid),
    .writeRelease_9                                      (pipe_out_18_valid),
    .writeRelease_10                                     (pipe_out_20_valid),
    .writeRelease_11                                     (pipe_out_22_valid),
    .writeRelease_12                                     (pipe_out_24_valid),
    .writeRelease_13                                     (pipe_out_26_valid),
    .writeRelease_14                                     (pipe_out_28_valid),
    .writeRelease_15                                     (pipe_out_30_valid),
    .dataInWriteQueue_0                                  (_lsu_dataInWriteQueue_0),
    .dataInWriteQueue_1                                  (_lsu_dataInWriteQueue_1),
    .dataInWriteQueue_2                                  (_lsu_dataInWriteQueue_2),
    .dataInWriteQueue_3                                  (_lsu_dataInWriteQueue_3),
    .dataInWriteQueue_4                                  (_lsu_dataInWriteQueue_4),
    .dataInWriteQueue_5                                  (_lsu_dataInWriteQueue_5),
    .dataInWriteQueue_6                                  (_lsu_dataInWriteQueue_6),
    .dataInWriteQueue_7                                  (_lsu_dataInWriteQueue_7),
    .dataInWriteQueue_8                                  (_lsu_dataInWriteQueue_8),
    .dataInWriteQueue_9                                  (_lsu_dataInWriteQueue_9),
    .dataInWriteQueue_10                                 (_lsu_dataInWriteQueue_10),
    .dataInWriteQueue_11                                 (_lsu_dataInWriteQueue_11),
    .dataInWriteQueue_12                                 (_lsu_dataInWriteQueue_12),
    .dataInWriteQueue_13                                 (_lsu_dataInWriteQueue_13),
    .dataInWriteQueue_14                                 (_lsu_dataInWriteQueue_14),
    .dataInWriteQueue_15                                 (_lsu_dataInWriteQueue_15),
    .csrInterface_vl                                     (evlForLsu[11:0]),
    .csrInterface_vStart                                 (requestRegCSR_vStart),
    .csrInterface_vlmul                                  (requestRegCSR_vlmul),
    .csrInterface_vSew                                   (requestRegCSR_vSew),
    .csrInterface_vxrm                                   (requestRegCSR_vxrm),
    .csrInterface_vta                                    (requestRegCSR_vta),
    .csrInterface_vma                                    (requestRegCSR_vma),
    .offsetReadResult_0_valid                            (_laneVec_0_maskUnitRequest_valid & _laneVec_0_maskRequestToLSU),
    .offsetReadResult_0_bits                             (_laneVec_0_maskUnitRequest_bits_source2),
    .offsetReadResult_1_valid                            (_laneVec_1_maskUnitRequest_valid & _laneVec_1_maskRequestToLSU),
    .offsetReadResult_1_bits                             (_laneVec_1_maskUnitRequest_bits_source2),
    .offsetReadResult_2_valid                            (_laneVec_2_maskUnitRequest_valid & _laneVec_2_maskRequestToLSU),
    .offsetReadResult_2_bits                             (_laneVec_2_maskUnitRequest_bits_source2),
    .offsetReadResult_3_valid                            (_laneVec_3_maskUnitRequest_valid & _laneVec_3_maskRequestToLSU),
    .offsetReadResult_3_bits                             (_laneVec_3_maskUnitRequest_bits_source2),
    .offsetReadResult_4_valid                            (_laneVec_4_maskUnitRequest_valid & _laneVec_4_maskRequestToLSU),
    .offsetReadResult_4_bits                             (_laneVec_4_maskUnitRequest_bits_source2),
    .offsetReadResult_5_valid                            (_laneVec_5_maskUnitRequest_valid & _laneVec_5_maskRequestToLSU),
    .offsetReadResult_5_bits                             (_laneVec_5_maskUnitRequest_bits_source2),
    .offsetReadResult_6_valid                            (_laneVec_6_maskUnitRequest_valid & _laneVec_6_maskRequestToLSU),
    .offsetReadResult_6_bits                             (_laneVec_6_maskUnitRequest_bits_source2),
    .offsetReadResult_7_valid                            (_laneVec_7_maskUnitRequest_valid & _laneVec_7_maskRequestToLSU),
    .offsetReadResult_7_bits                             (_laneVec_7_maskUnitRequest_bits_source2),
    .offsetReadResult_8_valid                            (_laneVec_8_maskUnitRequest_valid & _laneVec_8_maskRequestToLSU),
    .offsetReadResult_8_bits                             (_laneVec_8_maskUnitRequest_bits_source2),
    .offsetReadResult_9_valid                            (_laneVec_9_maskUnitRequest_valid & _laneVec_9_maskRequestToLSU),
    .offsetReadResult_9_bits                             (_laneVec_9_maskUnitRequest_bits_source2),
    .offsetReadResult_10_valid                           (_laneVec_10_maskUnitRequest_valid & _laneVec_10_maskRequestToLSU),
    .offsetReadResult_10_bits                            (_laneVec_10_maskUnitRequest_bits_source2),
    .offsetReadResult_11_valid                           (_laneVec_11_maskUnitRequest_valid & _laneVec_11_maskRequestToLSU),
    .offsetReadResult_11_bits                            (_laneVec_11_maskUnitRequest_bits_source2),
    .offsetReadResult_12_valid                           (_laneVec_12_maskUnitRequest_valid & _laneVec_12_maskRequestToLSU),
    .offsetReadResult_12_bits                            (_laneVec_12_maskUnitRequest_bits_source2),
    .offsetReadResult_13_valid                           (_laneVec_13_maskUnitRequest_valid & _laneVec_13_maskRequestToLSU),
    .offsetReadResult_13_bits                            (_laneVec_13_maskUnitRequest_bits_source2),
    .offsetReadResult_14_valid                           (_laneVec_14_maskUnitRequest_valid & _laneVec_14_maskRequestToLSU),
    .offsetReadResult_14_bits                            (_laneVec_14_maskUnitRequest_bits_source2),
    .offsetReadResult_15_valid                           (_laneVec_15_maskUnitRequest_valid & _laneVec_15_maskRequestToLSU),
    .offsetReadResult_15_bits                            (_laneVec_15_maskUnitRequest_bits_source2),
    .lastReport                                          (_lsu_lastReport),
    .tokenIO_offsetGroupRelease                          (_lsu_tokenIO_offsetGroupRelease)
  );
  VectorDecoder decode (
    .decodeInput                        (issue_bits_instruction_0),
    .decodeResult_orderReduce           (_decode_decodeResult_orderReduce),
    .decodeResult_floatMul              (_decode_decodeResult_floatMul),
    .decodeResult_fpExecutionType       (_decode_decodeResult_fpExecutionType),
    .decodeResult_float                 (_decode_decodeResult_float),
    .decodeResult_specialSlot           (_decode_decodeResult_specialSlot),
    .decodeResult_topUop                (_decode_decodeResult_topUop),
    .decodeResult_popCount              (_decode_decodeResult_popCount),
    .decodeResult_ffo                   (_decode_decodeResult_ffo),
    .decodeResult_average               (_decode_decodeResult_average),
    .decodeResult_reverse               (_decode_decodeResult_reverse),
    .decodeResult_dontNeedExecuteInLane (_decode_decodeResult_dontNeedExecuteInLane),
    .decodeResult_scheduler             (_decode_decodeResult_scheduler),
    .decodeResult_sReadVD               (_decode_decodeResult_sReadVD),
    .decodeResult_vtype                 (_decode_decodeResult_vtype),
    .decodeResult_sWrite                (_decode_decodeResult_sWrite),
    .decodeResult_crossRead             (_decode_decodeResult_crossRead),
    .decodeResult_crossWrite            (_decode_decodeResult_crossWrite),
    .decodeResult_maskUnit              (_decode_decodeResult_maskUnit),
    .decodeResult_special               (_decode_decodeResult_special),
    .decodeResult_saturate              (_decode_decodeResult_saturate),
    .decodeResult_vwmacc                (_decode_decodeResult_vwmacc),
    .decodeResult_readOnly              (_decode_decodeResult_readOnly),
    .decodeResult_maskSource            (_decode_decodeResult_maskSource),
    .decodeResult_maskDestination       (_decode_decodeResult_maskDestination),
    .decodeResult_maskLogic             (_decode_decodeResult_maskLogic),
    .decodeResult_uop                   (_decode_decodeResult_uop),
    .decodeResult_iota                  (_decode_decodeResult_iota),
    .decodeResult_mv                    (_decode_decodeResult_mv),
    .decodeResult_extend                (_decode_decodeResult_extend),
    .decodeResult_unOrderWrite          (_decode_decodeResult_unOrderWrite),
    .decodeResult_compress              (_decode_decodeResult_compress),
    .decodeResult_gather16              (_decode_decodeResult_gather16),
    .decodeResult_gather                (_decode_decodeResult_gather),
    .decodeResult_slid                  (_decode_decodeResult_slid),
    .decodeResult_targetRd              (_decode_decodeResult_targetRd),
    .decodeResult_widenReduce           (_decode_decodeResult_widenReduce),
    .decodeResult_red                   (_decode_decodeResult_red),
    .decodeResult_nr                    (_decode_decodeResult_nr),
    .decodeResult_itype                 (_decode_decodeResult_itype),
    .decodeResult_unsigned1             (_decode_decodeResult_unsigned1),
    .decodeResult_unsigned0             (_decode_decodeResult_unsigned0),
    .decodeResult_other                 (_decode_decodeResult_other),
    .decodeResult_multiCycle            (_decode_decodeResult_multiCycle),
    .decodeResult_divider               (_decode_decodeResult_divider),
    .decodeResult_multiplier            (_decode_decodeResult_multiplier),
    .decodeResult_shift                 (_decode_decodeResult_shift),
    .decodeResult_adder                 (_decode_decodeResult_adder),
    .decodeResult_logic                 (_decode_decodeResult_logic)
  );
  MaskUnit maskUnit (
    .clock                                           (clock),
    .reset                                           (reset),
    .instReq_valid                                   (maskUnit_gatherData_ready & requestReg_bits_decodeResult_maskUnit),
    .instReq_bits_instructionIndex                   (requestReg_bits_instructionIndex),
    .instReq_bits_decodeResult_orderReduce           (requestReg_bits_decodeResult_orderReduce),
    .instReq_bits_decodeResult_floatMul              (requestReg_bits_decodeResult_floatMul),
    .instReq_bits_decodeResult_fpExecutionType       (requestReg_bits_decodeResult_fpExecutionType),
    .instReq_bits_decodeResult_float                 (requestReg_bits_decodeResult_float),
    .instReq_bits_decodeResult_specialSlot           (requestReg_bits_decodeResult_specialSlot),
    .instReq_bits_decodeResult_topUop                (requestReg_bits_decodeResult_topUop),
    .instReq_bits_decodeResult_popCount              (requestReg_bits_decodeResult_popCount),
    .instReq_bits_decodeResult_ffo                   (requestReg_bits_decodeResult_ffo),
    .instReq_bits_decodeResult_average               (requestReg_bits_decodeResult_average),
    .instReq_bits_decodeResult_reverse               (requestReg_bits_decodeResult_reverse),
    .instReq_bits_decodeResult_dontNeedExecuteInLane (requestReg_bits_decodeResult_dontNeedExecuteInLane),
    .instReq_bits_decodeResult_scheduler             (requestReg_bits_decodeResult_scheduler),
    .instReq_bits_decodeResult_sReadVD               (requestReg_bits_decodeResult_sReadVD),
    .instReq_bits_decodeResult_vtype                 (requestReg_bits_decodeResult_vtype),
    .instReq_bits_decodeResult_sWrite                (requestReg_bits_decodeResult_sWrite),
    .instReq_bits_decodeResult_crossRead             (requestReg_bits_decodeResult_crossRead),
    .instReq_bits_decodeResult_crossWrite            (requestReg_bits_decodeResult_crossWrite),
    .instReq_bits_decodeResult_maskUnit              (requestReg_bits_decodeResult_maskUnit),
    .instReq_bits_decodeResult_special               (requestReg_bits_decodeResult_special),
    .instReq_bits_decodeResult_saturate              (requestReg_bits_decodeResult_saturate),
    .instReq_bits_decodeResult_vwmacc                (requestReg_bits_decodeResult_vwmacc),
    .instReq_bits_decodeResult_readOnly              (requestReg_bits_decodeResult_readOnly),
    .instReq_bits_decodeResult_maskSource            (requestReg_bits_decodeResult_maskSource),
    .instReq_bits_decodeResult_maskDestination       (requestReg_bits_decodeResult_maskDestination),
    .instReq_bits_decodeResult_maskLogic             (requestReg_bits_decodeResult_maskLogic),
    .instReq_bits_decodeResult_uop                   (requestReg_bits_decodeResult_uop),
    .instReq_bits_decodeResult_iota                  (requestReg_bits_decodeResult_iota),
    .instReq_bits_decodeResult_mv                    (requestReg_bits_decodeResult_mv),
    .instReq_bits_decodeResult_extend                (requestReg_bits_decodeResult_extend),
    .instReq_bits_decodeResult_unOrderWrite          (requestReg_bits_decodeResult_unOrderWrite),
    .instReq_bits_decodeResult_compress              (requestReg_bits_decodeResult_compress),
    .instReq_bits_decodeResult_gather16              (requestReg_bits_decodeResult_gather16),
    .instReq_bits_decodeResult_gather                (requestReg_bits_decodeResult_gather),
    .instReq_bits_decodeResult_slid                  (requestReg_bits_decodeResult_slid),
    .instReq_bits_decodeResult_targetRd              (requestReg_bits_decodeResult_targetRd),
    .instReq_bits_decodeResult_widenReduce           (requestReg_bits_decodeResult_widenReduce),
    .instReq_bits_decodeResult_red                   (requestReg_bits_decodeResult_red),
    .instReq_bits_decodeResult_nr                    (requestReg_bits_decodeResult_nr),
    .instReq_bits_decodeResult_itype                 (requestReg_bits_decodeResult_itype),
    .instReq_bits_decodeResult_unsigned1             (requestReg_bits_decodeResult_unsigned1),
    .instReq_bits_decodeResult_unsigned0             (requestReg_bits_decodeResult_unsigned0),
    .instReq_bits_decodeResult_other                 (requestReg_bits_decodeResult_other),
    .instReq_bits_decodeResult_multiCycle            (requestReg_bits_decodeResult_multiCycle),
    .instReq_bits_decodeResult_divider               (requestReg_bits_decodeResult_divider),
    .instReq_bits_decodeResult_multiplier            (requestReg_bits_decodeResult_multiplier),
    .instReq_bits_decodeResult_shift                 (requestReg_bits_decodeResult_shift),
    .instReq_bits_decodeResult_adder                 (requestReg_bits_decodeResult_adder),
    .instReq_bits_decodeResult_logic                 (requestReg_bits_decodeResult_logic),
    .instReq_bits_readFromScala                      (requestReg_bits_decodeResult_itype ? {27'h0, imm} : requestRegDequeue_bits_rs1Data),
    .instReq_bits_sew                                (requestRegCSR_vSew),
    .instReq_bits_vlmul                              (requestRegCSR_vlmul),
    .instReq_bits_maskType                           (maskType),
    .instReq_bits_vxrm                               ({1'h0, requestRegCSR_vxrm}),
    .instReq_bits_vs2                                (requestRegDequeue_bits_instruction[24:20]),
    .instReq_bits_vs1                                (requestRegDequeue_bits_instruction[19:15]),
    .instReq_bits_vd                                 (requestRegDequeue_bits_instruction[11:7]),
    .instReq_bits_vl                                 (requestRegCSR_vl),
    .exeReq_0_valid                                  (_laneVec_0_maskUnitRequest_valid & ~_laneVec_0_maskRequestToLSU),
    .exeReq_0_bits_source1                           (_laneVec_0_maskUnitRequest_bits_source1),
    .exeReq_0_bits_source2                           (_laneVec_0_maskUnitRequest_bits_source2),
    .exeReq_0_bits_index                             (_laneVec_0_maskUnitRequest_bits_index),
    .exeReq_0_bits_ffo                               (_laneVec_0_maskUnitRequest_bits_ffo),
    .exeReq_0_bits_fpReduceValid                     (_laneVec_0_maskUnitRequest_bits_fpReduceValid),
    .exeReq_1_valid                                  (_laneVec_1_maskUnitRequest_valid & ~_laneVec_1_maskRequestToLSU),
    .exeReq_1_bits_source1                           (_laneVec_1_maskUnitRequest_bits_source1),
    .exeReq_1_bits_source2                           (_laneVec_1_maskUnitRequest_bits_source2),
    .exeReq_1_bits_index                             (_laneVec_1_maskUnitRequest_bits_index),
    .exeReq_1_bits_ffo                               (_laneVec_1_maskUnitRequest_bits_ffo),
    .exeReq_1_bits_fpReduceValid                     (_laneVec_1_maskUnitRequest_bits_fpReduceValid),
    .exeReq_2_valid                                  (_laneVec_2_maskUnitRequest_valid & ~_laneVec_2_maskRequestToLSU),
    .exeReq_2_bits_source1                           (_laneVec_2_maskUnitRequest_bits_source1),
    .exeReq_2_bits_source2                           (_laneVec_2_maskUnitRequest_bits_source2),
    .exeReq_2_bits_index                             (_laneVec_2_maskUnitRequest_bits_index),
    .exeReq_2_bits_ffo                               (_laneVec_2_maskUnitRequest_bits_ffo),
    .exeReq_2_bits_fpReduceValid                     (_laneVec_2_maskUnitRequest_bits_fpReduceValid),
    .exeReq_3_valid                                  (_laneVec_3_maskUnitRequest_valid & ~_laneVec_3_maskRequestToLSU),
    .exeReq_3_bits_source1                           (_laneVec_3_maskUnitRequest_bits_source1),
    .exeReq_3_bits_source2                           (_laneVec_3_maskUnitRequest_bits_source2),
    .exeReq_3_bits_index                             (_laneVec_3_maskUnitRequest_bits_index),
    .exeReq_3_bits_ffo                               (_laneVec_3_maskUnitRequest_bits_ffo),
    .exeReq_3_bits_fpReduceValid                     (_laneVec_3_maskUnitRequest_bits_fpReduceValid),
    .exeReq_4_valid                                  (_laneVec_4_maskUnitRequest_valid & ~_laneVec_4_maskRequestToLSU),
    .exeReq_4_bits_source1                           (_laneVec_4_maskUnitRequest_bits_source1),
    .exeReq_4_bits_source2                           (_laneVec_4_maskUnitRequest_bits_source2),
    .exeReq_4_bits_index                             (_laneVec_4_maskUnitRequest_bits_index),
    .exeReq_4_bits_ffo                               (_laneVec_4_maskUnitRequest_bits_ffo),
    .exeReq_4_bits_fpReduceValid                     (_laneVec_4_maskUnitRequest_bits_fpReduceValid),
    .exeReq_5_valid                                  (_laneVec_5_maskUnitRequest_valid & ~_laneVec_5_maskRequestToLSU),
    .exeReq_5_bits_source1                           (_laneVec_5_maskUnitRequest_bits_source1),
    .exeReq_5_bits_source2                           (_laneVec_5_maskUnitRequest_bits_source2),
    .exeReq_5_bits_index                             (_laneVec_5_maskUnitRequest_bits_index),
    .exeReq_5_bits_ffo                               (_laneVec_5_maskUnitRequest_bits_ffo),
    .exeReq_5_bits_fpReduceValid                     (_laneVec_5_maskUnitRequest_bits_fpReduceValid),
    .exeReq_6_valid                                  (_laneVec_6_maskUnitRequest_valid & ~_laneVec_6_maskRequestToLSU),
    .exeReq_6_bits_source1                           (_laneVec_6_maskUnitRequest_bits_source1),
    .exeReq_6_bits_source2                           (_laneVec_6_maskUnitRequest_bits_source2),
    .exeReq_6_bits_index                             (_laneVec_6_maskUnitRequest_bits_index),
    .exeReq_6_bits_ffo                               (_laneVec_6_maskUnitRequest_bits_ffo),
    .exeReq_6_bits_fpReduceValid                     (_laneVec_6_maskUnitRequest_bits_fpReduceValid),
    .exeReq_7_valid                                  (_laneVec_7_maskUnitRequest_valid & ~_laneVec_7_maskRequestToLSU),
    .exeReq_7_bits_source1                           (_laneVec_7_maskUnitRequest_bits_source1),
    .exeReq_7_bits_source2                           (_laneVec_7_maskUnitRequest_bits_source2),
    .exeReq_7_bits_index                             (_laneVec_7_maskUnitRequest_bits_index),
    .exeReq_7_bits_ffo                               (_laneVec_7_maskUnitRequest_bits_ffo),
    .exeReq_7_bits_fpReduceValid                     (_laneVec_7_maskUnitRequest_bits_fpReduceValid),
    .exeReq_8_valid                                  (_laneVec_8_maskUnitRequest_valid & ~_laneVec_8_maskRequestToLSU),
    .exeReq_8_bits_source1                           (_laneVec_8_maskUnitRequest_bits_source1),
    .exeReq_8_bits_source2                           (_laneVec_8_maskUnitRequest_bits_source2),
    .exeReq_8_bits_index                             (_laneVec_8_maskUnitRequest_bits_index),
    .exeReq_8_bits_ffo                               (_laneVec_8_maskUnitRequest_bits_ffo),
    .exeReq_8_bits_fpReduceValid                     (_laneVec_8_maskUnitRequest_bits_fpReduceValid),
    .exeReq_9_valid                                  (_laneVec_9_maskUnitRequest_valid & ~_laneVec_9_maskRequestToLSU),
    .exeReq_9_bits_source1                           (_laneVec_9_maskUnitRequest_bits_source1),
    .exeReq_9_bits_source2                           (_laneVec_9_maskUnitRequest_bits_source2),
    .exeReq_9_bits_index                             (_laneVec_9_maskUnitRequest_bits_index),
    .exeReq_9_bits_ffo                               (_laneVec_9_maskUnitRequest_bits_ffo),
    .exeReq_9_bits_fpReduceValid                     (_laneVec_9_maskUnitRequest_bits_fpReduceValid),
    .exeReq_10_valid                                 (_laneVec_10_maskUnitRequest_valid & ~_laneVec_10_maskRequestToLSU),
    .exeReq_10_bits_source1                          (_laneVec_10_maskUnitRequest_bits_source1),
    .exeReq_10_bits_source2                          (_laneVec_10_maskUnitRequest_bits_source2),
    .exeReq_10_bits_index                            (_laneVec_10_maskUnitRequest_bits_index),
    .exeReq_10_bits_ffo                              (_laneVec_10_maskUnitRequest_bits_ffo),
    .exeReq_10_bits_fpReduceValid                    (_laneVec_10_maskUnitRequest_bits_fpReduceValid),
    .exeReq_11_valid                                 (_laneVec_11_maskUnitRequest_valid & ~_laneVec_11_maskRequestToLSU),
    .exeReq_11_bits_source1                          (_laneVec_11_maskUnitRequest_bits_source1),
    .exeReq_11_bits_source2                          (_laneVec_11_maskUnitRequest_bits_source2),
    .exeReq_11_bits_index                            (_laneVec_11_maskUnitRequest_bits_index),
    .exeReq_11_bits_ffo                              (_laneVec_11_maskUnitRequest_bits_ffo),
    .exeReq_11_bits_fpReduceValid                    (_laneVec_11_maskUnitRequest_bits_fpReduceValid),
    .exeReq_12_valid                                 (_laneVec_12_maskUnitRequest_valid & ~_laneVec_12_maskRequestToLSU),
    .exeReq_12_bits_source1                          (_laneVec_12_maskUnitRequest_bits_source1),
    .exeReq_12_bits_source2                          (_laneVec_12_maskUnitRequest_bits_source2),
    .exeReq_12_bits_index                            (_laneVec_12_maskUnitRequest_bits_index),
    .exeReq_12_bits_ffo                              (_laneVec_12_maskUnitRequest_bits_ffo),
    .exeReq_12_bits_fpReduceValid                    (_laneVec_12_maskUnitRequest_bits_fpReduceValid),
    .exeReq_13_valid                                 (_laneVec_13_maskUnitRequest_valid & ~_laneVec_13_maskRequestToLSU),
    .exeReq_13_bits_source1                          (_laneVec_13_maskUnitRequest_bits_source1),
    .exeReq_13_bits_source2                          (_laneVec_13_maskUnitRequest_bits_source2),
    .exeReq_13_bits_index                            (_laneVec_13_maskUnitRequest_bits_index),
    .exeReq_13_bits_ffo                              (_laneVec_13_maskUnitRequest_bits_ffo),
    .exeReq_13_bits_fpReduceValid                    (_laneVec_13_maskUnitRequest_bits_fpReduceValid),
    .exeReq_14_valid                                 (_laneVec_14_maskUnitRequest_valid & ~_laneVec_14_maskRequestToLSU),
    .exeReq_14_bits_source1                          (_laneVec_14_maskUnitRequest_bits_source1),
    .exeReq_14_bits_source2                          (_laneVec_14_maskUnitRequest_bits_source2),
    .exeReq_14_bits_index                            (_laneVec_14_maskUnitRequest_bits_index),
    .exeReq_14_bits_ffo                              (_laneVec_14_maskUnitRequest_bits_ffo),
    .exeReq_14_bits_fpReduceValid                    (_laneVec_14_maskUnitRequest_bits_fpReduceValid),
    .exeReq_15_valid                                 (_laneVec_15_maskUnitRequest_valid & ~_laneVec_15_maskRequestToLSU),
    .exeReq_15_bits_source1                          (_laneVec_15_maskUnitRequest_bits_source1),
    .exeReq_15_bits_source2                          (_laneVec_15_maskUnitRequest_bits_source2),
    .exeReq_15_bits_index                            (_laneVec_15_maskUnitRequest_bits_index),
    .exeReq_15_bits_ffo                              (_laneVec_15_maskUnitRequest_bits_ffo),
    .exeReq_15_bits_fpReduceValid                    (_laneVec_15_maskUnitRequest_bits_fpReduceValid),
    .exeResp_0_ready                                 (x22_0_ready),
    .exeResp_0_valid                                 (_maskUnit_exeResp_0_valid),
    .exeResp_0_bits_vd                               (x22_0_bits_vd),
    .exeResp_0_bits_offset                           (x22_0_bits_offset),
    .exeResp_0_bits_mask                             (_maskUnit_exeResp_0_bits_mask),
    .exeResp_0_bits_data                             (x22_0_bits_data),
    .exeResp_0_bits_instructionIndex                 (_maskUnit_exeResp_0_bits_instructionIndex),
    .exeResp_1_ready                                 (x22_1_0_ready),
    .exeResp_1_valid                                 (_maskUnit_exeResp_1_valid),
    .exeResp_1_bits_vd                               (x22_1_0_bits_vd),
    .exeResp_1_bits_offset                           (x22_1_0_bits_offset),
    .exeResp_1_bits_mask                             (_maskUnit_exeResp_1_bits_mask),
    .exeResp_1_bits_data                             (x22_1_0_bits_data),
    .exeResp_1_bits_instructionIndex                 (_maskUnit_exeResp_1_bits_instructionIndex),
    .exeResp_2_ready                                 (x22_2_0_ready),
    .exeResp_2_valid                                 (_maskUnit_exeResp_2_valid),
    .exeResp_2_bits_vd                               (x22_2_0_bits_vd),
    .exeResp_2_bits_offset                           (x22_2_0_bits_offset),
    .exeResp_2_bits_mask                             (_maskUnit_exeResp_2_bits_mask),
    .exeResp_2_bits_data                             (x22_2_0_bits_data),
    .exeResp_2_bits_instructionIndex                 (_maskUnit_exeResp_2_bits_instructionIndex),
    .exeResp_3_ready                                 (x22_3_0_ready),
    .exeResp_3_valid                                 (_maskUnit_exeResp_3_valid),
    .exeResp_3_bits_vd                               (x22_3_0_bits_vd),
    .exeResp_3_bits_offset                           (x22_3_0_bits_offset),
    .exeResp_3_bits_mask                             (_maskUnit_exeResp_3_bits_mask),
    .exeResp_3_bits_data                             (x22_3_0_bits_data),
    .exeResp_3_bits_instructionIndex                 (_maskUnit_exeResp_3_bits_instructionIndex),
    .exeResp_4_ready                                 (x22_4_0_ready),
    .exeResp_4_valid                                 (_maskUnit_exeResp_4_valid),
    .exeResp_4_bits_vd                               (x22_4_0_bits_vd),
    .exeResp_4_bits_offset                           (x22_4_0_bits_offset),
    .exeResp_4_bits_mask                             (_maskUnit_exeResp_4_bits_mask),
    .exeResp_4_bits_data                             (x22_4_0_bits_data),
    .exeResp_4_bits_instructionIndex                 (_maskUnit_exeResp_4_bits_instructionIndex),
    .exeResp_5_ready                                 (x22_5_0_ready),
    .exeResp_5_valid                                 (_maskUnit_exeResp_5_valid),
    .exeResp_5_bits_vd                               (x22_5_0_bits_vd),
    .exeResp_5_bits_offset                           (x22_5_0_bits_offset),
    .exeResp_5_bits_mask                             (_maskUnit_exeResp_5_bits_mask),
    .exeResp_5_bits_data                             (x22_5_0_bits_data),
    .exeResp_5_bits_instructionIndex                 (_maskUnit_exeResp_5_bits_instructionIndex),
    .exeResp_6_ready                                 (x22_6_0_ready),
    .exeResp_6_valid                                 (_maskUnit_exeResp_6_valid),
    .exeResp_6_bits_vd                               (x22_6_0_bits_vd),
    .exeResp_6_bits_offset                           (x22_6_0_bits_offset),
    .exeResp_6_bits_mask                             (_maskUnit_exeResp_6_bits_mask),
    .exeResp_6_bits_data                             (x22_6_0_bits_data),
    .exeResp_6_bits_instructionIndex                 (_maskUnit_exeResp_6_bits_instructionIndex),
    .exeResp_7_ready                                 (x22_7_0_ready),
    .exeResp_7_valid                                 (_maskUnit_exeResp_7_valid),
    .exeResp_7_bits_vd                               (x22_7_0_bits_vd),
    .exeResp_7_bits_offset                           (x22_7_0_bits_offset),
    .exeResp_7_bits_mask                             (_maskUnit_exeResp_7_bits_mask),
    .exeResp_7_bits_data                             (x22_7_0_bits_data),
    .exeResp_7_bits_instructionIndex                 (_maskUnit_exeResp_7_bits_instructionIndex),
    .exeResp_8_ready                                 (x22_8_0_ready),
    .exeResp_8_valid                                 (_maskUnit_exeResp_8_valid),
    .exeResp_8_bits_vd                               (x22_8_0_bits_vd),
    .exeResp_8_bits_offset                           (x22_8_0_bits_offset),
    .exeResp_8_bits_mask                             (_maskUnit_exeResp_8_bits_mask),
    .exeResp_8_bits_data                             (x22_8_0_bits_data),
    .exeResp_8_bits_instructionIndex                 (_maskUnit_exeResp_8_bits_instructionIndex),
    .exeResp_9_ready                                 (x22_9_0_ready),
    .exeResp_9_valid                                 (_maskUnit_exeResp_9_valid),
    .exeResp_9_bits_vd                               (x22_9_0_bits_vd),
    .exeResp_9_bits_offset                           (x22_9_0_bits_offset),
    .exeResp_9_bits_mask                             (_maskUnit_exeResp_9_bits_mask),
    .exeResp_9_bits_data                             (x22_9_0_bits_data),
    .exeResp_9_bits_instructionIndex                 (_maskUnit_exeResp_9_bits_instructionIndex),
    .exeResp_10_ready                                (x22_10_0_ready),
    .exeResp_10_valid                                (_maskUnit_exeResp_10_valid),
    .exeResp_10_bits_vd                              (x22_10_0_bits_vd),
    .exeResp_10_bits_offset                          (x22_10_0_bits_offset),
    .exeResp_10_bits_mask                            (_maskUnit_exeResp_10_bits_mask),
    .exeResp_10_bits_data                            (x22_10_0_bits_data),
    .exeResp_10_bits_instructionIndex                (_maskUnit_exeResp_10_bits_instructionIndex),
    .exeResp_11_ready                                (x22_11_0_ready),
    .exeResp_11_valid                                (_maskUnit_exeResp_11_valid),
    .exeResp_11_bits_vd                              (x22_11_0_bits_vd),
    .exeResp_11_bits_offset                          (x22_11_0_bits_offset),
    .exeResp_11_bits_mask                            (_maskUnit_exeResp_11_bits_mask),
    .exeResp_11_bits_data                            (x22_11_0_bits_data),
    .exeResp_11_bits_instructionIndex                (_maskUnit_exeResp_11_bits_instructionIndex),
    .exeResp_12_ready                                (x22_12_0_ready),
    .exeResp_12_valid                                (_maskUnit_exeResp_12_valid),
    .exeResp_12_bits_vd                              (x22_12_0_bits_vd),
    .exeResp_12_bits_offset                          (x22_12_0_bits_offset),
    .exeResp_12_bits_mask                            (_maskUnit_exeResp_12_bits_mask),
    .exeResp_12_bits_data                            (x22_12_0_bits_data),
    .exeResp_12_bits_instructionIndex                (_maskUnit_exeResp_12_bits_instructionIndex),
    .exeResp_13_ready                                (x22_13_0_ready),
    .exeResp_13_valid                                (_maskUnit_exeResp_13_valid),
    .exeResp_13_bits_vd                              (x22_13_0_bits_vd),
    .exeResp_13_bits_offset                          (x22_13_0_bits_offset),
    .exeResp_13_bits_mask                            (_maskUnit_exeResp_13_bits_mask),
    .exeResp_13_bits_data                            (x22_13_0_bits_data),
    .exeResp_13_bits_instructionIndex                (_maskUnit_exeResp_13_bits_instructionIndex),
    .exeResp_14_ready                                (x22_14_0_ready),
    .exeResp_14_valid                                (_maskUnit_exeResp_14_valid),
    .exeResp_14_bits_vd                              (x22_14_0_bits_vd),
    .exeResp_14_bits_offset                          (x22_14_0_bits_offset),
    .exeResp_14_bits_mask                            (_maskUnit_exeResp_14_bits_mask),
    .exeResp_14_bits_data                            (x22_14_0_bits_data),
    .exeResp_14_bits_instructionIndex                (_maskUnit_exeResp_14_bits_instructionIndex),
    .exeResp_15_ready                                (x22_15_0_ready),
    .exeResp_15_valid                                (_maskUnit_exeResp_15_valid),
    .exeResp_15_bits_vd                              (x22_15_0_bits_vd),
    .exeResp_15_bits_offset                          (x22_15_0_bits_offset),
    .exeResp_15_bits_mask                            (_maskUnit_exeResp_15_bits_mask),
    .exeResp_15_bits_data                            (x22_15_0_bits_data),
    .exeResp_15_bits_instructionIndex                (_maskUnit_exeResp_15_bits_instructionIndex),
    .writeRelease_0                                  (view__writeRelease_0_pipe_out_valid),
    .writeRelease_1                                  (view__writeRelease_1_pipe_out_valid),
    .writeRelease_2                                  (view__writeRelease_2_pipe_out_valid),
    .writeRelease_3                                  (view__writeRelease_3_pipe_out_valid),
    .writeRelease_4                                  (view__writeRelease_4_pipe_out_valid),
    .writeRelease_5                                  (view__writeRelease_5_pipe_out_valid),
    .writeRelease_6                                  (view__writeRelease_6_pipe_out_valid),
    .writeRelease_7                                  (view__writeRelease_7_pipe_out_valid),
    .writeRelease_8                                  (view__writeRelease_8_pipe_out_valid),
    .writeRelease_9                                  (view__writeRelease_9_pipe_out_valid),
    .writeRelease_10                                 (view__writeRelease_10_pipe_out_valid),
    .writeRelease_11                                 (view__writeRelease_11_pipe_out_valid),
    .writeRelease_12                                 (view__writeRelease_12_pipe_out_valid),
    .writeRelease_13                                 (view__writeRelease_13_pipe_out_valid),
    .writeRelease_14                                 (view__writeRelease_14_pipe_out_valid),
    .writeRelease_15                                 (view__writeRelease_15_pipe_out_valid),
    .tokenIO_0_maskRequestRelease                    (_maskUnit_tokenIO_0_maskRequestRelease),
    .tokenIO_1_maskRequestRelease                    (_maskUnit_tokenIO_1_maskRequestRelease),
    .tokenIO_2_maskRequestRelease                    (_maskUnit_tokenIO_2_maskRequestRelease),
    .tokenIO_3_maskRequestRelease                    (_maskUnit_tokenIO_3_maskRequestRelease),
    .tokenIO_4_maskRequestRelease                    (_maskUnit_tokenIO_4_maskRequestRelease),
    .tokenIO_5_maskRequestRelease                    (_maskUnit_tokenIO_5_maskRequestRelease),
    .tokenIO_6_maskRequestRelease                    (_maskUnit_tokenIO_6_maskRequestRelease),
    .tokenIO_7_maskRequestRelease                    (_maskUnit_tokenIO_7_maskRequestRelease),
    .tokenIO_8_maskRequestRelease                    (_maskUnit_tokenIO_8_maskRequestRelease),
    .tokenIO_9_maskRequestRelease                    (_maskUnit_tokenIO_9_maskRequestRelease),
    .tokenIO_10_maskRequestRelease                   (_maskUnit_tokenIO_10_maskRequestRelease),
    .tokenIO_11_maskRequestRelease                   (_maskUnit_tokenIO_11_maskRequestRelease),
    .tokenIO_12_maskRequestRelease                   (_maskUnit_tokenIO_12_maskRequestRelease),
    .tokenIO_13_maskRequestRelease                   (_maskUnit_tokenIO_13_maskRequestRelease),
    .tokenIO_14_maskRequestRelease                   (_maskUnit_tokenIO_14_maskRequestRelease),
    .tokenIO_15_maskRequestRelease                   (_maskUnit_tokenIO_15_maskRequestRelease),
    .readChannel_0_ready                             (x13_0_ready),
    .readChannel_0_valid                             (x13_0_valid),
    .readChannel_0_bits_vs                           (x13_0_bits_vs),
    .readChannel_0_bits_offset                       (x13_0_bits_offset),
    .readChannel_0_bits_instructionIndex             (x13_0_bits_instructionIndex),
    .readChannel_1_ready                             (x13_1_0_ready),
    .readChannel_1_valid                             (x13_1_0_valid),
    .readChannel_1_bits_vs                           (x13_1_0_bits_vs),
    .readChannel_1_bits_offset                       (x13_1_0_bits_offset),
    .readChannel_1_bits_instructionIndex             (x13_1_0_bits_instructionIndex),
    .readChannel_2_ready                             (x13_2_0_ready),
    .readChannel_2_valid                             (x13_2_0_valid),
    .readChannel_2_bits_vs                           (x13_2_0_bits_vs),
    .readChannel_2_bits_offset                       (x13_2_0_bits_offset),
    .readChannel_2_bits_instructionIndex             (x13_2_0_bits_instructionIndex),
    .readChannel_3_ready                             (x13_3_0_ready),
    .readChannel_3_valid                             (x13_3_0_valid),
    .readChannel_3_bits_vs                           (x13_3_0_bits_vs),
    .readChannel_3_bits_offset                       (x13_3_0_bits_offset),
    .readChannel_3_bits_instructionIndex             (x13_3_0_bits_instructionIndex),
    .readChannel_4_ready                             (x13_4_0_ready),
    .readChannel_4_valid                             (x13_4_0_valid),
    .readChannel_4_bits_vs                           (x13_4_0_bits_vs),
    .readChannel_4_bits_offset                       (x13_4_0_bits_offset),
    .readChannel_4_bits_instructionIndex             (x13_4_0_bits_instructionIndex),
    .readChannel_5_ready                             (x13_5_0_ready),
    .readChannel_5_valid                             (x13_5_0_valid),
    .readChannel_5_bits_vs                           (x13_5_0_bits_vs),
    .readChannel_5_bits_offset                       (x13_5_0_bits_offset),
    .readChannel_5_bits_instructionIndex             (x13_5_0_bits_instructionIndex),
    .readChannel_6_ready                             (x13_6_0_ready),
    .readChannel_6_valid                             (x13_6_0_valid),
    .readChannel_6_bits_vs                           (x13_6_0_bits_vs),
    .readChannel_6_bits_offset                       (x13_6_0_bits_offset),
    .readChannel_6_bits_instructionIndex             (x13_6_0_bits_instructionIndex),
    .readChannel_7_ready                             (x13_7_0_ready),
    .readChannel_7_valid                             (x13_7_0_valid),
    .readChannel_7_bits_vs                           (x13_7_0_bits_vs),
    .readChannel_7_bits_offset                       (x13_7_0_bits_offset),
    .readChannel_7_bits_instructionIndex             (x13_7_0_bits_instructionIndex),
    .readChannel_8_ready                             (x13_8_0_ready),
    .readChannel_8_valid                             (x13_8_0_valid),
    .readChannel_8_bits_vs                           (x13_8_0_bits_vs),
    .readChannel_8_bits_offset                       (x13_8_0_bits_offset),
    .readChannel_8_bits_instructionIndex             (x13_8_0_bits_instructionIndex),
    .readChannel_9_ready                             (x13_9_0_ready),
    .readChannel_9_valid                             (x13_9_0_valid),
    .readChannel_9_bits_vs                           (x13_9_0_bits_vs),
    .readChannel_9_bits_offset                       (x13_9_0_bits_offset),
    .readChannel_9_bits_instructionIndex             (x13_9_0_bits_instructionIndex),
    .readChannel_10_ready                            (x13_10_0_ready),
    .readChannel_10_valid                            (x13_10_0_valid),
    .readChannel_10_bits_vs                          (x13_10_0_bits_vs),
    .readChannel_10_bits_offset                      (x13_10_0_bits_offset),
    .readChannel_10_bits_instructionIndex            (x13_10_0_bits_instructionIndex),
    .readChannel_11_ready                            (x13_11_0_ready),
    .readChannel_11_valid                            (x13_11_0_valid),
    .readChannel_11_bits_vs                          (x13_11_0_bits_vs),
    .readChannel_11_bits_offset                      (x13_11_0_bits_offset),
    .readChannel_11_bits_instructionIndex            (x13_11_0_bits_instructionIndex),
    .readChannel_12_ready                            (x13_12_0_ready),
    .readChannel_12_valid                            (x13_12_0_valid),
    .readChannel_12_bits_vs                          (x13_12_0_bits_vs),
    .readChannel_12_bits_offset                      (x13_12_0_bits_offset),
    .readChannel_12_bits_instructionIndex            (x13_12_0_bits_instructionIndex),
    .readChannel_13_ready                            (x13_13_0_ready),
    .readChannel_13_valid                            (x13_13_0_valid),
    .readChannel_13_bits_vs                          (x13_13_0_bits_vs),
    .readChannel_13_bits_offset                      (x13_13_0_bits_offset),
    .readChannel_13_bits_instructionIndex            (x13_13_0_bits_instructionIndex),
    .readChannel_14_ready                            (x13_14_0_ready),
    .readChannel_14_valid                            (x13_14_0_valid),
    .readChannel_14_bits_vs                          (x13_14_0_bits_vs),
    .readChannel_14_bits_offset                      (x13_14_0_bits_offset),
    .readChannel_14_bits_instructionIndex            (x13_14_0_bits_instructionIndex),
    .readChannel_15_ready                            (x13_15_0_ready),
    .readChannel_15_valid                            (x13_15_0_valid),
    .readChannel_15_bits_vs                          (x13_15_0_bits_vs),
    .readChannel_15_bits_offset                      (x13_15_0_bits_offset),
    .readChannel_15_bits_instructionIndex            (x13_15_0_bits_instructionIndex),
    .readResult_0_valid                              (shifterReg_16_0_valid),
    .readResult_0_bits                               (shifterReg_16_0_bits),
    .readResult_1_valid                              (shifterReg_18_0_valid),
    .readResult_1_bits                               (shifterReg_18_0_bits),
    .readResult_2_valid                              (shifterReg_20_0_valid),
    .readResult_2_bits                               (shifterReg_20_0_bits),
    .readResult_3_valid                              (shifterReg_22_0_valid),
    .readResult_3_bits                               (shifterReg_22_0_bits),
    .readResult_4_valid                              (shifterReg_24_0_valid),
    .readResult_4_bits                               (shifterReg_24_0_bits),
    .readResult_5_valid                              (shifterReg_26_0_valid),
    .readResult_5_bits                               (shifterReg_26_0_bits),
    .readResult_6_valid                              (shifterReg_28_0_valid),
    .readResult_6_bits                               (shifterReg_28_0_bits),
    .readResult_7_valid                              (shifterReg_30_0_valid),
    .readResult_7_bits                               (shifterReg_30_0_bits),
    .readResult_8_valid                              (shifterReg_32_0_valid),
    .readResult_8_bits                               (shifterReg_32_0_bits),
    .readResult_9_valid                              (shifterReg_34_0_valid),
    .readResult_9_bits                               (shifterReg_34_0_bits),
    .readResult_10_valid                             (shifterReg_36_0_valid),
    .readResult_10_bits                              (shifterReg_36_0_bits),
    .readResult_11_valid                             (shifterReg_38_0_valid),
    .readResult_11_bits                              (shifterReg_38_0_bits),
    .readResult_12_valid                             (shifterReg_40_0_valid),
    .readResult_12_bits                              (shifterReg_40_0_bits),
    .readResult_13_valid                             (shifterReg_42_0_valid),
    .readResult_13_bits                              (shifterReg_42_0_bits),
    .readResult_14_valid                             (shifterReg_44_0_valid),
    .readResult_14_bits                              (shifterReg_44_0_bits),
    .readResult_15_valid                             (shifterReg_46_0_valid),
    .readResult_15_bits                              (shifterReg_46_0_bits),
    .lastReport                                      (_maskUnit_lastReport),
    .laneMaskInput_0                                 (_maskUnit_laneMaskInput_0),
    .laneMaskInput_1                                 (_maskUnit_laneMaskInput_1),
    .laneMaskInput_2                                 (_maskUnit_laneMaskInput_2),
    .laneMaskInput_3                                 (_maskUnit_laneMaskInput_3),
    .laneMaskInput_4                                 (_maskUnit_laneMaskInput_4),
    .laneMaskInput_5                                 (_maskUnit_laneMaskInput_5),
    .laneMaskInput_6                                 (_maskUnit_laneMaskInput_6),
    .laneMaskInput_7                                 (_maskUnit_laneMaskInput_7),
    .laneMaskInput_8                                 (_maskUnit_laneMaskInput_8),
    .laneMaskInput_9                                 (_maskUnit_laneMaskInput_9),
    .laneMaskInput_10                                (_maskUnit_laneMaskInput_10),
    .laneMaskInput_11                                (_maskUnit_laneMaskInput_11),
    .laneMaskInput_12                                (_maskUnit_laneMaskInput_12),
    .laneMaskInput_13                                (_maskUnit_laneMaskInput_13),
    .laneMaskInput_14                                (_maskUnit_laneMaskInput_14),
    .laneMaskInput_15                                (_maskUnit_laneMaskInput_15),
    .laneMaskSelect_0                                (view__laneMaskSelect_0_pipe_pipe_out_bits),
    .laneMaskSelect_1                                (view__laneMaskSelect_1_pipe_pipe_out_bits),
    .laneMaskSelect_2                                (view__laneMaskSelect_2_pipe_pipe_out_bits),
    .laneMaskSelect_3                                (view__laneMaskSelect_3_pipe_pipe_out_bits),
    .laneMaskSelect_4                                (view__laneMaskSelect_4_pipe_pipe_out_bits),
    .laneMaskSelect_5                                (view__laneMaskSelect_5_pipe_pipe_out_bits),
    .laneMaskSelect_6                                (view__laneMaskSelect_6_pipe_pipe_out_bits),
    .laneMaskSelect_7                                (view__laneMaskSelect_7_pipe_pipe_out_bits),
    .laneMaskSelect_8                                (view__laneMaskSelect_8_pipe_pipe_out_bits),
    .laneMaskSelect_9                                (view__laneMaskSelect_9_pipe_pipe_out_bits),
    .laneMaskSelect_10                               (view__laneMaskSelect_10_pipe_pipe_out_bits),
    .laneMaskSelect_11                               (view__laneMaskSelect_11_pipe_pipe_out_bits),
    .laneMaskSelect_12                               (view__laneMaskSelect_12_pipe_pipe_out_bits),
    .laneMaskSelect_13                               (view__laneMaskSelect_13_pipe_pipe_out_bits),
    .laneMaskSelect_14                               (view__laneMaskSelect_14_pipe_pipe_out_bits),
    .laneMaskSelect_15                               (view__laneMaskSelect_15_pipe_pipe_out_bits),
    .laneMaskSewSelect_0                             (view__laneMaskSewSelect_0_pipe_pipe_out_bits),
    .laneMaskSewSelect_1                             (view__laneMaskSewSelect_1_pipe_pipe_out_bits),
    .laneMaskSewSelect_2                             (view__laneMaskSewSelect_2_pipe_pipe_out_bits),
    .laneMaskSewSelect_3                             (view__laneMaskSewSelect_3_pipe_pipe_out_bits),
    .laneMaskSewSelect_4                             (view__laneMaskSewSelect_4_pipe_pipe_out_bits),
    .laneMaskSewSelect_5                             (view__laneMaskSewSelect_5_pipe_pipe_out_bits),
    .laneMaskSewSelect_6                             (view__laneMaskSewSelect_6_pipe_pipe_out_bits),
    .laneMaskSewSelect_7                             (view__laneMaskSewSelect_7_pipe_pipe_out_bits),
    .laneMaskSewSelect_8                             (view__laneMaskSewSelect_8_pipe_pipe_out_bits),
    .laneMaskSewSelect_9                             (view__laneMaskSewSelect_9_pipe_pipe_out_bits),
    .laneMaskSewSelect_10                            (view__laneMaskSewSelect_10_pipe_pipe_out_bits),
    .laneMaskSewSelect_11                            (view__laneMaskSewSelect_11_pipe_pipe_out_bits),
    .laneMaskSewSelect_12                            (view__laneMaskSewSelect_12_pipe_pipe_out_bits),
    .laneMaskSewSelect_13                            (view__laneMaskSewSelect_13_pipe_pipe_out_bits),
    .laneMaskSewSelect_14                            (view__laneMaskSewSelect_14_pipe_pipe_out_bits),
    .laneMaskSewSelect_15                            (view__laneMaskSewSelect_15_pipe_pipe_out_bits),
    .v0UpdateVec_0_valid                             (_laneVec_0_v0Update_valid),
    .v0UpdateVec_0_bits_data                         (_laneVec_0_v0Update_bits_data),
    .v0UpdateVec_0_bits_offset                       (_laneVec_0_v0Update_bits_offset),
    .v0UpdateVec_0_bits_mask                         (_laneVec_0_v0Update_bits_mask),
    .v0UpdateVec_1_valid                             (_laneVec_1_v0Update_valid),
    .v0UpdateVec_1_bits_data                         (_laneVec_1_v0Update_bits_data),
    .v0UpdateVec_1_bits_offset                       (_laneVec_1_v0Update_bits_offset),
    .v0UpdateVec_1_bits_mask                         (_laneVec_1_v0Update_bits_mask),
    .v0UpdateVec_2_valid                             (_laneVec_2_v0Update_valid),
    .v0UpdateVec_2_bits_data                         (_laneVec_2_v0Update_bits_data),
    .v0UpdateVec_2_bits_offset                       (_laneVec_2_v0Update_bits_offset),
    .v0UpdateVec_2_bits_mask                         (_laneVec_2_v0Update_bits_mask),
    .v0UpdateVec_3_valid                             (_laneVec_3_v0Update_valid),
    .v0UpdateVec_3_bits_data                         (_laneVec_3_v0Update_bits_data),
    .v0UpdateVec_3_bits_offset                       (_laneVec_3_v0Update_bits_offset),
    .v0UpdateVec_3_bits_mask                         (_laneVec_3_v0Update_bits_mask),
    .v0UpdateVec_4_valid                             (_laneVec_4_v0Update_valid),
    .v0UpdateVec_4_bits_data                         (_laneVec_4_v0Update_bits_data),
    .v0UpdateVec_4_bits_offset                       (_laneVec_4_v0Update_bits_offset),
    .v0UpdateVec_4_bits_mask                         (_laneVec_4_v0Update_bits_mask),
    .v0UpdateVec_5_valid                             (_laneVec_5_v0Update_valid),
    .v0UpdateVec_5_bits_data                         (_laneVec_5_v0Update_bits_data),
    .v0UpdateVec_5_bits_offset                       (_laneVec_5_v0Update_bits_offset),
    .v0UpdateVec_5_bits_mask                         (_laneVec_5_v0Update_bits_mask),
    .v0UpdateVec_6_valid                             (_laneVec_6_v0Update_valid),
    .v0UpdateVec_6_bits_data                         (_laneVec_6_v0Update_bits_data),
    .v0UpdateVec_6_bits_offset                       (_laneVec_6_v0Update_bits_offset),
    .v0UpdateVec_6_bits_mask                         (_laneVec_6_v0Update_bits_mask),
    .v0UpdateVec_7_valid                             (_laneVec_7_v0Update_valid),
    .v0UpdateVec_7_bits_data                         (_laneVec_7_v0Update_bits_data),
    .v0UpdateVec_7_bits_offset                       (_laneVec_7_v0Update_bits_offset),
    .v0UpdateVec_7_bits_mask                         (_laneVec_7_v0Update_bits_mask),
    .v0UpdateVec_8_valid                             (_laneVec_8_v0Update_valid),
    .v0UpdateVec_8_bits_data                         (_laneVec_8_v0Update_bits_data),
    .v0UpdateVec_8_bits_offset                       (_laneVec_8_v0Update_bits_offset),
    .v0UpdateVec_8_bits_mask                         (_laneVec_8_v0Update_bits_mask),
    .v0UpdateVec_9_valid                             (_laneVec_9_v0Update_valid),
    .v0UpdateVec_9_bits_data                         (_laneVec_9_v0Update_bits_data),
    .v0UpdateVec_9_bits_offset                       (_laneVec_9_v0Update_bits_offset),
    .v0UpdateVec_9_bits_mask                         (_laneVec_9_v0Update_bits_mask),
    .v0UpdateVec_10_valid                            (_laneVec_10_v0Update_valid),
    .v0UpdateVec_10_bits_data                        (_laneVec_10_v0Update_bits_data),
    .v0UpdateVec_10_bits_offset                      (_laneVec_10_v0Update_bits_offset),
    .v0UpdateVec_10_bits_mask                        (_laneVec_10_v0Update_bits_mask),
    .v0UpdateVec_11_valid                            (_laneVec_11_v0Update_valid),
    .v0UpdateVec_11_bits_data                        (_laneVec_11_v0Update_bits_data),
    .v0UpdateVec_11_bits_offset                      (_laneVec_11_v0Update_bits_offset),
    .v0UpdateVec_11_bits_mask                        (_laneVec_11_v0Update_bits_mask),
    .v0UpdateVec_12_valid                            (_laneVec_12_v0Update_valid),
    .v0UpdateVec_12_bits_data                        (_laneVec_12_v0Update_bits_data),
    .v0UpdateVec_12_bits_offset                      (_laneVec_12_v0Update_bits_offset),
    .v0UpdateVec_12_bits_mask                        (_laneVec_12_v0Update_bits_mask),
    .v0UpdateVec_13_valid                            (_laneVec_13_v0Update_valid),
    .v0UpdateVec_13_bits_data                        (_laneVec_13_v0Update_bits_data),
    .v0UpdateVec_13_bits_offset                      (_laneVec_13_v0Update_bits_offset),
    .v0UpdateVec_13_bits_mask                        (_laneVec_13_v0Update_bits_mask),
    .v0UpdateVec_14_valid                            (_laneVec_14_v0Update_valid),
    .v0UpdateVec_14_bits_data                        (_laneVec_14_v0Update_bits_data),
    .v0UpdateVec_14_bits_offset                      (_laneVec_14_v0Update_bits_offset),
    .v0UpdateVec_14_bits_mask                        (_laneVec_14_v0Update_bits_mask),
    .v0UpdateVec_15_valid                            (_laneVec_15_v0Update_valid),
    .v0UpdateVec_15_bits_data                        (_laneVec_15_v0Update_bits_data),
    .v0UpdateVec_15_bits_offset                      (_laneVec_15_v0Update_bits_offset),
    .v0UpdateVec_15_bits_mask                        (_laneVec_15_v0Update_bits_mask),
    .writeRDData                                     (retire_rd_bits_rdData_0),
    .gatherData_ready                                (maskUnit_gatherData_ready),
    .gatherData_valid                                (_maskUnit_gatherData_valid),
    .gatherData_bits                                 (_maskUnit_gatherData_bits),
    .gatherRead                                      (gatherNeedRead)
  );
  T1TokenManager tokenManager (
    .clock                                  (clock),
    .reset                                  (reset),
    .instructionIssue_valid                 (maskUnit_gatherData_ready),
    .instructionIssue_bits_instructionIndex (requestReg_bits_instructionIndex),
    .instructionIssue_bits_writeV0          (~requestReg_bits_decodeResult_targetRd & ~isStoreType & requestReg_bits_vdIsV0),
    .instructionIssue_bits_useV0AsMask      (maskType),
    .instructionIssue_bits_toLane           (~noOffsetReadLoadStore & ~maskUnitInstruction),
    .instructionIssue_bits_toMask           (requestReg_bits_decodeResult_maskUnit),
    .lsuWriteV0_0_valid                     (x22_1_ready & _lsu_vrfWritePort_0_valid & _lsu_vrfWritePort_0_bits_vd == 5'h0 & (|_lsu_vrfWritePort_0_bits_mask)),
    .lsuWriteV0_0_bits                      (_lsu_vrfWritePort_0_bits_instructionIndex),
    .lsuWriteV0_1_valid                     (x22_1_1_ready & _lsu_vrfWritePort_1_valid & _lsu_vrfWritePort_1_bits_vd == 5'h0 & (|_lsu_vrfWritePort_1_bits_mask)),
    .lsuWriteV0_1_bits                      (_lsu_vrfWritePort_1_bits_instructionIndex),
    .lsuWriteV0_2_valid                     (x22_2_1_ready & _lsu_vrfWritePort_2_valid & _lsu_vrfWritePort_2_bits_vd == 5'h0 & (|_lsu_vrfWritePort_2_bits_mask)),
    .lsuWriteV0_2_bits                      (_lsu_vrfWritePort_2_bits_instructionIndex),
    .lsuWriteV0_3_valid                     (x22_3_1_ready & _lsu_vrfWritePort_3_valid & _lsu_vrfWritePort_3_bits_vd == 5'h0 & (|_lsu_vrfWritePort_3_bits_mask)),
    .lsuWriteV0_3_bits                      (_lsu_vrfWritePort_3_bits_instructionIndex),
    .lsuWriteV0_4_valid                     (x22_4_1_ready & _lsu_vrfWritePort_4_valid & _lsu_vrfWritePort_4_bits_vd == 5'h0 & (|_lsu_vrfWritePort_4_bits_mask)),
    .lsuWriteV0_4_bits                      (_lsu_vrfWritePort_4_bits_instructionIndex),
    .lsuWriteV0_5_valid                     (x22_5_1_ready & _lsu_vrfWritePort_5_valid & _lsu_vrfWritePort_5_bits_vd == 5'h0 & (|_lsu_vrfWritePort_5_bits_mask)),
    .lsuWriteV0_5_bits                      (_lsu_vrfWritePort_5_bits_instructionIndex),
    .lsuWriteV0_6_valid                     (x22_6_1_ready & _lsu_vrfWritePort_6_valid & _lsu_vrfWritePort_6_bits_vd == 5'h0 & (|_lsu_vrfWritePort_6_bits_mask)),
    .lsuWriteV0_6_bits                      (_lsu_vrfWritePort_6_bits_instructionIndex),
    .lsuWriteV0_7_valid                     (x22_7_1_ready & _lsu_vrfWritePort_7_valid & _lsu_vrfWritePort_7_bits_vd == 5'h0 & (|_lsu_vrfWritePort_7_bits_mask)),
    .lsuWriteV0_7_bits                      (_lsu_vrfWritePort_7_bits_instructionIndex),
    .lsuWriteV0_8_valid                     (x22_8_1_ready & _lsu_vrfWritePort_8_valid & _lsu_vrfWritePort_8_bits_vd == 5'h0 & (|_lsu_vrfWritePort_8_bits_mask)),
    .lsuWriteV0_8_bits                      (_lsu_vrfWritePort_8_bits_instructionIndex),
    .lsuWriteV0_9_valid                     (x22_9_1_ready & _lsu_vrfWritePort_9_valid & _lsu_vrfWritePort_9_bits_vd == 5'h0 & (|_lsu_vrfWritePort_9_bits_mask)),
    .lsuWriteV0_9_bits                      (_lsu_vrfWritePort_9_bits_instructionIndex),
    .lsuWriteV0_10_valid                    (x22_10_1_ready & _lsu_vrfWritePort_10_valid & _lsu_vrfWritePort_10_bits_vd == 5'h0 & (|_lsu_vrfWritePort_10_bits_mask)),
    .lsuWriteV0_10_bits                     (_lsu_vrfWritePort_10_bits_instructionIndex),
    .lsuWriteV0_11_valid                    (x22_11_1_ready & _lsu_vrfWritePort_11_valid & _lsu_vrfWritePort_11_bits_vd == 5'h0 & (|_lsu_vrfWritePort_11_bits_mask)),
    .lsuWriteV0_11_bits                     (_lsu_vrfWritePort_11_bits_instructionIndex),
    .lsuWriteV0_12_valid                    (x22_12_1_ready & _lsu_vrfWritePort_12_valid & _lsu_vrfWritePort_12_bits_vd == 5'h0 & (|_lsu_vrfWritePort_12_bits_mask)),
    .lsuWriteV0_12_bits                     (_lsu_vrfWritePort_12_bits_instructionIndex),
    .lsuWriteV0_13_valid                    (x22_13_1_ready & _lsu_vrfWritePort_13_valid & _lsu_vrfWritePort_13_bits_vd == 5'h0 & (|_lsu_vrfWritePort_13_bits_mask)),
    .lsuWriteV0_13_bits                     (_lsu_vrfWritePort_13_bits_instructionIndex),
    .lsuWriteV0_14_valid                    (x22_14_1_ready & _lsu_vrfWritePort_14_valid & _lsu_vrfWritePort_14_bits_vd == 5'h0 & (|_lsu_vrfWritePort_14_bits_mask)),
    .lsuWriteV0_14_bits                     (_lsu_vrfWritePort_14_bits_instructionIndex),
    .lsuWriteV0_15_valid                    (x22_15_1_ready & _lsu_vrfWritePort_15_valid & _lsu_vrfWritePort_15_bits_vd == 5'h0 & (|_lsu_vrfWritePort_15_bits_mask)),
    .lsuWriteV0_15_bits                     (_lsu_vrfWritePort_15_bits_instructionIndex),
    .issueAllow                             (_tokenManager_issueAllow),
    .instructionFinish_0                    (instructionFinishedPipe_pipe_out_bits),
    .instructionFinish_1                    (instructionFinishedPipe_pipe_out_1_bits),
    .instructionFinish_2                    (instructionFinishedPipe_pipe_out_2_bits),
    .instructionFinish_3                    (instructionFinishedPipe_pipe_out_3_bits),
    .instructionFinish_4                    (instructionFinishedPipe_pipe_out_4_bits),
    .instructionFinish_5                    (instructionFinishedPipe_pipe_out_5_bits),
    .instructionFinish_6                    (instructionFinishedPipe_pipe_out_6_bits),
    .instructionFinish_7                    (instructionFinishedPipe_pipe_out_7_bits),
    .instructionFinish_8                    (instructionFinishedPipe_pipe_out_8_bits),
    .instructionFinish_9                    (instructionFinishedPipe_pipe_out_9_bits),
    .instructionFinish_10                   (instructionFinishedPipe_pipe_out_10_bits),
    .instructionFinish_11                   (instructionFinishedPipe_pipe_out_11_bits),
    .instructionFinish_12                   (instructionFinishedPipe_pipe_out_12_bits),
    .instructionFinish_13                   (instructionFinishedPipe_pipe_out_13_bits),
    .instructionFinish_14                   (instructionFinishedPipe_pipe_out_14_bits),
    .instructionFinish_15                   (instructionFinishedPipe_pipe_out_15_bits),
    .v0WriteValid                           (_tokenManager_v0WriteValid),
    .maskUnitFree                           (slots_3_state_idle)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_enq_ready & queue_enq_valid & ~(_queue_fifo_empty & queue_deq_ready))),
    .pop_req_n    (~(queue_deq_ready & ~_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn),
    .empty        (_queue_fifo_empty),
    .almost_empty (queue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_almostFull),
    .full         (_queue_fifo_full),
    .error        (_queue_fifo_error),
    .data_out     (_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_1_enq_ready & queue_1_enq_valid & ~(_queue_fifo_1_empty & queue_1_deq_ready))),
    .pop_req_n    (~(queue_1_deq_ready & ~_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_1),
    .empty        (_queue_fifo_1_empty),
    .almost_empty (queue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_1_almostFull),
    .full         (_queue_fifo_1_full),
    .error        (_queue_fifo_1_error),
    .data_out     (_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_2_enq_ready & queue_2_enq_valid & ~(_queue_fifo_2_empty & queue_2_deq_ready))),
    .pop_req_n    (~(queue_2_deq_ready & ~_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_2),
    .empty        (_queue_fifo_2_empty),
    .almost_empty (queue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_2_almostFull),
    .full         (_queue_fifo_2_full),
    .error        (_queue_fifo_2_error),
    .data_out     (_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_3_enq_ready & queue_3_enq_valid & ~(_queue_fifo_3_empty & queue_3_deq_ready))),
    .pop_req_n    (~(queue_3_deq_ready & ~_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_3),
    .empty        (_queue_fifo_3_empty),
    .almost_empty (queue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_3_almostFull),
    .full         (_queue_fifo_3_full),
    .error        (_queue_fifo_3_error),
    .data_out     (_queue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_4_enq_ready & queue_4_enq_valid & ~(_queue_fifo_4_empty & queue_4_deq_ready))),
    .pop_req_n    (~(queue_4_deq_ready & ~_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_4),
    .empty        (_queue_fifo_4_empty),
    .almost_empty (queue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_4_almostFull),
    .full         (_queue_fifo_4_full),
    .error        (_queue_fifo_4_error),
    .data_out     (_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_5_enq_ready & queue_5_enq_valid & ~(_queue_fifo_5_empty & queue_5_deq_ready))),
    .pop_req_n    (~(queue_5_deq_ready & ~_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_5),
    .empty        (_queue_fifo_5_empty),
    .almost_empty (queue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_5_almostFull),
    .full         (_queue_fifo_5_full),
    .error        (_queue_fifo_5_error),
    .data_out     (_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_6_enq_ready & queue_6_enq_valid & ~(_queue_fifo_6_empty & queue_6_deq_ready))),
    .pop_req_n    (~(queue_6_deq_ready & ~_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_6),
    .empty        (_queue_fifo_6_empty),
    .almost_empty (queue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_6_almostFull),
    .full         (_queue_fifo_6_full),
    .error        (_queue_fifo_6_error),
    .data_out     (_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_7_enq_ready & queue_7_enq_valid & ~(_queue_fifo_7_empty & queue_7_deq_ready))),
    .pop_req_n    (~(queue_7_deq_ready & ~_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_7),
    .empty        (_queue_fifo_7_empty),
    .almost_empty (queue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_7_almostFull),
    .full         (_queue_fifo_7_full),
    .error        (_queue_fifo_7_error),
    .data_out     (_queue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_8_enq_ready & queue_8_enq_valid & ~(_queue_fifo_8_empty & queue_8_deq_ready))),
    .pop_req_n    (~(queue_8_deq_ready & ~_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_8),
    .empty        (_queue_fifo_8_empty),
    .almost_empty (queue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_8_almostFull),
    .full         (_queue_fifo_8_full),
    .error        (_queue_fifo_8_error),
    .data_out     (_queue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_9_enq_ready & queue_9_enq_valid & ~(_queue_fifo_9_empty & queue_9_deq_ready))),
    .pop_req_n    (~(queue_9_deq_ready & ~_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_9),
    .empty        (_queue_fifo_9_empty),
    .almost_empty (queue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_9_almostFull),
    .full         (_queue_fifo_9_full),
    .error        (_queue_fifo_9_error),
    .data_out     (_queue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_10_enq_ready & queue_10_enq_valid & ~(_queue_fifo_10_empty & queue_10_deq_ready))),
    .pop_req_n    (~(queue_10_deq_ready & ~_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_10),
    .empty        (_queue_fifo_10_empty),
    .almost_empty (queue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_10_almostFull),
    .full         (_queue_fifo_10_full),
    .error        (_queue_fifo_10_error),
    .data_out     (_queue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_11_enq_ready & queue_11_enq_valid & ~(_queue_fifo_11_empty & queue_11_deq_ready))),
    .pop_req_n    (~(queue_11_deq_ready & ~_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_11),
    .empty        (_queue_fifo_11_empty),
    .almost_empty (queue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_11_almostFull),
    .full         (_queue_fifo_11_full),
    .error        (_queue_fifo_11_error),
    .data_out     (_queue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_12_enq_ready & queue_12_enq_valid & ~(_queue_fifo_12_empty & queue_12_deq_ready))),
    .pop_req_n    (~(queue_12_deq_ready & ~_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_12),
    .empty        (_queue_fifo_12_empty),
    .almost_empty (queue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_12_almostFull),
    .full         (_queue_fifo_12_full),
    .error        (_queue_fifo_12_error),
    .data_out     (_queue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_13_enq_ready & queue_13_enq_valid & ~(_queue_fifo_13_empty & queue_13_deq_ready))),
    .pop_req_n    (~(queue_13_deq_ready & ~_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_13),
    .empty        (_queue_fifo_13_empty),
    .almost_empty (queue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_13_almostFull),
    .full         (_queue_fifo_13_full),
    .error        (_queue_fifo_13_error),
    .data_out     (_queue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_14_enq_ready & queue_14_enq_valid & ~(_queue_fifo_14_empty & queue_14_deq_ready))),
    .pop_req_n    (~(queue_14_deq_ready & ~_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_14),
    .empty        (_queue_fifo_14_empty),
    .almost_empty (queue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_14_almostFull),
    .full         (_queue_fifo_14_full),
    .error        (_queue_fifo_14_error),
    .data_out     (_queue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(150)
  ) queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_15_enq_ready & queue_15_enq_valid & ~(_queue_fifo_15_empty & queue_15_deq_ready))),
    .pop_req_n    (~(queue_15_deq_ready & ~_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_15),
    .empty        (_queue_fifo_15_empty),
    .almost_empty (queue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_15_almostFull),
    .full         (_queue_fifo_15_full),
    .error        (_queue_fifo_15_error),
    .data_out     (_queue_fifo_15_data_out)
  );
  Lane laneVec_0 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h0),
    .readBusPort_0_enq_valid                             (shifterReg_48_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_48_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_0_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_0_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_0_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_32_valid),
    .readBusPort_1_enq_valid                             (shifterReg_50_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_50_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_0_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_0_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_0_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_64_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_49_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_49_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_49_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_49_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_49_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_0_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_0_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_0_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_0_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_0_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_0_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_33_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_81_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_81_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_81_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_81_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_81_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_0_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_0_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_0_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_0_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_0_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_0_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_35_valid),
    .laneRequest_ready                                   (_laneVec_0_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_0_valid & laneRequestSinkWire_0_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_0_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_0_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_0_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_0_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_0_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_0_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_0_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_0_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_0_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_0_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_0_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_0_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_0_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_0_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_0_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_0_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_0_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_0_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_0_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_0_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_0_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_0_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_0_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_0_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_0_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_0_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_0_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_0_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_0_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_0_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_0_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_0_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_0_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_0_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_0_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_0_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_0_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_0_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_0_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_0_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_0_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_0_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_0_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_0_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_0_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_0_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_0_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_0_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_0_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_0_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_0_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_0_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_0_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_0_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_0_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_0_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_0_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_0_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_0_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_0_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_0_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_0_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_0_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_0_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_0_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_0_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_0_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_0_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_0_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_0_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_0_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_0_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_0_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_0_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_0_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_0_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[0]),
    .vrfReadAddressChannel_ready                         (sinkWire_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_0_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_1_ready),
    .vrfWriteChannel_valid                               (sinkWire_1_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_1_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_1_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_1_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_1_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_1_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_1_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_0_valid_T),
    .instructionFinished                                 (_laneVec_0_instructionFinished),
    .vxsatReport                                         (_laneVec_0_vxsatReport),
    .v0Update_valid                                      (_laneVec_0_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_0_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_0_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_0_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_bits),
    .maskSelect                                          (_laneVec_0_maskSelect),
    .maskSelectSew                                       (_laneVec_0_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_bits | maskLastPipe_pipe_out_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_0),
    .writeCount                                          (pipe_out_1_bits),
    .writeQueueValid                                     (dataInWritePipeVec_0)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_enq_ready & sinkVec_queue_enq_valid & ~(_sinkVec_queue_fifo_empty & sinkVec_queue_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_deq_ready & ~_sinkVec_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn),
    .empty        (_sinkVec_queue_fifo_empty),
    .almost_empty (sinkVec_queue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_almostFull),
    .full         (_sinkVec_queue_fifo_full),
    .error        (_sinkVec_queue_fifo_error),
    .data_out     (_sinkVec_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_1_enq_ready & sinkVec_queue_1_enq_valid & ~(_sinkVec_queue_fifo_1_empty & sinkVec_queue_1_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_1_deq_ready & ~_sinkVec_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_1),
    .empty        (_sinkVec_queue_fifo_1_empty),
    .almost_empty (sinkVec_queue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_1_almostFull),
    .full         (_sinkVec_queue_fifo_1_full),
    .error        (_sinkVec_queue_fifo_1_error),
    .data_out     (_sinkVec_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_2_enq_ready & sinkVec_queue_2_enq_valid & ~(_sinkVec_queue_fifo_2_empty & sinkVec_queue_2_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_2_deq_ready & ~_sinkVec_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_2),
    .empty        (_sinkVec_queue_fifo_2_empty),
    .almost_empty (sinkVec_queue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_2_almostFull),
    .full         (_sinkVec_queue_fifo_2_full),
    .error        (_sinkVec_queue_fifo_2_error),
    .data_out     (_sinkVec_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_3_enq_ready & sinkVec_queue_3_enq_valid & ~(_sinkVec_queue_fifo_3_empty & sinkVec_queue_3_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_3_deq_ready & ~_sinkVec_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_3),
    .empty        (_sinkVec_queue_fifo_3_empty),
    .almost_empty (sinkVec_queue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_3_almostFull),
    .full         (_sinkVec_queue_fifo_3_full),
    .error        (_sinkVec_queue_fifo_3_error),
    .data_out     (_sinkVec_queue_fifo_3_data_out)
  );
  Lane laneVec_1 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h1),
    .readBusPort_0_enq_valid                             (shifterReg_52_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_52_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_1_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_1_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_1_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_34_valid),
    .readBusPort_1_enq_valid                             (shifterReg_54_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_54_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_1_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_1_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_1_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_66_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_51_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_51_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_51_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_51_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_51_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_1_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_1_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_1_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_1_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_1_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_1_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_37_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_83_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_83_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_83_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_83_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_83_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_1_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_1_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_1_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_1_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_1_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_1_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_39_valid),
    .laneRequest_ready                                   (_laneVec_1_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_1_valid & laneRequestSinkWire_1_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_1_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_1_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_1_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_1_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_1_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_1_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_1_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_1_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_1_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_1_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_1_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_1_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_1_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_1_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_1_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_1_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_1_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_1_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_1_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_1_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_1_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_1_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_1_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_1_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_1_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_1_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_1_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_1_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_1_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_1_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_1_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_1_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_1_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_1_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_1_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_1_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_1_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_1_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_1_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_1_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_1_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_1_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_1_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_1_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_1_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_1_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_1_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_1_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_1_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_1_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_1_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_1_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_1_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_1_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_1_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_1_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_1_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_1_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_1_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_1_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_1_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_1_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_1_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_1_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_1_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_1_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_1_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_1_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_1_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_1_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_1_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_1_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_1_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_1_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_1_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_1_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[1]),
    .vrfReadAddressChannel_ready                         (sinkWire_2_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_2_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_2_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_2_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_2_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_2_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_1_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_3_ready),
    .vrfWriteChannel_valid                               (sinkWire_3_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_3_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_3_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_3_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_3_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_3_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_3_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_1_valid_T),
    .instructionFinished                                 (_laneVec_1_instructionFinished),
    .vxsatReport                                         (_laneVec_1_vxsatReport),
    .v0Update_valid                                      (_laneVec_1_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_1_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_1_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_1_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_1_bits),
    .maskSelect                                          (_laneVec_1_maskSelect),
    .maskSelectSew                                       (_laneVec_1_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_1_bits | maskLastPipe_pipe_out_1_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_1),
    .writeCount                                          (pipe_out_3_bits),
    .writeQueueValid                                     (dataInWritePipeVec_1)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_4_enq_ready & sinkVec_queue_4_enq_valid & ~(_sinkVec_queue_fifo_4_empty & sinkVec_queue_4_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_4_deq_ready & ~_sinkVec_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_4),
    .empty        (_sinkVec_queue_fifo_4_empty),
    .almost_empty (sinkVec_queue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_4_almostFull),
    .full         (_sinkVec_queue_fifo_4_full),
    .error        (_sinkVec_queue_fifo_4_error),
    .data_out     (_sinkVec_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_5_enq_ready & sinkVec_queue_5_enq_valid & ~(_sinkVec_queue_fifo_5_empty & sinkVec_queue_5_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_5_deq_ready & ~_sinkVec_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_5),
    .empty        (_sinkVec_queue_fifo_5_empty),
    .almost_empty (sinkVec_queue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_5_almostFull),
    .full         (_sinkVec_queue_fifo_5_full),
    .error        (_sinkVec_queue_fifo_5_error),
    .data_out     (_sinkVec_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_6_enq_ready & sinkVec_queue_6_enq_valid & ~(_sinkVec_queue_fifo_6_empty & sinkVec_queue_6_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_6_deq_ready & ~_sinkVec_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_6),
    .empty        (_sinkVec_queue_fifo_6_empty),
    .almost_empty (sinkVec_queue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_6_almostFull),
    .full         (_sinkVec_queue_fifo_6_full),
    .error        (_sinkVec_queue_fifo_6_error),
    .data_out     (_sinkVec_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_7_enq_ready & sinkVec_queue_7_enq_valid & ~(_sinkVec_queue_fifo_7_empty & sinkVec_queue_7_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_7_deq_ready & ~_sinkVec_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_7),
    .empty        (_sinkVec_queue_fifo_7_empty),
    .almost_empty (sinkVec_queue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_7_almostFull),
    .full         (_sinkVec_queue_fifo_7_full),
    .error        (_sinkVec_queue_fifo_7_error),
    .data_out     (_sinkVec_queue_fifo_7_data_out)
  );
  Lane laneVec_2 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h2),
    .readBusPort_0_enq_valid                             (shifterReg_56_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_56_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_2_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_2_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_2_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_36_valid),
    .readBusPort_1_enq_valid                             (shifterReg_58_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_58_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_2_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_2_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_2_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_68_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_53_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_53_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_53_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_53_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_53_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_2_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_2_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_2_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_2_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_2_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_2_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_41_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_85_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_85_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_85_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_85_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_85_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_2_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_2_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_2_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_2_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_2_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_2_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_43_valid),
    .laneRequest_ready                                   (_laneVec_2_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_2_valid & laneRequestSinkWire_2_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_2_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_2_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_2_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_2_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_2_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_2_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_2_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_2_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_2_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_2_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_2_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_2_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_2_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_2_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_2_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_2_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_2_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_2_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_2_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_2_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_2_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_2_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_2_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_2_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_2_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_2_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_2_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_2_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_2_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_2_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_2_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_2_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_2_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_2_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_2_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_2_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_2_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_2_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_2_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_2_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_2_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_2_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_2_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_2_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_2_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_2_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_2_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_2_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_2_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_2_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_2_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_2_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_2_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_2_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_2_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_2_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_2_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_2_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_2_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_2_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_2_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_2_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_2_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_2_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_2_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_2_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_2_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_2_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_2_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_2_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_2_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_2_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_2_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_2_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_2_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_2_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[2]),
    .vrfReadAddressChannel_ready                         (sinkWire_4_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_4_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_4_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_4_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_4_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_4_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_2_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_5_ready),
    .vrfWriteChannel_valid                               (sinkWire_5_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_5_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_5_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_5_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_5_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_5_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_5_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_2_valid_T),
    .instructionFinished                                 (_laneVec_2_instructionFinished),
    .vxsatReport                                         (_laneVec_2_vxsatReport),
    .v0Update_valid                                      (_laneVec_2_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_2_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_2_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_2_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_2_bits),
    .maskSelect                                          (_laneVec_2_maskSelect),
    .maskSelectSew                                       (_laneVec_2_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_2_bits | maskLastPipe_pipe_out_2_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_2),
    .writeCount                                          (pipe_out_5_bits),
    .writeQueueValid                                     (dataInWritePipeVec_2)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_8_enq_ready & sinkVec_queue_8_enq_valid & ~(_sinkVec_queue_fifo_8_empty & sinkVec_queue_8_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_8_deq_ready & ~_sinkVec_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_8),
    .empty        (_sinkVec_queue_fifo_8_empty),
    .almost_empty (sinkVec_queue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_8_almostFull),
    .full         (_sinkVec_queue_fifo_8_full),
    .error        (_sinkVec_queue_fifo_8_error),
    .data_out     (_sinkVec_queue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_9_enq_ready & sinkVec_queue_9_enq_valid & ~(_sinkVec_queue_fifo_9_empty & sinkVec_queue_9_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_9_deq_ready & ~_sinkVec_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_9),
    .empty        (_sinkVec_queue_fifo_9_empty),
    .almost_empty (sinkVec_queue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_9_almostFull),
    .full         (_sinkVec_queue_fifo_9_full),
    .error        (_sinkVec_queue_fifo_9_error),
    .data_out     (_sinkVec_queue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_10_enq_ready & sinkVec_queue_10_enq_valid & ~(_sinkVec_queue_fifo_10_empty & sinkVec_queue_10_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_10_deq_ready & ~_sinkVec_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_10),
    .empty        (_sinkVec_queue_fifo_10_empty),
    .almost_empty (sinkVec_queue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_10_almostFull),
    .full         (_sinkVec_queue_fifo_10_full),
    .error        (_sinkVec_queue_fifo_10_error),
    .data_out     (_sinkVec_queue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_11_enq_ready & sinkVec_queue_11_enq_valid & ~(_sinkVec_queue_fifo_11_empty & sinkVec_queue_11_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_11_deq_ready & ~_sinkVec_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_11),
    .empty        (_sinkVec_queue_fifo_11_empty),
    .almost_empty (sinkVec_queue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_11_almostFull),
    .full         (_sinkVec_queue_fifo_11_full),
    .error        (_sinkVec_queue_fifo_11_error),
    .data_out     (_sinkVec_queue_fifo_11_data_out)
  );
  Lane laneVec_3 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h3),
    .readBusPort_0_enq_valid                             (shifterReg_60_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_60_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_3_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_3_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_3_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_38_valid),
    .readBusPort_1_enq_valid                             (shifterReg_62_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_62_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_3_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_3_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_3_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_70_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_55_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_55_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_55_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_55_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_55_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_3_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_3_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_3_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_3_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_3_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_3_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_45_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_87_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_87_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_87_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_87_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_87_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_3_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_3_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_3_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_3_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_3_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_3_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_47_valid),
    .laneRequest_ready                                   (_laneVec_3_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_3_valid & laneRequestSinkWire_3_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_3_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_3_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_3_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_3_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_3_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_3_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_3_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_3_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_3_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_3_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_3_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_3_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_3_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_3_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_3_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_3_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_3_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_3_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_3_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_3_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_3_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_3_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_3_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_3_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_3_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_3_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_3_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_3_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_3_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_3_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_3_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_3_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_3_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_3_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_3_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_3_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_3_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_3_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_3_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_3_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_3_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_3_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_3_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_3_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_3_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_3_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_3_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_3_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_3_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_3_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_3_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_3_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_3_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_3_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_3_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_3_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_3_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_3_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_3_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_3_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_3_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_3_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_3_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_3_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_3_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_3_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_3_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_3_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_3_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_3_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_3_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_3_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_3_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_3_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_3_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_3_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[3]),
    .vrfReadAddressChannel_ready                         (sinkWire_6_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_6_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_6_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_6_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_6_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_6_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_3_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_7_ready),
    .vrfWriteChannel_valid                               (sinkWire_7_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_7_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_7_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_7_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_7_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_7_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_7_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_3_valid_T),
    .instructionFinished                                 (_laneVec_3_instructionFinished),
    .vxsatReport                                         (_laneVec_3_vxsatReport),
    .v0Update_valid                                      (_laneVec_3_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_3_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_3_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_3_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_3_bits),
    .maskSelect                                          (_laneVec_3_maskSelect),
    .maskSelectSew                                       (_laneVec_3_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_3_bits | maskLastPipe_pipe_out_3_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_3),
    .writeCount                                          (pipe_out_7_bits),
    .writeQueueValid                                     (dataInWritePipeVec_3)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_12_enq_ready & sinkVec_queue_12_enq_valid & ~(_sinkVec_queue_fifo_12_empty & sinkVec_queue_12_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_12_deq_ready & ~_sinkVec_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_12),
    .empty        (_sinkVec_queue_fifo_12_empty),
    .almost_empty (sinkVec_queue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_12_almostFull),
    .full         (_sinkVec_queue_fifo_12_full),
    .error        (_sinkVec_queue_fifo_12_error),
    .data_out     (_sinkVec_queue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_13_enq_ready & sinkVec_queue_13_enq_valid & ~(_sinkVec_queue_fifo_13_empty & sinkVec_queue_13_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_13_deq_ready & ~_sinkVec_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_13),
    .empty        (_sinkVec_queue_fifo_13_empty),
    .almost_empty (sinkVec_queue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_13_almostFull),
    .full         (_sinkVec_queue_fifo_13_full),
    .error        (_sinkVec_queue_fifo_13_error),
    .data_out     (_sinkVec_queue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_14_enq_ready & sinkVec_queue_14_enq_valid & ~(_sinkVec_queue_fifo_14_empty & sinkVec_queue_14_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_14_deq_ready & ~_sinkVec_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_14),
    .empty        (_sinkVec_queue_fifo_14_empty),
    .almost_empty (sinkVec_queue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_14_almostFull),
    .full         (_sinkVec_queue_fifo_14_full),
    .error        (_sinkVec_queue_fifo_14_error),
    .data_out     (_sinkVec_queue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_15_enq_ready & sinkVec_queue_15_enq_valid & ~(_sinkVec_queue_fifo_15_empty & sinkVec_queue_15_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_15_deq_ready & ~_sinkVec_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_15),
    .empty        (_sinkVec_queue_fifo_15_empty),
    .almost_empty (sinkVec_queue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_15_almostFull),
    .full         (_sinkVec_queue_fifo_15_full),
    .error        (_sinkVec_queue_fifo_15_error),
    .data_out     (_sinkVec_queue_fifo_15_data_out)
  );
  Lane laneVec_4 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h4),
    .readBusPort_0_enq_valid                             (shifterReg_64_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_64_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_4_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_4_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_4_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_40_valid),
    .readBusPort_1_enq_valid                             (shifterReg_66_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_66_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_4_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_4_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_4_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_72_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_57_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_57_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_57_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_57_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_57_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_4_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_4_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_4_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_4_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_4_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_4_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_49_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_89_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_89_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_89_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_89_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_89_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_4_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_4_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_4_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_4_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_4_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_4_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_51_valid),
    .laneRequest_ready                                   (_laneVec_4_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_4_valid & laneRequestSinkWire_4_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_4_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_4_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_4_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_4_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_4_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_4_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_4_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_4_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_4_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_4_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_4_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_4_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_4_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_4_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_4_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_4_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_4_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_4_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_4_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_4_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_4_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_4_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_4_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_4_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_4_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_4_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_4_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_4_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_4_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_4_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_4_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_4_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_4_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_4_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_4_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_4_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_4_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_4_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_4_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_4_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_4_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_4_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_4_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_4_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_4_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_4_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_4_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_4_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_4_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_4_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_4_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_4_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_4_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_4_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_4_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_4_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_4_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_4_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_4_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_4_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_4_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_4_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_4_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_4_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_4_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_4_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_4_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_4_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_4_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_4_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_4_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_4_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_4_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_4_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_4_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_4_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[4]),
    .vrfReadAddressChannel_ready                         (sinkWire_8_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_8_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_8_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_8_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_8_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_8_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_4_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_9_ready),
    .vrfWriteChannel_valid                               (sinkWire_9_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_9_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_9_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_9_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_9_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_9_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_9_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_4_valid_T),
    .instructionFinished                                 (_laneVec_4_instructionFinished),
    .vxsatReport                                         (_laneVec_4_vxsatReport),
    .v0Update_valid                                      (_laneVec_4_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_4_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_4_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_4_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_4_bits),
    .maskSelect                                          (_laneVec_4_maskSelect),
    .maskSelectSew                                       (_laneVec_4_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_4_bits | maskLastPipe_pipe_out_4_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_4),
    .writeCount                                          (pipe_out_9_bits),
    .writeQueueValid                                     (dataInWritePipeVec_4)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_16_enq_ready & sinkVec_queue_16_enq_valid & ~(_sinkVec_queue_fifo_16_empty & sinkVec_queue_16_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_16_deq_ready & ~_sinkVec_queue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_16),
    .empty        (_sinkVec_queue_fifo_16_empty),
    .almost_empty (sinkVec_queue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_16_almostFull),
    .full         (_sinkVec_queue_fifo_16_full),
    .error        (_sinkVec_queue_fifo_16_error),
    .data_out     (_sinkVec_queue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_17_enq_ready & sinkVec_queue_17_enq_valid & ~(_sinkVec_queue_fifo_17_empty & sinkVec_queue_17_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_17_deq_ready & ~_sinkVec_queue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_17),
    .empty        (_sinkVec_queue_fifo_17_empty),
    .almost_empty (sinkVec_queue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_17_almostFull),
    .full         (_sinkVec_queue_fifo_17_full),
    .error        (_sinkVec_queue_fifo_17_error),
    .data_out     (_sinkVec_queue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_18_enq_ready & sinkVec_queue_18_enq_valid & ~(_sinkVec_queue_fifo_18_empty & sinkVec_queue_18_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_18_deq_ready & ~_sinkVec_queue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_18),
    .empty        (_sinkVec_queue_fifo_18_empty),
    .almost_empty (sinkVec_queue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_18_almostFull),
    .full         (_sinkVec_queue_fifo_18_full),
    .error        (_sinkVec_queue_fifo_18_error),
    .data_out     (_sinkVec_queue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_19_enq_ready & sinkVec_queue_19_enq_valid & ~(_sinkVec_queue_fifo_19_empty & sinkVec_queue_19_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_19_deq_ready & ~_sinkVec_queue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_19),
    .empty        (_sinkVec_queue_fifo_19_empty),
    .almost_empty (sinkVec_queue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_19_almostFull),
    .full         (_sinkVec_queue_fifo_19_full),
    .error        (_sinkVec_queue_fifo_19_error),
    .data_out     (_sinkVec_queue_fifo_19_data_out)
  );
  Lane laneVec_5 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h5),
    .readBusPort_0_enq_valid                             (shifterReg_68_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_68_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_5_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_5_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_5_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_42_valid),
    .readBusPort_1_enq_valid                             (shifterReg_70_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_70_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_5_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_5_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_5_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_74_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_59_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_59_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_59_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_59_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_59_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_5_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_5_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_5_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_5_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_5_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_5_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_53_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_91_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_91_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_91_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_91_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_91_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_5_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_5_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_5_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_5_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_5_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_5_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_55_valid),
    .laneRequest_ready                                   (_laneVec_5_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_5_valid & laneRequestSinkWire_5_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_5_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_5_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_5_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_5_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_5_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_5_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_5_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_5_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_5_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_5_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_5_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_5_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_5_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_5_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_5_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_5_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_5_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_5_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_5_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_5_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_5_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_5_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_5_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_5_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_5_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_5_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_5_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_5_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_5_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_5_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_5_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_5_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_5_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_5_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_5_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_5_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_5_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_5_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_5_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_5_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_5_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_5_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_5_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_5_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_5_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_5_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_5_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_5_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_5_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_5_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_5_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_5_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_5_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_5_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_5_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_5_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_5_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_5_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_5_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_5_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_5_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_5_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_5_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_5_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_5_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_5_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_5_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_5_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_5_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_5_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_5_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_5_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_5_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_5_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_5_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_5_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[5]),
    .vrfReadAddressChannel_ready                         (sinkWire_10_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_10_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_10_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_10_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_10_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_10_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_5_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_11_ready),
    .vrfWriteChannel_valid                               (sinkWire_11_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_11_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_11_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_11_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_11_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_11_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_11_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_5_valid_T),
    .instructionFinished                                 (_laneVec_5_instructionFinished),
    .vxsatReport                                         (_laneVec_5_vxsatReport),
    .v0Update_valid                                      (_laneVec_5_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_5_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_5_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_5_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_5_bits),
    .maskSelect                                          (_laneVec_5_maskSelect),
    .maskSelectSew                                       (_laneVec_5_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_5_bits | maskLastPipe_pipe_out_5_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_5),
    .writeCount                                          (pipe_out_11_bits),
    .writeQueueValid                                     (dataInWritePipeVec_5)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_20_enq_ready & sinkVec_queue_20_enq_valid & ~(_sinkVec_queue_fifo_20_empty & sinkVec_queue_20_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_20_deq_ready & ~_sinkVec_queue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_20),
    .empty        (_sinkVec_queue_fifo_20_empty),
    .almost_empty (sinkVec_queue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_20_almostFull),
    .full         (_sinkVec_queue_fifo_20_full),
    .error        (_sinkVec_queue_fifo_20_error),
    .data_out     (_sinkVec_queue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_21_enq_ready & sinkVec_queue_21_enq_valid & ~(_sinkVec_queue_fifo_21_empty & sinkVec_queue_21_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_21_deq_ready & ~_sinkVec_queue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_21),
    .empty        (_sinkVec_queue_fifo_21_empty),
    .almost_empty (sinkVec_queue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_21_almostFull),
    .full         (_sinkVec_queue_fifo_21_full),
    .error        (_sinkVec_queue_fifo_21_error),
    .data_out     (_sinkVec_queue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_22_enq_ready & sinkVec_queue_22_enq_valid & ~(_sinkVec_queue_fifo_22_empty & sinkVec_queue_22_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_22_deq_ready & ~_sinkVec_queue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_22),
    .empty        (_sinkVec_queue_fifo_22_empty),
    .almost_empty (sinkVec_queue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_22_almostFull),
    .full         (_sinkVec_queue_fifo_22_full),
    .error        (_sinkVec_queue_fifo_22_error),
    .data_out     (_sinkVec_queue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_23_enq_ready & sinkVec_queue_23_enq_valid & ~(_sinkVec_queue_fifo_23_empty & sinkVec_queue_23_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_23_deq_ready & ~_sinkVec_queue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_23),
    .empty        (_sinkVec_queue_fifo_23_empty),
    .almost_empty (sinkVec_queue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_23_almostFull),
    .full         (_sinkVec_queue_fifo_23_full),
    .error        (_sinkVec_queue_fifo_23_error),
    .data_out     (_sinkVec_queue_fifo_23_data_out)
  );
  Lane laneVec_6 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h6),
    .readBusPort_0_enq_valid                             (shifterReg_72_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_72_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_6_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_6_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_6_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_44_valid),
    .readBusPort_1_enq_valid                             (shifterReg_74_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_74_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_6_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_6_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_6_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_76_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_61_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_61_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_61_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_61_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_61_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_6_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_6_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_6_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_6_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_6_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_6_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_57_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_93_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_93_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_93_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_93_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_93_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_6_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_6_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_6_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_6_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_6_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_6_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_59_valid),
    .laneRequest_ready                                   (_laneVec_6_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_6_valid & laneRequestSinkWire_6_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_6_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_6_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_6_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_6_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_6_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_6_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_6_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_6_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_6_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_6_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_6_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_6_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_6_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_6_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_6_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_6_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_6_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_6_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_6_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_6_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_6_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_6_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_6_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_6_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_6_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_6_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_6_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_6_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_6_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_6_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_6_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_6_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_6_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_6_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_6_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_6_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_6_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_6_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_6_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_6_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_6_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_6_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_6_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_6_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_6_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_6_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_6_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_6_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_6_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_6_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_6_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_6_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_6_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_6_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_6_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_6_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_6_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_6_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_6_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_6_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_6_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_6_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_6_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_6_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_6_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_6_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_6_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_6_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_6_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_6_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_6_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_6_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_6_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_6_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_6_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_6_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[6]),
    .vrfReadAddressChannel_ready                         (sinkWire_12_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_12_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_12_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_12_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_12_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_12_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_6_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_13_ready),
    .vrfWriteChannel_valid                               (sinkWire_13_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_13_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_13_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_13_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_13_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_13_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_13_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_6_valid_T),
    .instructionFinished                                 (_laneVec_6_instructionFinished),
    .vxsatReport                                         (_laneVec_6_vxsatReport),
    .v0Update_valid                                      (_laneVec_6_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_6_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_6_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_6_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_6_bits),
    .maskSelect                                          (_laneVec_6_maskSelect),
    .maskSelectSew                                       (_laneVec_6_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_6_bits | maskLastPipe_pipe_out_6_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_6),
    .writeCount                                          (pipe_out_13_bits),
    .writeQueueValid                                     (dataInWritePipeVec_6)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_24_enq_ready & sinkVec_queue_24_enq_valid & ~(_sinkVec_queue_fifo_24_empty & sinkVec_queue_24_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_24_deq_ready & ~_sinkVec_queue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_24),
    .empty        (_sinkVec_queue_fifo_24_empty),
    .almost_empty (sinkVec_queue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_24_almostFull),
    .full         (_sinkVec_queue_fifo_24_full),
    .error        (_sinkVec_queue_fifo_24_error),
    .data_out     (_sinkVec_queue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_25_enq_ready & sinkVec_queue_25_enq_valid & ~(_sinkVec_queue_fifo_25_empty & sinkVec_queue_25_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_25_deq_ready & ~_sinkVec_queue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_25),
    .empty        (_sinkVec_queue_fifo_25_empty),
    .almost_empty (sinkVec_queue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_25_almostFull),
    .full         (_sinkVec_queue_fifo_25_full),
    .error        (_sinkVec_queue_fifo_25_error),
    .data_out     (_sinkVec_queue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_26_enq_ready & sinkVec_queue_26_enq_valid & ~(_sinkVec_queue_fifo_26_empty & sinkVec_queue_26_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_26_deq_ready & ~_sinkVec_queue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_26),
    .empty        (_sinkVec_queue_fifo_26_empty),
    .almost_empty (sinkVec_queue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_26_almostFull),
    .full         (_sinkVec_queue_fifo_26_full),
    .error        (_sinkVec_queue_fifo_26_error),
    .data_out     (_sinkVec_queue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_27_enq_ready & sinkVec_queue_27_enq_valid & ~(_sinkVec_queue_fifo_27_empty & sinkVec_queue_27_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_27_deq_ready & ~_sinkVec_queue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_27),
    .empty        (_sinkVec_queue_fifo_27_empty),
    .almost_empty (sinkVec_queue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_27_almostFull),
    .full         (_sinkVec_queue_fifo_27_full),
    .error        (_sinkVec_queue_fifo_27_error),
    .data_out     (_sinkVec_queue_fifo_27_data_out)
  );
  Lane laneVec_7 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h7),
    .readBusPort_0_enq_valid                             (shifterReg_76_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_76_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_7_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_7_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_7_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_46_valid),
    .readBusPort_1_enq_valid                             (shifterReg_78_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_78_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_7_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_7_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_7_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_78_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_63_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_63_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_63_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_63_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_63_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_7_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_7_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_7_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_7_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_7_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_7_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_61_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_95_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_95_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_95_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_95_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_95_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_7_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_7_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_7_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_7_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_7_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_7_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_63_valid),
    .laneRequest_ready                                   (_laneVec_7_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_7_valid & laneRequestSinkWire_7_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_7_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_7_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_7_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_7_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_7_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_7_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_7_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_7_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_7_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_7_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_7_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_7_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_7_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_7_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_7_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_7_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_7_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_7_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_7_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_7_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_7_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_7_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_7_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_7_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_7_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_7_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_7_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_7_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_7_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_7_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_7_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_7_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_7_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_7_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_7_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_7_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_7_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_7_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_7_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_7_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_7_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_7_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_7_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_7_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_7_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_7_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_7_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_7_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_7_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_7_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_7_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_7_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_7_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_7_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_7_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_7_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_7_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_7_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_7_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_7_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_7_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_7_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_7_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_7_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_7_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_7_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_7_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_7_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_7_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_7_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_7_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_7_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_7_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_7_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_7_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_7_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[7]),
    .vrfReadAddressChannel_ready                         (sinkWire_14_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_14_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_14_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_14_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_14_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_14_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_7_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_15_ready),
    .vrfWriteChannel_valid                               (sinkWire_15_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_15_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_15_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_15_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_15_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_15_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_15_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_7_valid_T),
    .instructionFinished                                 (_laneVec_7_instructionFinished),
    .vxsatReport                                         (_laneVec_7_vxsatReport),
    .v0Update_valid                                      (_laneVec_7_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_7_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_7_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_7_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_7_bits),
    .maskSelect                                          (_laneVec_7_maskSelect),
    .maskSelectSew                                       (_laneVec_7_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_7_bits | maskLastPipe_pipe_out_7_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_7),
    .writeCount                                          (pipe_out_15_bits),
    .writeQueueValid                                     (dataInWritePipeVec_7)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_28_enq_ready & sinkVec_queue_28_enq_valid & ~(_sinkVec_queue_fifo_28_empty & sinkVec_queue_28_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_28_deq_ready & ~_sinkVec_queue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_28),
    .empty        (_sinkVec_queue_fifo_28_empty),
    .almost_empty (sinkVec_queue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_28_almostFull),
    .full         (_sinkVec_queue_fifo_28_full),
    .error        (_sinkVec_queue_fifo_28_error),
    .data_out     (_sinkVec_queue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_29_enq_ready & sinkVec_queue_29_enq_valid & ~(_sinkVec_queue_fifo_29_empty & sinkVec_queue_29_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_29_deq_ready & ~_sinkVec_queue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_29),
    .empty        (_sinkVec_queue_fifo_29_empty),
    .almost_empty (sinkVec_queue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_29_almostFull),
    .full         (_sinkVec_queue_fifo_29_full),
    .error        (_sinkVec_queue_fifo_29_error),
    .data_out     (_sinkVec_queue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_30_enq_ready & sinkVec_queue_30_enq_valid & ~(_sinkVec_queue_fifo_30_empty & sinkVec_queue_30_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_30_deq_ready & ~_sinkVec_queue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_30),
    .empty        (_sinkVec_queue_fifo_30_empty),
    .almost_empty (sinkVec_queue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_30_almostFull),
    .full         (_sinkVec_queue_fifo_30_full),
    .error        (_sinkVec_queue_fifo_30_error),
    .data_out     (_sinkVec_queue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_31_enq_ready & sinkVec_queue_31_enq_valid & ~(_sinkVec_queue_fifo_31_empty & sinkVec_queue_31_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_31_deq_ready & ~_sinkVec_queue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_31),
    .empty        (_sinkVec_queue_fifo_31_empty),
    .almost_empty (sinkVec_queue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_31_almostFull),
    .full         (_sinkVec_queue_fifo_31_full),
    .error        (_sinkVec_queue_fifo_31_error),
    .data_out     (_sinkVec_queue_fifo_31_data_out)
  );
  Lane laneVec_8 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h8),
    .readBusPort_0_enq_valid                             (shifterReg_80_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_80_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_8_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_8_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_8_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_48_valid),
    .readBusPort_1_enq_valid                             (shifterReg_82_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_82_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_8_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_8_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_8_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_80_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_65_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_65_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_65_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_65_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_65_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_8_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_8_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_8_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_8_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_8_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_8_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_65_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_97_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_97_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_97_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_97_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_97_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_8_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_8_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_8_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_8_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_8_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_8_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_67_valid),
    .laneRequest_ready                                   (_laneVec_8_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_8_valid & laneRequestSinkWire_8_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_8_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_8_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_8_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_8_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_8_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_8_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_8_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_8_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_8_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_8_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_8_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_8_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_8_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_8_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_8_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_8_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_8_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_8_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_8_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_8_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_8_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_8_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_8_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_8_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_8_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_8_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_8_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_8_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_8_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_8_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_8_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_8_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_8_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_8_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_8_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_8_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_8_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_8_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_8_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_8_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_8_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_8_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_8_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_8_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_8_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_8_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_8_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_8_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_8_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_8_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_8_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_8_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_8_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_8_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_8_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_8_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_8_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_8_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_8_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_8_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_8_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_8_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_8_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_8_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_8_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_8_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_8_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_8_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_8_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_8_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_8_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_8_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_8_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_8_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_8_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_8_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[8]),
    .vrfReadAddressChannel_ready                         (sinkWire_16_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_16_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_16_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_16_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_16_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_16_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_8_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_17_ready),
    .vrfWriteChannel_valid                               (sinkWire_17_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_17_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_17_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_17_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_17_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_17_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_17_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_8_valid_T),
    .instructionFinished                                 (_laneVec_8_instructionFinished),
    .vxsatReport                                         (_laneVec_8_vxsatReport),
    .v0Update_valid                                      (_laneVec_8_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_8_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_8_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_8_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_8_bits),
    .maskSelect                                          (_laneVec_8_maskSelect),
    .maskSelectSew                                       (_laneVec_8_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_8_bits | maskLastPipe_pipe_out_8_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_8),
    .writeCount                                          (pipe_out_17_bits),
    .writeQueueValid                                     (dataInWritePipeVec_8)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_32 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_32_enq_ready & sinkVec_queue_32_enq_valid & ~(_sinkVec_queue_fifo_32_empty & sinkVec_queue_32_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_32_deq_ready & ~_sinkVec_queue_fifo_32_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_32),
    .empty        (_sinkVec_queue_fifo_32_empty),
    .almost_empty (sinkVec_queue_32_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_32_almostFull),
    .full         (_sinkVec_queue_fifo_32_full),
    .error        (_sinkVec_queue_fifo_32_error),
    .data_out     (_sinkVec_queue_fifo_32_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_33 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_33_enq_ready & sinkVec_queue_33_enq_valid & ~(_sinkVec_queue_fifo_33_empty & sinkVec_queue_33_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_33_deq_ready & ~_sinkVec_queue_fifo_33_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_33),
    .empty        (_sinkVec_queue_fifo_33_empty),
    .almost_empty (sinkVec_queue_33_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_33_almostFull),
    .full         (_sinkVec_queue_fifo_33_full),
    .error        (_sinkVec_queue_fifo_33_error),
    .data_out     (_sinkVec_queue_fifo_33_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_34 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_34_enq_ready & sinkVec_queue_34_enq_valid & ~(_sinkVec_queue_fifo_34_empty & sinkVec_queue_34_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_34_deq_ready & ~_sinkVec_queue_fifo_34_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_34),
    .empty        (_sinkVec_queue_fifo_34_empty),
    .almost_empty (sinkVec_queue_34_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_34_almostFull),
    .full         (_sinkVec_queue_fifo_34_full),
    .error        (_sinkVec_queue_fifo_34_error),
    .data_out     (_sinkVec_queue_fifo_34_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_35 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_35_enq_ready & sinkVec_queue_35_enq_valid & ~(_sinkVec_queue_fifo_35_empty & sinkVec_queue_35_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_35_deq_ready & ~_sinkVec_queue_fifo_35_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_35),
    .empty        (_sinkVec_queue_fifo_35_empty),
    .almost_empty (sinkVec_queue_35_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_35_almostFull),
    .full         (_sinkVec_queue_fifo_35_full),
    .error        (_sinkVec_queue_fifo_35_error),
    .data_out     (_sinkVec_queue_fifo_35_data_out)
  );
  Lane laneVec_9 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'h9),
    .readBusPort_0_enq_valid                             (shifterReg_84_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_84_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_9_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_9_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_9_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_50_valid),
    .readBusPort_1_enq_valid                             (shifterReg_86_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_86_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_9_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_9_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_9_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_82_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_67_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_67_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_67_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_67_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_67_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_9_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_9_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_9_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_9_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_9_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_9_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_69_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_99_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_99_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_99_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_99_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_99_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_9_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_9_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_9_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_9_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_9_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_9_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_71_valid),
    .laneRequest_ready                                   (_laneVec_9_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_9_valid & laneRequestSinkWire_9_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_9_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_9_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_9_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_9_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_9_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_9_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_9_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_9_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_9_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_9_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_9_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_9_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_9_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_9_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_9_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_9_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_9_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_9_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_9_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_9_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_9_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_9_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_9_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_9_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_9_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_9_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_9_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_9_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_9_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_9_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_9_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_9_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_9_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_9_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_9_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_9_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_9_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_9_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_9_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_9_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_9_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_9_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_9_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_9_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_9_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_9_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_9_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_9_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_9_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_9_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_9_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_9_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_9_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_9_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_9_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_9_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_9_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_9_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_9_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_9_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_9_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_9_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_9_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_9_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_9_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_9_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_9_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_9_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_9_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_9_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_9_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_9_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_9_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_9_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_9_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_9_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[9]),
    .vrfReadAddressChannel_ready                         (sinkWire_18_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_18_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_18_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_18_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_18_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_18_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_9_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_19_ready),
    .vrfWriteChannel_valid                               (sinkWire_19_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_19_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_19_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_19_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_19_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_19_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_19_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_9_valid_T),
    .instructionFinished                                 (_laneVec_9_instructionFinished),
    .vxsatReport                                         (_laneVec_9_vxsatReport),
    .v0Update_valid                                      (_laneVec_9_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_9_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_9_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_9_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_9_bits),
    .maskSelect                                          (_laneVec_9_maskSelect),
    .maskSelectSew                                       (_laneVec_9_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_9_bits | maskLastPipe_pipe_out_9_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_9),
    .writeCount                                          (pipe_out_19_bits),
    .writeQueueValid                                     (dataInWritePipeVec_9)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_36 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_36_enq_ready & sinkVec_queue_36_enq_valid & ~(_sinkVec_queue_fifo_36_empty & sinkVec_queue_36_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_36_deq_ready & ~_sinkVec_queue_fifo_36_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_36),
    .empty        (_sinkVec_queue_fifo_36_empty),
    .almost_empty (sinkVec_queue_36_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_36_almostFull),
    .full         (_sinkVec_queue_fifo_36_full),
    .error        (_sinkVec_queue_fifo_36_error),
    .data_out     (_sinkVec_queue_fifo_36_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_37 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_37_enq_ready & sinkVec_queue_37_enq_valid & ~(_sinkVec_queue_fifo_37_empty & sinkVec_queue_37_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_37_deq_ready & ~_sinkVec_queue_fifo_37_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_37),
    .empty        (_sinkVec_queue_fifo_37_empty),
    .almost_empty (sinkVec_queue_37_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_37_almostFull),
    .full         (_sinkVec_queue_fifo_37_full),
    .error        (_sinkVec_queue_fifo_37_error),
    .data_out     (_sinkVec_queue_fifo_37_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_38 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_38_enq_ready & sinkVec_queue_38_enq_valid & ~(_sinkVec_queue_fifo_38_empty & sinkVec_queue_38_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_38_deq_ready & ~_sinkVec_queue_fifo_38_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_38),
    .empty        (_sinkVec_queue_fifo_38_empty),
    .almost_empty (sinkVec_queue_38_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_38_almostFull),
    .full         (_sinkVec_queue_fifo_38_full),
    .error        (_sinkVec_queue_fifo_38_error),
    .data_out     (_sinkVec_queue_fifo_38_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_39 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_39_enq_ready & sinkVec_queue_39_enq_valid & ~(_sinkVec_queue_fifo_39_empty & sinkVec_queue_39_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_39_deq_ready & ~_sinkVec_queue_fifo_39_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_39),
    .empty        (_sinkVec_queue_fifo_39_empty),
    .almost_empty (sinkVec_queue_39_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_39_almostFull),
    .full         (_sinkVec_queue_fifo_39_full),
    .error        (_sinkVec_queue_fifo_39_error),
    .data_out     (_sinkVec_queue_fifo_39_data_out)
  );
  Lane laneVec_10 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hA),
    .readBusPort_0_enq_valid                             (shifterReg_88_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_88_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_10_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_10_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_10_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_52_valid),
    .readBusPort_1_enq_valid                             (shifterReg_90_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_90_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_10_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_10_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_10_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_84_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_69_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_69_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_69_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_69_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_69_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_10_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_10_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_10_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_10_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_10_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_10_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_73_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_101_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_101_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_101_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_101_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_101_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_10_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_10_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_10_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_10_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_10_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_10_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_75_valid),
    .laneRequest_ready                                   (_laneVec_10_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_10_valid & laneRequestSinkWire_10_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_10_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_10_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_10_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_10_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_10_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_10_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_10_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_10_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_10_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_10_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_10_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_10_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_10_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_10_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_10_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_10_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_10_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_10_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_10_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_10_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_10_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_10_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_10_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_10_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_10_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_10_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_10_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_10_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_10_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_10_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_10_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_10_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_10_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_10_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_10_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_10_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_10_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_10_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_10_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_10_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_10_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_10_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_10_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_10_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_10_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_10_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_10_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_10_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_10_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_10_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_10_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_10_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_10_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_10_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_10_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_10_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_10_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_10_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_10_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_10_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_10_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_10_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_10_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_10_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_10_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_10_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_10_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_10_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_10_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_10_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_10_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_10_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_10_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_10_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_10_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_10_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[10]),
    .vrfReadAddressChannel_ready                         (sinkWire_20_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_20_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_20_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_20_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_20_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_20_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_10_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_21_ready),
    .vrfWriteChannel_valid                               (sinkWire_21_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_21_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_21_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_21_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_21_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_21_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_21_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_10_valid_T),
    .instructionFinished                                 (_laneVec_10_instructionFinished),
    .vxsatReport                                         (_laneVec_10_vxsatReport),
    .v0Update_valid                                      (_laneVec_10_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_10_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_10_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_10_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_10_bits),
    .maskSelect                                          (_laneVec_10_maskSelect),
    .maskSelectSew                                       (_laneVec_10_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_10_bits | maskLastPipe_pipe_out_10_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_10),
    .writeCount                                          (pipe_out_21_bits),
    .writeQueueValid                                     (dataInWritePipeVec_10)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_40 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_40_enq_ready & sinkVec_queue_40_enq_valid & ~(_sinkVec_queue_fifo_40_empty & sinkVec_queue_40_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_40_deq_ready & ~_sinkVec_queue_fifo_40_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_40),
    .empty        (_sinkVec_queue_fifo_40_empty),
    .almost_empty (sinkVec_queue_40_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_40_almostFull),
    .full         (_sinkVec_queue_fifo_40_full),
    .error        (_sinkVec_queue_fifo_40_error),
    .data_out     (_sinkVec_queue_fifo_40_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_41 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_41_enq_ready & sinkVec_queue_41_enq_valid & ~(_sinkVec_queue_fifo_41_empty & sinkVec_queue_41_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_41_deq_ready & ~_sinkVec_queue_fifo_41_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_41),
    .empty        (_sinkVec_queue_fifo_41_empty),
    .almost_empty (sinkVec_queue_41_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_41_almostFull),
    .full         (_sinkVec_queue_fifo_41_full),
    .error        (_sinkVec_queue_fifo_41_error),
    .data_out     (_sinkVec_queue_fifo_41_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_42 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_42_enq_ready & sinkVec_queue_42_enq_valid & ~(_sinkVec_queue_fifo_42_empty & sinkVec_queue_42_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_42_deq_ready & ~_sinkVec_queue_fifo_42_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_42),
    .empty        (_sinkVec_queue_fifo_42_empty),
    .almost_empty (sinkVec_queue_42_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_42_almostFull),
    .full         (_sinkVec_queue_fifo_42_full),
    .error        (_sinkVec_queue_fifo_42_error),
    .data_out     (_sinkVec_queue_fifo_42_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_43 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_43_enq_ready & sinkVec_queue_43_enq_valid & ~(_sinkVec_queue_fifo_43_empty & sinkVec_queue_43_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_43_deq_ready & ~_sinkVec_queue_fifo_43_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_43),
    .empty        (_sinkVec_queue_fifo_43_empty),
    .almost_empty (sinkVec_queue_43_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_43_almostFull),
    .full         (_sinkVec_queue_fifo_43_full),
    .error        (_sinkVec_queue_fifo_43_error),
    .data_out     (_sinkVec_queue_fifo_43_data_out)
  );
  Lane laneVec_11 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hB),
    .readBusPort_0_enq_valid                             (shifterReg_92_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_92_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_11_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_11_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_11_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_54_valid),
    .readBusPort_1_enq_valid                             (shifterReg_94_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_94_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_11_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_11_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_11_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_86_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_71_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_71_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_71_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_71_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_71_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_11_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_11_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_11_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_11_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_11_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_11_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_77_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_103_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_103_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_103_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_103_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_103_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_11_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_11_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_11_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_11_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_11_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_11_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_79_valid),
    .laneRequest_ready                                   (_laneVec_11_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_11_valid & laneRequestSinkWire_11_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_11_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_11_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_11_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_11_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_11_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_11_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_11_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_11_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_11_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_11_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_11_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_11_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_11_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_11_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_11_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_11_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_11_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_11_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_11_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_11_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_11_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_11_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_11_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_11_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_11_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_11_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_11_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_11_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_11_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_11_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_11_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_11_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_11_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_11_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_11_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_11_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_11_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_11_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_11_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_11_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_11_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_11_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_11_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_11_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_11_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_11_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_11_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_11_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_11_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_11_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_11_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_11_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_11_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_11_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_11_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_11_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_11_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_11_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_11_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_11_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_11_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_11_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_11_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_11_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_11_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_11_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_11_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_11_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_11_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_11_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_11_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_11_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_11_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_11_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_11_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_11_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[11]),
    .vrfReadAddressChannel_ready                         (sinkWire_22_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_22_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_22_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_22_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_22_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_22_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_11_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_23_ready),
    .vrfWriteChannel_valid                               (sinkWire_23_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_23_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_23_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_23_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_23_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_23_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_23_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_11_valid_T),
    .instructionFinished                                 (_laneVec_11_instructionFinished),
    .vxsatReport                                         (_laneVec_11_vxsatReport),
    .v0Update_valid                                      (_laneVec_11_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_11_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_11_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_11_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_11_bits),
    .maskSelect                                          (_laneVec_11_maskSelect),
    .maskSelectSew                                       (_laneVec_11_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_11_bits | maskLastPipe_pipe_out_11_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_11),
    .writeCount                                          (pipe_out_23_bits),
    .writeQueueValid                                     (dataInWritePipeVec_11)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_44 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_44_enq_ready & sinkVec_queue_44_enq_valid & ~(_sinkVec_queue_fifo_44_empty & sinkVec_queue_44_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_44_deq_ready & ~_sinkVec_queue_fifo_44_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_44),
    .empty        (_sinkVec_queue_fifo_44_empty),
    .almost_empty (sinkVec_queue_44_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_44_almostFull),
    .full         (_sinkVec_queue_fifo_44_full),
    .error        (_sinkVec_queue_fifo_44_error),
    .data_out     (_sinkVec_queue_fifo_44_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_45 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_45_enq_ready & sinkVec_queue_45_enq_valid & ~(_sinkVec_queue_fifo_45_empty & sinkVec_queue_45_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_45_deq_ready & ~_sinkVec_queue_fifo_45_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_45),
    .empty        (_sinkVec_queue_fifo_45_empty),
    .almost_empty (sinkVec_queue_45_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_45_almostFull),
    .full         (_sinkVec_queue_fifo_45_full),
    .error        (_sinkVec_queue_fifo_45_error),
    .data_out     (_sinkVec_queue_fifo_45_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_46 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_46_enq_ready & sinkVec_queue_46_enq_valid & ~(_sinkVec_queue_fifo_46_empty & sinkVec_queue_46_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_46_deq_ready & ~_sinkVec_queue_fifo_46_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_46),
    .empty        (_sinkVec_queue_fifo_46_empty),
    .almost_empty (sinkVec_queue_46_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_46_almostFull),
    .full         (_sinkVec_queue_fifo_46_full),
    .error        (_sinkVec_queue_fifo_46_error),
    .data_out     (_sinkVec_queue_fifo_46_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_47 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_47_enq_ready & sinkVec_queue_47_enq_valid & ~(_sinkVec_queue_fifo_47_empty & sinkVec_queue_47_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_47_deq_ready & ~_sinkVec_queue_fifo_47_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_47),
    .empty        (_sinkVec_queue_fifo_47_empty),
    .almost_empty (sinkVec_queue_47_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_47_almostFull),
    .full         (_sinkVec_queue_fifo_47_full),
    .error        (_sinkVec_queue_fifo_47_error),
    .data_out     (_sinkVec_queue_fifo_47_data_out)
  );
  Lane laneVec_12 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hC),
    .readBusPort_0_enq_valid                             (shifterReg_96_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_96_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_12_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_12_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_12_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_56_valid),
    .readBusPort_1_enq_valid                             (shifterReg_98_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_98_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_12_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_12_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_12_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_88_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_73_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_73_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_73_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_73_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_73_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_12_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_12_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_12_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_12_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_12_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_12_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_81_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_105_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_105_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_105_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_105_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_105_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_12_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_12_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_12_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_12_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_12_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_12_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_83_valid),
    .laneRequest_ready                                   (_laneVec_12_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_12_valid & laneRequestSinkWire_12_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_12_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_12_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_12_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_12_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_12_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_12_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_12_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_12_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_12_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_12_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_12_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_12_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_12_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_12_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_12_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_12_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_12_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_12_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_12_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_12_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_12_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_12_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_12_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_12_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_12_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_12_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_12_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_12_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_12_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_12_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_12_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_12_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_12_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_12_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_12_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_12_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_12_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_12_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_12_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_12_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_12_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_12_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_12_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_12_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_12_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_12_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_12_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_12_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_12_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_12_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_12_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_12_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_12_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_12_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_12_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_12_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_12_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_12_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_12_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_12_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_12_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_12_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_12_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_12_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_12_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_12_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_12_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_12_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_12_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_12_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_12_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_12_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_12_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_12_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_12_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_12_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[12]),
    .vrfReadAddressChannel_ready                         (sinkWire_24_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_24_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_24_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_24_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_24_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_24_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_12_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_25_ready),
    .vrfWriteChannel_valid                               (sinkWire_25_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_25_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_25_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_25_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_25_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_25_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_25_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_12_valid_T),
    .instructionFinished                                 (_laneVec_12_instructionFinished),
    .vxsatReport                                         (_laneVec_12_vxsatReport),
    .v0Update_valid                                      (_laneVec_12_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_12_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_12_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_12_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_12_bits),
    .maskSelect                                          (_laneVec_12_maskSelect),
    .maskSelectSew                                       (_laneVec_12_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_12_bits | maskLastPipe_pipe_out_12_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_12),
    .writeCount                                          (pipe_out_25_bits),
    .writeQueueValid                                     (dataInWritePipeVec_12)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_48 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_48_enq_ready & sinkVec_queue_48_enq_valid & ~(_sinkVec_queue_fifo_48_empty & sinkVec_queue_48_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_48_deq_ready & ~_sinkVec_queue_fifo_48_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_48),
    .empty        (_sinkVec_queue_fifo_48_empty),
    .almost_empty (sinkVec_queue_48_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_48_almostFull),
    .full         (_sinkVec_queue_fifo_48_full),
    .error        (_sinkVec_queue_fifo_48_error),
    .data_out     (_sinkVec_queue_fifo_48_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_49 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_49_enq_ready & sinkVec_queue_49_enq_valid & ~(_sinkVec_queue_fifo_49_empty & sinkVec_queue_49_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_49_deq_ready & ~_sinkVec_queue_fifo_49_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_49),
    .empty        (_sinkVec_queue_fifo_49_empty),
    .almost_empty (sinkVec_queue_49_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_49_almostFull),
    .full         (_sinkVec_queue_fifo_49_full),
    .error        (_sinkVec_queue_fifo_49_error),
    .data_out     (_sinkVec_queue_fifo_49_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_50 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_50_enq_ready & sinkVec_queue_50_enq_valid & ~(_sinkVec_queue_fifo_50_empty & sinkVec_queue_50_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_50_deq_ready & ~_sinkVec_queue_fifo_50_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_50),
    .empty        (_sinkVec_queue_fifo_50_empty),
    .almost_empty (sinkVec_queue_50_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_50_almostFull),
    .full         (_sinkVec_queue_fifo_50_full),
    .error        (_sinkVec_queue_fifo_50_error),
    .data_out     (_sinkVec_queue_fifo_50_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_51 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_51_enq_ready & sinkVec_queue_51_enq_valid & ~(_sinkVec_queue_fifo_51_empty & sinkVec_queue_51_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_51_deq_ready & ~_sinkVec_queue_fifo_51_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_51),
    .empty        (_sinkVec_queue_fifo_51_empty),
    .almost_empty (sinkVec_queue_51_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_51_almostFull),
    .full         (_sinkVec_queue_fifo_51_full),
    .error        (_sinkVec_queue_fifo_51_error),
    .data_out     (_sinkVec_queue_fifo_51_data_out)
  );
  Lane laneVec_13 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hD),
    .readBusPort_0_enq_valid                             (shifterReg_100_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_100_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_13_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_13_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_13_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_58_valid),
    .readBusPort_1_enq_valid                             (shifterReg_102_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_102_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_13_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_13_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_13_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_90_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_75_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_75_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_75_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_75_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_75_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_13_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_13_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_13_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_13_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_13_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_13_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_85_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_107_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_107_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_107_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_107_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_107_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_13_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_13_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_13_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_13_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_13_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_13_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_87_valid),
    .laneRequest_ready                                   (_laneVec_13_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_13_valid & laneRequestSinkWire_13_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_13_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_13_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_13_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_13_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_13_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_13_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_13_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_13_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_13_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_13_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_13_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_13_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_13_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_13_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_13_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_13_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_13_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_13_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_13_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_13_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_13_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_13_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_13_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_13_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_13_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_13_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_13_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_13_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_13_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_13_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_13_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_13_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_13_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_13_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_13_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_13_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_13_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_13_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_13_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_13_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_13_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_13_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_13_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_13_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_13_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_13_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_13_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_13_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_13_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_13_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_13_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_13_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_13_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_13_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_13_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_13_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_13_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_13_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_13_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_13_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_13_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_13_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_13_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_13_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_13_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_13_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_13_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_13_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_13_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_13_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_13_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_13_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_13_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_13_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_13_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_13_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[13]),
    .vrfReadAddressChannel_ready                         (sinkWire_26_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_26_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_26_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_26_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_26_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_26_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_13_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_27_ready),
    .vrfWriteChannel_valid                               (sinkWire_27_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_27_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_27_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_27_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_27_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_27_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_27_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_13_valid_T),
    .instructionFinished                                 (_laneVec_13_instructionFinished),
    .vxsatReport                                         (_laneVec_13_vxsatReport),
    .v0Update_valid                                      (_laneVec_13_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_13_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_13_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_13_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_13_bits),
    .maskSelect                                          (_laneVec_13_maskSelect),
    .maskSelectSew                                       (_laneVec_13_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_13_bits | maskLastPipe_pipe_out_13_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_13),
    .writeCount                                          (pipe_out_27_bits),
    .writeQueueValid                                     (dataInWritePipeVec_13)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_52 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_52_enq_ready & sinkVec_queue_52_enq_valid & ~(_sinkVec_queue_fifo_52_empty & sinkVec_queue_52_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_52_deq_ready & ~_sinkVec_queue_fifo_52_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_52),
    .empty        (_sinkVec_queue_fifo_52_empty),
    .almost_empty (sinkVec_queue_52_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_52_almostFull),
    .full         (_sinkVec_queue_fifo_52_full),
    .error        (_sinkVec_queue_fifo_52_error),
    .data_out     (_sinkVec_queue_fifo_52_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_53 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_53_enq_ready & sinkVec_queue_53_enq_valid & ~(_sinkVec_queue_fifo_53_empty & sinkVec_queue_53_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_53_deq_ready & ~_sinkVec_queue_fifo_53_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_53),
    .empty        (_sinkVec_queue_fifo_53_empty),
    .almost_empty (sinkVec_queue_53_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_53_almostFull),
    .full         (_sinkVec_queue_fifo_53_full),
    .error        (_sinkVec_queue_fifo_53_error),
    .data_out     (_sinkVec_queue_fifo_53_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_54 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_54_enq_ready & sinkVec_queue_54_enq_valid & ~(_sinkVec_queue_fifo_54_empty & sinkVec_queue_54_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_54_deq_ready & ~_sinkVec_queue_fifo_54_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_54),
    .empty        (_sinkVec_queue_fifo_54_empty),
    .almost_empty (sinkVec_queue_54_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_54_almostFull),
    .full         (_sinkVec_queue_fifo_54_full),
    .error        (_sinkVec_queue_fifo_54_error),
    .data_out     (_sinkVec_queue_fifo_54_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_55 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_55_enq_ready & sinkVec_queue_55_enq_valid & ~(_sinkVec_queue_fifo_55_empty & sinkVec_queue_55_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_55_deq_ready & ~_sinkVec_queue_fifo_55_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_55),
    .empty        (_sinkVec_queue_fifo_55_empty),
    .almost_empty (sinkVec_queue_55_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_55_almostFull),
    .full         (_sinkVec_queue_fifo_55_full),
    .error        (_sinkVec_queue_fifo_55_error),
    .data_out     (_sinkVec_queue_fifo_55_data_out)
  );
  Lane laneVec_14 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hE),
    .readBusPort_0_enq_valid                             (shifterReg_104_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_104_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_14_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_14_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_14_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_60_valid),
    .readBusPort_1_enq_valid                             (shifterReg_106_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_106_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_14_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_14_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_14_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_92_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_77_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_77_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_77_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_77_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_77_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_14_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_14_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_14_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_14_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_14_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_14_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_89_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_109_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_109_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_109_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_109_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_109_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_14_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_14_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_14_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_14_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_14_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_14_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_91_valid),
    .laneRequest_ready                                   (_laneVec_14_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_14_valid & laneRequestSinkWire_14_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_14_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_14_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_14_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_14_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_14_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_14_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_14_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_14_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_14_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_14_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_14_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_14_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_14_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_14_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_14_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_14_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_14_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_14_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_14_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_14_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_14_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_14_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_14_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_14_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_14_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_14_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_14_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_14_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_14_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_14_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_14_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_14_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_14_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_14_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_14_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_14_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_14_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_14_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_14_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_14_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_14_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_14_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_14_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_14_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_14_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_14_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_14_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_14_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_14_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_14_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_14_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_14_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_14_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_14_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_14_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_14_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_14_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_14_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_14_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_14_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_14_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_14_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_14_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_14_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_14_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_14_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_14_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_14_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_14_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_14_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_14_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_14_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_14_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_14_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_14_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_14_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[14]),
    .vrfReadAddressChannel_ready                         (sinkWire_28_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_28_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_28_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_28_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_28_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_28_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_14_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_29_ready),
    .vrfWriteChannel_valid                               (sinkWire_29_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_29_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_29_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_29_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_29_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_29_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_29_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_14_valid_T),
    .instructionFinished                                 (_laneVec_14_instructionFinished),
    .vxsatReport                                         (_laneVec_14_vxsatReport),
    .v0Update_valid                                      (_laneVec_14_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_14_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_14_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_14_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_14_bits),
    .maskSelect                                          (_laneVec_14_maskSelect),
    .maskSelectSew                                       (_laneVec_14_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_14_bits | maskLastPipe_pipe_out_14_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_14),
    .writeCount                                          (pipe_out_29_bits),
    .writeQueueValid                                     (dataInWritePipeVec_14)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_56 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_56_enq_ready & sinkVec_queue_56_enq_valid & ~(_sinkVec_queue_fifo_56_empty & sinkVec_queue_56_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_56_deq_ready & ~_sinkVec_queue_fifo_56_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_56),
    .empty        (_sinkVec_queue_fifo_56_empty),
    .almost_empty (sinkVec_queue_56_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_56_almostFull),
    .full         (_sinkVec_queue_fifo_56_full),
    .error        (_sinkVec_queue_fifo_56_error),
    .data_out     (_sinkVec_queue_fifo_56_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_57 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_57_enq_ready & sinkVec_queue_57_enq_valid & ~(_sinkVec_queue_fifo_57_empty & sinkVec_queue_57_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_57_deq_ready & ~_sinkVec_queue_fifo_57_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_57),
    .empty        (_sinkVec_queue_fifo_57_empty),
    .almost_empty (sinkVec_queue_57_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_57_almostFull),
    .full         (_sinkVec_queue_fifo_57_full),
    .error        (_sinkVec_queue_fifo_57_error),
    .data_out     (_sinkVec_queue_fifo_57_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_58 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_58_enq_ready & sinkVec_queue_58_enq_valid & ~(_sinkVec_queue_fifo_58_empty & sinkVec_queue_58_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_58_deq_ready & ~_sinkVec_queue_fifo_58_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_58),
    .empty        (_sinkVec_queue_fifo_58_empty),
    .almost_empty (sinkVec_queue_58_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_58_almostFull),
    .full         (_sinkVec_queue_fifo_58_full),
    .error        (_sinkVec_queue_fifo_58_error),
    .data_out     (_sinkVec_queue_fifo_58_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_59 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_59_enq_ready & sinkVec_queue_59_enq_valid & ~(_sinkVec_queue_fifo_59_empty & sinkVec_queue_59_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_59_deq_ready & ~_sinkVec_queue_fifo_59_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_59),
    .empty        (_sinkVec_queue_fifo_59_empty),
    .almost_empty (sinkVec_queue_59_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_59_almostFull),
    .full         (_sinkVec_queue_fifo_59_full),
    .error        (_sinkVec_queue_fifo_59_error),
    .data_out     (_sinkVec_queue_fifo_59_data_out)
  );
  Lane laneVec_15 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (4'hF),
    .readBusPort_0_enq_valid                             (shifterReg_108_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_108_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_15_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_15_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_15_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_62_valid),
    .readBusPort_1_enq_valid                             (shifterReg_110_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_110_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_15_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_15_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_15_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_94_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_79_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_79_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_79_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_79_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_79_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_15_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_15_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_15_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_15_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_15_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_15_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_93_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_111_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_111_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_111_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_111_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_111_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_15_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_15_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_15_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_15_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_15_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_15_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_95_valid),
    .laneRequest_ready                                   (_laneVec_15_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_15_valid & laneRequestSinkWire_15_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_15_bits_instructionIndex),
    .laneRequest_bits_decodeResult_orderReduce           (laneRequestSinkWire_15_bits_decodeResult_orderReduce),
    .laneRequest_bits_decodeResult_floatMul              (laneRequestSinkWire_15_bits_decodeResult_floatMul),
    .laneRequest_bits_decodeResult_fpExecutionType       (laneRequestSinkWire_15_bits_decodeResult_fpExecutionType),
    .laneRequest_bits_decodeResult_float                 (laneRequestSinkWire_15_bits_decodeResult_float),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_15_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_15_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_15_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_15_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_15_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_15_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_15_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_15_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_15_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_15_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_15_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_15_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_15_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_15_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_15_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_15_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_15_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_15_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_15_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_15_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_15_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_15_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_15_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_15_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_15_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_15_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_15_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_15_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_15_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_15_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_15_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_15_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_15_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_15_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_15_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_15_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_15_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_15_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_15_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_15_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_15_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_15_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_15_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_15_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_15_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_15_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_15_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_15_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_15_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_15_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_15_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_15_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_15_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_15_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_15_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_15_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_15_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_15_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_15_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_15_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_15_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_15_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_15_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_15_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_15_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_15_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_15_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_15_maskUnitRequest_bits_ffo),
    .maskUnitRequest_bits_fpReduceValid                  (_laneVec_15_maskUnitRequest_bits_fpReduceValid),
    .maskRequestToLSU                                    (_laneVec_15_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_15_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[15]),
    .vrfReadAddressChannel_ready                         (sinkWire_30_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_30_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_30_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_30_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_30_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_30_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_15_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_31_ready),
    .vrfWriteChannel_valid                               (sinkWire_31_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_31_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_31_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_31_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_31_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_31_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_31_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_15_valid_T),
    .instructionFinished                                 (_laneVec_15_instructionFinished),
    .vxsatReport                                         (_laneVec_15_vxsatReport),
    .v0Update_valid                                      (_laneVec_15_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_15_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_15_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_15_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_15_bits),
    .maskSelect                                          (_laneVec_15_maskSelect),
    .maskSelectSew                                       (_laneVec_15_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_15_bits | maskLastPipe_pipe_out_15_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_15),
    .writeCount                                          (pipe_out_31_bits),
    .writeQueueValid                                     (dataInWritePipeVec_15)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_60 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_60_enq_ready & sinkVec_queue_60_enq_valid & ~(_sinkVec_queue_fifo_60_empty & sinkVec_queue_60_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_60_deq_ready & ~_sinkVec_queue_fifo_60_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_60),
    .empty        (_sinkVec_queue_fifo_60_empty),
    .almost_empty (sinkVec_queue_60_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_60_almostFull),
    .full         (_sinkVec_queue_fifo_60_full),
    .error        (_sinkVec_queue_fifo_60_error),
    .data_out     (_sinkVec_queue_fifo_60_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sinkVec_queue_fifo_61 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_61_enq_ready & sinkVec_queue_61_enq_valid & ~(_sinkVec_queue_fifo_61_empty & sinkVec_queue_61_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_61_deq_ready & ~_sinkVec_queue_fifo_61_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_61),
    .empty        (_sinkVec_queue_fifo_61_empty),
    .almost_empty (sinkVec_queue_61_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_61_almostFull),
    .full         (_sinkVec_queue_fifo_61_full),
    .error        (_sinkVec_queue_fifo_61_error),
    .data_out     (_sinkVec_queue_fifo_61_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_62 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_62_enq_ready & sinkVec_queue_62_enq_valid & ~(_sinkVec_queue_fifo_62_empty & sinkVec_queue_62_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_62_deq_ready & ~_sinkVec_queue_fifo_62_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_62),
    .empty        (_sinkVec_queue_fifo_62_empty),
    .almost_empty (sinkVec_queue_62_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_62_almostFull),
    .full         (_sinkVec_queue_fifo_62_full),
    .error        (_sinkVec_queue_fifo_62_error),
    .data_out     (_sinkVec_queue_fifo_62_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(47)
  ) sinkVec_queue_fifo_63 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_63_enq_ready & sinkVec_queue_63_enq_valid & ~(_sinkVec_queue_fifo_63_empty & sinkVec_queue_63_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_63_deq_ready & ~_sinkVec_queue_fifo_63_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_63),
    .empty        (_sinkVec_queue_fifo_63_empty),
    .almost_empty (sinkVec_queue_63_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_63_almostFull),
    .full         (_sinkVec_queue_fifo_63_full),
    .error        (_sinkVec_queue_fifo_63_error),
    .data_out     (_sinkVec_queue_fifo_63_data_out)
  );
  assign indexedLoadStorePort_aw_valid = indexedLoadStorePort_aw_valid_0;
  assign indexedLoadStorePort_aw_bits_id = indexedLoadStorePort_aw_bits_id_0;
  assign indexedLoadStorePort_aw_bits_addr = indexedLoadStorePort_aw_bits_addr_0;
  assign indexedLoadStorePort_aw_bits_len = 8'h0;
  assign indexedLoadStorePort_aw_bits_size = indexedLoadStorePort_aw_bits_size_0;
  assign indexedLoadStorePort_aw_bits_burst = 2'h1;
  assign indexedLoadStorePort_aw_bits_lock = 1'h0;
  assign indexedLoadStorePort_aw_bits_cache = 4'h0;
  assign indexedLoadStorePort_aw_bits_prot = 3'h0;
  assign indexedLoadStorePort_aw_bits_qos = 4'h0;
  assign indexedLoadStorePort_aw_bits_region = 4'h0;
  assign indexedLoadStorePort_w_valid = indexedLoadStorePort_w_valid_0;
  assign indexedLoadStorePort_w_bits_data = indexedLoadStorePort_w_bits_data_0;
  assign indexedLoadStorePort_w_bits_strb = indexedLoadStorePort_w_bits_strb_0;
  assign indexedLoadStorePort_w_bits_last = 1'h1;
  assign indexedLoadStorePort_b_ready = 1'h1;
  assign indexedLoadStorePort_ar_valid = indexedLoadStorePort_ar_valid_0;
  assign indexedLoadStorePort_ar_bits_id = 2'h0;
  assign indexedLoadStorePort_ar_bits_addr = indexedLoadStorePort_ar_bits_addr_0;
  assign indexedLoadStorePort_ar_bits_len = 8'h0;
  assign indexedLoadStorePort_ar_bits_size = 3'h2;
  assign indexedLoadStorePort_ar_bits_burst = 2'h1;
  assign indexedLoadStorePort_ar_bits_lock = 1'h0;
  assign indexedLoadStorePort_ar_bits_cache = 4'h0;
  assign indexedLoadStorePort_ar_bits_prot = 3'h0;
  assign indexedLoadStorePort_ar_bits_qos = 4'h0;
  assign indexedLoadStorePort_ar_bits_region = 4'h0;
  assign indexedLoadStorePort_r_ready = indexedLoadStorePort_r_ready_0;
  assign highBandwidthLoadStorePort_aw_valid = highBandwidthLoadStorePort_aw_valid_0;
  assign highBandwidthLoadStorePort_aw_bits_id = highBandwidthLoadStorePort_aw_bits_id_0;
  assign highBandwidthLoadStorePort_aw_bits_addr = highBandwidthLoadStorePort_aw_bits_addr_0;
  assign highBandwidthLoadStorePort_aw_bits_len = 8'h0;
  assign highBandwidthLoadStorePort_aw_bits_size = 3'h6;
  assign highBandwidthLoadStorePort_aw_bits_burst = 2'h1;
  assign highBandwidthLoadStorePort_aw_bits_lock = 1'h0;
  assign highBandwidthLoadStorePort_aw_bits_cache = 4'h0;
  assign highBandwidthLoadStorePort_aw_bits_prot = 3'h0;
  assign highBandwidthLoadStorePort_aw_bits_qos = 4'h0;
  assign highBandwidthLoadStorePort_aw_bits_region = 4'h0;
  assign highBandwidthLoadStorePort_w_valid = highBandwidthLoadStorePort_w_valid_0;
  assign highBandwidthLoadStorePort_w_bits_data = highBandwidthLoadStorePort_w_bits_data_0;
  assign highBandwidthLoadStorePort_w_bits_strb = highBandwidthLoadStorePort_w_bits_strb_0;
  assign highBandwidthLoadStorePort_w_bits_last = 1'h1;
  assign highBandwidthLoadStorePort_b_ready = 1'h1;
  assign highBandwidthLoadStorePort_ar_valid = highBandwidthLoadStorePort_ar_valid_0;
  assign highBandwidthLoadStorePort_ar_bits_id = 2'h0;
  assign highBandwidthLoadStorePort_ar_bits_addr = highBandwidthLoadStorePort_ar_bits_addr_0;
  assign highBandwidthLoadStorePort_ar_bits_len = 8'h0;
  assign highBandwidthLoadStorePort_ar_bits_size = 3'h6;
  assign highBandwidthLoadStorePort_ar_bits_burst = 2'h1;
  assign highBandwidthLoadStorePort_ar_bits_lock = 1'h0;
  assign highBandwidthLoadStorePort_ar_bits_cache = 4'h0;
  assign highBandwidthLoadStorePort_ar_bits_prot = 3'h0;
  assign highBandwidthLoadStorePort_ar_bits_qos = 4'h0;
  assign highBandwidthLoadStorePort_ar_bits_region = 4'h0;
  assign highBandwidthLoadStorePort_r_ready = highBandwidthLoadStorePort_r_ready_0;
  assign retire_rd_valid = retire_rd_valid_0;
  assign retire_rd_bits_rdAddress = retire_rd_bits_rdAddress_0;
  assign retire_rd_bits_rdData = retire_rd_bits_rdData_0;
  assign retire_rd_bits_isFp = retire_rd_bits_isFp_0;
  assign retire_csr_valid = 1'h0;
  assign retire_csr_bits_vxsat = retire_csr_bits_vxsat_0;
  assign retire_csr_bits_fflag = 32'h0;
  assign retire_mem_valid = retire_mem_valid_0;
  assign issue_ready = issue_ready_0;
endmodule

