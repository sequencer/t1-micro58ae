module MaskExtend(
  input  [1:0]    in_eew,
  input  [2:0]    in_uop,
  input  [1023:0] in_source2,
  input  [5:0]    in_groupCounter,
  output [1023:0] out
);

  wire [3:0]    _eew1H_T = 4'h1 << in_eew;
  wire [2:0]    eew1H = _eew1H_T[2:0];
  wire          isMaskDestination = in_uop == 3'h0;
  wire [31:0]   sourceDataVec_0 = in_source2[31:0];
  wire [31:0]   sourceDataVec_1 = in_source2[63:32];
  wire [31:0]   sourceDataVec_2 = in_source2[95:64];
  wire [31:0]   sourceDataVec_3 = in_source2[127:96];
  wire [31:0]   sourceDataVec_4 = in_source2[159:128];
  wire [31:0]   sourceDataVec_5 = in_source2[191:160];
  wire [31:0]   sourceDataVec_6 = in_source2[223:192];
  wire [31:0]   sourceDataVec_7 = in_source2[255:224];
  wire [31:0]   sourceDataVec_8 = in_source2[287:256];
  wire [31:0]   sourceDataVec_9 = in_source2[319:288];
  wire [31:0]   sourceDataVec_10 = in_source2[351:320];
  wire [31:0]   sourceDataVec_11 = in_source2[383:352];
  wire [31:0]   sourceDataVec_12 = in_source2[415:384];
  wire [31:0]   sourceDataVec_13 = in_source2[447:416];
  wire [31:0]   sourceDataVec_14 = in_source2[479:448];
  wire [31:0]   sourceDataVec_15 = in_source2[511:480];
  wire [31:0]   sourceDataVec_16 = in_source2[543:512];
  wire [31:0]   sourceDataVec_17 = in_source2[575:544];
  wire [31:0]   sourceDataVec_18 = in_source2[607:576];
  wire [31:0]   sourceDataVec_19 = in_source2[639:608];
  wire [31:0]   sourceDataVec_20 = in_source2[671:640];
  wire [31:0]   sourceDataVec_21 = in_source2[703:672];
  wire [31:0]   sourceDataVec_22 = in_source2[735:704];
  wire [31:0]   sourceDataVec_23 = in_source2[767:736];
  wire [31:0]   sourceDataVec_24 = in_source2[799:768];
  wire [31:0]   sourceDataVec_25 = in_source2[831:800];
  wire [31:0]   sourceDataVec_26 = in_source2[863:832];
  wire [31:0]   sourceDataVec_27 = in_source2[895:864];
  wire [31:0]   sourceDataVec_28 = in_source2[927:896];
  wire [31:0]   sourceDataVec_29 = in_source2[959:928];
  wire [31:0]   sourceDataVec_30 = in_source2[991:960];
  wire [31:0]   sourceDataVec_31 = in_source2[1023:992];
  wire [1:0]    maskDestinationResult_lo = sourceDataVec_0[1:0];
  wire [1:0]    maskDestinationResult_hi = sourceDataVec_0[3:2];
  wire [1:0]    maskDestinationResult_lo_1 = sourceDataVec_0[5:4];
  wire [1:0]    maskDestinationResult_hi_1 = sourceDataVec_0[7:6];
  wire [1:0]    maskDestinationResult_lo_2 = sourceDataVec_0[9:8];
  wire [1:0]    maskDestinationResult_hi_2 = sourceDataVec_0[11:10];
  wire [1:0]    maskDestinationResult_lo_3 = sourceDataVec_0[13:12];
  wire [1:0]    maskDestinationResult_hi_3 = sourceDataVec_0[15:14];
  wire [1:0]    maskDestinationResult_lo_4 = sourceDataVec_0[17:16];
  wire [1:0]    maskDestinationResult_hi_4 = sourceDataVec_0[19:18];
  wire [1:0]    maskDestinationResult_lo_5 = sourceDataVec_0[21:20];
  wire [1:0]    maskDestinationResult_hi_5 = sourceDataVec_0[23:22];
  wire [1:0]    maskDestinationResult_lo_6 = sourceDataVec_0[25:24];
  wire [1:0]    maskDestinationResult_hi_6 = sourceDataVec_0[27:26];
  wire [1:0]    maskDestinationResult_lo_7 = sourceDataVec_0[29:28];
  wire [1:0]    maskDestinationResult_hi_7 = sourceDataVec_0[31:30];
  wire [1:0]    maskDestinationResult_lo_8 = sourceDataVec_1[1:0];
  wire [1:0]    maskDestinationResult_hi_8 = sourceDataVec_1[3:2];
  wire [1:0]    maskDestinationResult_lo_9 = sourceDataVec_1[5:4];
  wire [1:0]    maskDestinationResult_hi_9 = sourceDataVec_1[7:6];
  wire [1:0]    maskDestinationResult_lo_10 = sourceDataVec_1[9:8];
  wire [1:0]    maskDestinationResult_hi_10 = sourceDataVec_1[11:10];
  wire [1:0]    maskDestinationResult_lo_11 = sourceDataVec_1[13:12];
  wire [1:0]    maskDestinationResult_hi_11 = sourceDataVec_1[15:14];
  wire [1:0]    maskDestinationResult_lo_12 = sourceDataVec_1[17:16];
  wire [1:0]    maskDestinationResult_hi_12 = sourceDataVec_1[19:18];
  wire [1:0]    maskDestinationResult_lo_13 = sourceDataVec_1[21:20];
  wire [1:0]    maskDestinationResult_hi_13 = sourceDataVec_1[23:22];
  wire [1:0]    maskDestinationResult_lo_14 = sourceDataVec_1[25:24];
  wire [1:0]    maskDestinationResult_hi_14 = sourceDataVec_1[27:26];
  wire [1:0]    maskDestinationResult_lo_15 = sourceDataVec_1[29:28];
  wire [1:0]    maskDestinationResult_hi_15 = sourceDataVec_1[31:30];
  wire [1:0]    maskDestinationResult_lo_16 = sourceDataVec_2[1:0];
  wire [1:0]    maskDestinationResult_hi_16 = sourceDataVec_2[3:2];
  wire [1:0]    maskDestinationResult_lo_17 = sourceDataVec_2[5:4];
  wire [1:0]    maskDestinationResult_hi_17 = sourceDataVec_2[7:6];
  wire [1:0]    maskDestinationResult_lo_18 = sourceDataVec_2[9:8];
  wire [1:0]    maskDestinationResult_hi_18 = sourceDataVec_2[11:10];
  wire [1:0]    maskDestinationResult_lo_19 = sourceDataVec_2[13:12];
  wire [1:0]    maskDestinationResult_hi_19 = sourceDataVec_2[15:14];
  wire [1:0]    maskDestinationResult_lo_20 = sourceDataVec_2[17:16];
  wire [1:0]    maskDestinationResult_hi_20 = sourceDataVec_2[19:18];
  wire [1:0]    maskDestinationResult_lo_21 = sourceDataVec_2[21:20];
  wire [1:0]    maskDestinationResult_hi_21 = sourceDataVec_2[23:22];
  wire [1:0]    maskDestinationResult_lo_22 = sourceDataVec_2[25:24];
  wire [1:0]    maskDestinationResult_hi_22 = sourceDataVec_2[27:26];
  wire [1:0]    maskDestinationResult_lo_23 = sourceDataVec_2[29:28];
  wire [1:0]    maskDestinationResult_hi_23 = sourceDataVec_2[31:30];
  wire [1:0]    maskDestinationResult_lo_24 = sourceDataVec_3[1:0];
  wire [1:0]    maskDestinationResult_hi_24 = sourceDataVec_3[3:2];
  wire [1:0]    maskDestinationResult_lo_25 = sourceDataVec_3[5:4];
  wire [1:0]    maskDestinationResult_hi_25 = sourceDataVec_3[7:6];
  wire [1:0]    maskDestinationResult_lo_26 = sourceDataVec_3[9:8];
  wire [1:0]    maskDestinationResult_hi_26 = sourceDataVec_3[11:10];
  wire [1:0]    maskDestinationResult_lo_27 = sourceDataVec_3[13:12];
  wire [1:0]    maskDestinationResult_hi_27 = sourceDataVec_3[15:14];
  wire [1:0]    maskDestinationResult_lo_28 = sourceDataVec_3[17:16];
  wire [1:0]    maskDestinationResult_hi_28 = sourceDataVec_3[19:18];
  wire [1:0]    maskDestinationResult_lo_29 = sourceDataVec_3[21:20];
  wire [1:0]    maskDestinationResult_hi_29 = sourceDataVec_3[23:22];
  wire [1:0]    maskDestinationResult_lo_30 = sourceDataVec_3[25:24];
  wire [1:0]    maskDestinationResult_hi_30 = sourceDataVec_3[27:26];
  wire [1:0]    maskDestinationResult_lo_31 = sourceDataVec_3[29:28];
  wire [1:0]    maskDestinationResult_hi_31 = sourceDataVec_3[31:30];
  wire [1:0]    maskDestinationResult_lo_32 = sourceDataVec_4[1:0];
  wire [1:0]    maskDestinationResult_hi_32 = sourceDataVec_4[3:2];
  wire [1:0]    maskDestinationResult_lo_33 = sourceDataVec_4[5:4];
  wire [1:0]    maskDestinationResult_hi_33 = sourceDataVec_4[7:6];
  wire [1:0]    maskDestinationResult_lo_34 = sourceDataVec_4[9:8];
  wire [1:0]    maskDestinationResult_hi_34 = sourceDataVec_4[11:10];
  wire [1:0]    maskDestinationResult_lo_35 = sourceDataVec_4[13:12];
  wire [1:0]    maskDestinationResult_hi_35 = sourceDataVec_4[15:14];
  wire [1:0]    maskDestinationResult_lo_36 = sourceDataVec_4[17:16];
  wire [1:0]    maskDestinationResult_hi_36 = sourceDataVec_4[19:18];
  wire [1:0]    maskDestinationResult_lo_37 = sourceDataVec_4[21:20];
  wire [1:0]    maskDestinationResult_hi_37 = sourceDataVec_4[23:22];
  wire [1:0]    maskDestinationResult_lo_38 = sourceDataVec_4[25:24];
  wire [1:0]    maskDestinationResult_hi_38 = sourceDataVec_4[27:26];
  wire [1:0]    maskDestinationResult_lo_39 = sourceDataVec_4[29:28];
  wire [1:0]    maskDestinationResult_hi_39 = sourceDataVec_4[31:30];
  wire [1:0]    maskDestinationResult_lo_40 = sourceDataVec_5[1:0];
  wire [1:0]    maskDestinationResult_hi_40 = sourceDataVec_5[3:2];
  wire [1:0]    maskDestinationResult_lo_41 = sourceDataVec_5[5:4];
  wire [1:0]    maskDestinationResult_hi_41 = sourceDataVec_5[7:6];
  wire [1:0]    maskDestinationResult_lo_42 = sourceDataVec_5[9:8];
  wire [1:0]    maskDestinationResult_hi_42 = sourceDataVec_5[11:10];
  wire [1:0]    maskDestinationResult_lo_43 = sourceDataVec_5[13:12];
  wire [1:0]    maskDestinationResult_hi_43 = sourceDataVec_5[15:14];
  wire [1:0]    maskDestinationResult_lo_44 = sourceDataVec_5[17:16];
  wire [1:0]    maskDestinationResult_hi_44 = sourceDataVec_5[19:18];
  wire [1:0]    maskDestinationResult_lo_45 = sourceDataVec_5[21:20];
  wire [1:0]    maskDestinationResult_hi_45 = sourceDataVec_5[23:22];
  wire [1:0]    maskDestinationResult_lo_46 = sourceDataVec_5[25:24];
  wire [1:0]    maskDestinationResult_hi_46 = sourceDataVec_5[27:26];
  wire [1:0]    maskDestinationResult_lo_47 = sourceDataVec_5[29:28];
  wire [1:0]    maskDestinationResult_hi_47 = sourceDataVec_5[31:30];
  wire [1:0]    maskDestinationResult_lo_48 = sourceDataVec_6[1:0];
  wire [1:0]    maskDestinationResult_hi_48 = sourceDataVec_6[3:2];
  wire [1:0]    maskDestinationResult_lo_49 = sourceDataVec_6[5:4];
  wire [1:0]    maskDestinationResult_hi_49 = sourceDataVec_6[7:6];
  wire [1:0]    maskDestinationResult_lo_50 = sourceDataVec_6[9:8];
  wire [1:0]    maskDestinationResult_hi_50 = sourceDataVec_6[11:10];
  wire [1:0]    maskDestinationResult_lo_51 = sourceDataVec_6[13:12];
  wire [1:0]    maskDestinationResult_hi_51 = sourceDataVec_6[15:14];
  wire [1:0]    maskDestinationResult_lo_52 = sourceDataVec_6[17:16];
  wire [1:0]    maskDestinationResult_hi_52 = sourceDataVec_6[19:18];
  wire [1:0]    maskDestinationResult_lo_53 = sourceDataVec_6[21:20];
  wire [1:0]    maskDestinationResult_hi_53 = sourceDataVec_6[23:22];
  wire [1:0]    maskDestinationResult_lo_54 = sourceDataVec_6[25:24];
  wire [1:0]    maskDestinationResult_hi_54 = sourceDataVec_6[27:26];
  wire [1:0]    maskDestinationResult_lo_55 = sourceDataVec_6[29:28];
  wire [1:0]    maskDestinationResult_hi_55 = sourceDataVec_6[31:30];
  wire [1:0]    maskDestinationResult_lo_56 = sourceDataVec_7[1:0];
  wire [1:0]    maskDestinationResult_hi_56 = sourceDataVec_7[3:2];
  wire [1:0]    maskDestinationResult_lo_57 = sourceDataVec_7[5:4];
  wire [1:0]    maskDestinationResult_hi_57 = sourceDataVec_7[7:6];
  wire [1:0]    maskDestinationResult_lo_58 = sourceDataVec_7[9:8];
  wire [1:0]    maskDestinationResult_hi_58 = sourceDataVec_7[11:10];
  wire [1:0]    maskDestinationResult_lo_59 = sourceDataVec_7[13:12];
  wire [1:0]    maskDestinationResult_hi_59 = sourceDataVec_7[15:14];
  wire [1:0]    maskDestinationResult_lo_60 = sourceDataVec_7[17:16];
  wire [1:0]    maskDestinationResult_hi_60 = sourceDataVec_7[19:18];
  wire [1:0]    maskDestinationResult_lo_61 = sourceDataVec_7[21:20];
  wire [1:0]    maskDestinationResult_hi_61 = sourceDataVec_7[23:22];
  wire [1:0]    maskDestinationResult_lo_62 = sourceDataVec_7[25:24];
  wire [1:0]    maskDestinationResult_hi_62 = sourceDataVec_7[27:26];
  wire [1:0]    maskDestinationResult_lo_63 = sourceDataVec_7[29:28];
  wire [1:0]    maskDestinationResult_hi_63 = sourceDataVec_7[31:30];
  wire [1:0]    maskDestinationResult_lo_64 = sourceDataVec_8[1:0];
  wire [1:0]    maskDestinationResult_hi_64 = sourceDataVec_8[3:2];
  wire [1:0]    maskDestinationResult_lo_65 = sourceDataVec_8[5:4];
  wire [1:0]    maskDestinationResult_hi_65 = sourceDataVec_8[7:6];
  wire [1:0]    maskDestinationResult_lo_66 = sourceDataVec_8[9:8];
  wire [1:0]    maskDestinationResult_hi_66 = sourceDataVec_8[11:10];
  wire [1:0]    maskDestinationResult_lo_67 = sourceDataVec_8[13:12];
  wire [1:0]    maskDestinationResult_hi_67 = sourceDataVec_8[15:14];
  wire [1:0]    maskDestinationResult_lo_68 = sourceDataVec_8[17:16];
  wire [1:0]    maskDestinationResult_hi_68 = sourceDataVec_8[19:18];
  wire [1:0]    maskDestinationResult_lo_69 = sourceDataVec_8[21:20];
  wire [1:0]    maskDestinationResult_hi_69 = sourceDataVec_8[23:22];
  wire [1:0]    maskDestinationResult_lo_70 = sourceDataVec_8[25:24];
  wire [1:0]    maskDestinationResult_hi_70 = sourceDataVec_8[27:26];
  wire [1:0]    maskDestinationResult_lo_71 = sourceDataVec_8[29:28];
  wire [1:0]    maskDestinationResult_hi_71 = sourceDataVec_8[31:30];
  wire [1:0]    maskDestinationResult_lo_72 = sourceDataVec_9[1:0];
  wire [1:0]    maskDestinationResult_hi_72 = sourceDataVec_9[3:2];
  wire [1:0]    maskDestinationResult_lo_73 = sourceDataVec_9[5:4];
  wire [1:0]    maskDestinationResult_hi_73 = sourceDataVec_9[7:6];
  wire [1:0]    maskDestinationResult_lo_74 = sourceDataVec_9[9:8];
  wire [1:0]    maskDestinationResult_hi_74 = sourceDataVec_9[11:10];
  wire [1:0]    maskDestinationResult_lo_75 = sourceDataVec_9[13:12];
  wire [1:0]    maskDestinationResult_hi_75 = sourceDataVec_9[15:14];
  wire [1:0]    maskDestinationResult_lo_76 = sourceDataVec_9[17:16];
  wire [1:0]    maskDestinationResult_hi_76 = sourceDataVec_9[19:18];
  wire [1:0]    maskDestinationResult_lo_77 = sourceDataVec_9[21:20];
  wire [1:0]    maskDestinationResult_hi_77 = sourceDataVec_9[23:22];
  wire [1:0]    maskDestinationResult_lo_78 = sourceDataVec_9[25:24];
  wire [1:0]    maskDestinationResult_hi_78 = sourceDataVec_9[27:26];
  wire [1:0]    maskDestinationResult_lo_79 = sourceDataVec_9[29:28];
  wire [1:0]    maskDestinationResult_hi_79 = sourceDataVec_9[31:30];
  wire [1:0]    maskDestinationResult_lo_80 = sourceDataVec_10[1:0];
  wire [1:0]    maskDestinationResult_hi_80 = sourceDataVec_10[3:2];
  wire [1:0]    maskDestinationResult_lo_81 = sourceDataVec_10[5:4];
  wire [1:0]    maskDestinationResult_hi_81 = sourceDataVec_10[7:6];
  wire [1:0]    maskDestinationResult_lo_82 = sourceDataVec_10[9:8];
  wire [1:0]    maskDestinationResult_hi_82 = sourceDataVec_10[11:10];
  wire [1:0]    maskDestinationResult_lo_83 = sourceDataVec_10[13:12];
  wire [1:0]    maskDestinationResult_hi_83 = sourceDataVec_10[15:14];
  wire [1:0]    maskDestinationResult_lo_84 = sourceDataVec_10[17:16];
  wire [1:0]    maskDestinationResult_hi_84 = sourceDataVec_10[19:18];
  wire [1:0]    maskDestinationResult_lo_85 = sourceDataVec_10[21:20];
  wire [1:0]    maskDestinationResult_hi_85 = sourceDataVec_10[23:22];
  wire [1:0]    maskDestinationResult_lo_86 = sourceDataVec_10[25:24];
  wire [1:0]    maskDestinationResult_hi_86 = sourceDataVec_10[27:26];
  wire [1:0]    maskDestinationResult_lo_87 = sourceDataVec_10[29:28];
  wire [1:0]    maskDestinationResult_hi_87 = sourceDataVec_10[31:30];
  wire [1:0]    maskDestinationResult_lo_88 = sourceDataVec_11[1:0];
  wire [1:0]    maskDestinationResult_hi_88 = sourceDataVec_11[3:2];
  wire [1:0]    maskDestinationResult_lo_89 = sourceDataVec_11[5:4];
  wire [1:0]    maskDestinationResult_hi_89 = sourceDataVec_11[7:6];
  wire [1:0]    maskDestinationResult_lo_90 = sourceDataVec_11[9:8];
  wire [1:0]    maskDestinationResult_hi_90 = sourceDataVec_11[11:10];
  wire [1:0]    maskDestinationResult_lo_91 = sourceDataVec_11[13:12];
  wire [1:0]    maskDestinationResult_hi_91 = sourceDataVec_11[15:14];
  wire [1:0]    maskDestinationResult_lo_92 = sourceDataVec_11[17:16];
  wire [1:0]    maskDestinationResult_hi_92 = sourceDataVec_11[19:18];
  wire [1:0]    maskDestinationResult_lo_93 = sourceDataVec_11[21:20];
  wire [1:0]    maskDestinationResult_hi_93 = sourceDataVec_11[23:22];
  wire [1:0]    maskDestinationResult_lo_94 = sourceDataVec_11[25:24];
  wire [1:0]    maskDestinationResult_hi_94 = sourceDataVec_11[27:26];
  wire [1:0]    maskDestinationResult_lo_95 = sourceDataVec_11[29:28];
  wire [1:0]    maskDestinationResult_hi_95 = sourceDataVec_11[31:30];
  wire [1:0]    maskDestinationResult_lo_96 = sourceDataVec_12[1:0];
  wire [1:0]    maskDestinationResult_hi_96 = sourceDataVec_12[3:2];
  wire [1:0]    maskDestinationResult_lo_97 = sourceDataVec_12[5:4];
  wire [1:0]    maskDestinationResult_hi_97 = sourceDataVec_12[7:6];
  wire [1:0]    maskDestinationResult_lo_98 = sourceDataVec_12[9:8];
  wire [1:0]    maskDestinationResult_hi_98 = sourceDataVec_12[11:10];
  wire [1:0]    maskDestinationResult_lo_99 = sourceDataVec_12[13:12];
  wire [1:0]    maskDestinationResult_hi_99 = sourceDataVec_12[15:14];
  wire [1:0]    maskDestinationResult_lo_100 = sourceDataVec_12[17:16];
  wire [1:0]    maskDestinationResult_hi_100 = sourceDataVec_12[19:18];
  wire [1:0]    maskDestinationResult_lo_101 = sourceDataVec_12[21:20];
  wire [1:0]    maskDestinationResult_hi_101 = sourceDataVec_12[23:22];
  wire [1:0]    maskDestinationResult_lo_102 = sourceDataVec_12[25:24];
  wire [1:0]    maskDestinationResult_hi_102 = sourceDataVec_12[27:26];
  wire [1:0]    maskDestinationResult_lo_103 = sourceDataVec_12[29:28];
  wire [1:0]    maskDestinationResult_hi_103 = sourceDataVec_12[31:30];
  wire [1:0]    maskDestinationResult_lo_104 = sourceDataVec_13[1:0];
  wire [1:0]    maskDestinationResult_hi_104 = sourceDataVec_13[3:2];
  wire [1:0]    maskDestinationResult_lo_105 = sourceDataVec_13[5:4];
  wire [1:0]    maskDestinationResult_hi_105 = sourceDataVec_13[7:6];
  wire [1:0]    maskDestinationResult_lo_106 = sourceDataVec_13[9:8];
  wire [1:0]    maskDestinationResult_hi_106 = sourceDataVec_13[11:10];
  wire [1:0]    maskDestinationResult_lo_107 = sourceDataVec_13[13:12];
  wire [1:0]    maskDestinationResult_hi_107 = sourceDataVec_13[15:14];
  wire [1:0]    maskDestinationResult_lo_108 = sourceDataVec_13[17:16];
  wire [1:0]    maskDestinationResult_hi_108 = sourceDataVec_13[19:18];
  wire [1:0]    maskDestinationResult_lo_109 = sourceDataVec_13[21:20];
  wire [1:0]    maskDestinationResult_hi_109 = sourceDataVec_13[23:22];
  wire [1:0]    maskDestinationResult_lo_110 = sourceDataVec_13[25:24];
  wire [1:0]    maskDestinationResult_hi_110 = sourceDataVec_13[27:26];
  wire [1:0]    maskDestinationResult_lo_111 = sourceDataVec_13[29:28];
  wire [1:0]    maskDestinationResult_hi_111 = sourceDataVec_13[31:30];
  wire [1:0]    maskDestinationResult_lo_112 = sourceDataVec_14[1:0];
  wire [1:0]    maskDestinationResult_hi_112 = sourceDataVec_14[3:2];
  wire [1:0]    maskDestinationResult_lo_113 = sourceDataVec_14[5:4];
  wire [1:0]    maskDestinationResult_hi_113 = sourceDataVec_14[7:6];
  wire [1:0]    maskDestinationResult_lo_114 = sourceDataVec_14[9:8];
  wire [1:0]    maskDestinationResult_hi_114 = sourceDataVec_14[11:10];
  wire [1:0]    maskDestinationResult_lo_115 = sourceDataVec_14[13:12];
  wire [1:0]    maskDestinationResult_hi_115 = sourceDataVec_14[15:14];
  wire [1:0]    maskDestinationResult_lo_116 = sourceDataVec_14[17:16];
  wire [1:0]    maskDestinationResult_hi_116 = sourceDataVec_14[19:18];
  wire [1:0]    maskDestinationResult_lo_117 = sourceDataVec_14[21:20];
  wire [1:0]    maskDestinationResult_hi_117 = sourceDataVec_14[23:22];
  wire [1:0]    maskDestinationResult_lo_118 = sourceDataVec_14[25:24];
  wire [1:0]    maskDestinationResult_hi_118 = sourceDataVec_14[27:26];
  wire [1:0]    maskDestinationResult_lo_119 = sourceDataVec_14[29:28];
  wire [1:0]    maskDestinationResult_hi_119 = sourceDataVec_14[31:30];
  wire [1:0]    maskDestinationResult_lo_120 = sourceDataVec_15[1:0];
  wire [1:0]    maskDestinationResult_hi_120 = sourceDataVec_15[3:2];
  wire [1:0]    maskDestinationResult_lo_121 = sourceDataVec_15[5:4];
  wire [1:0]    maskDestinationResult_hi_121 = sourceDataVec_15[7:6];
  wire [1:0]    maskDestinationResult_lo_122 = sourceDataVec_15[9:8];
  wire [1:0]    maskDestinationResult_hi_122 = sourceDataVec_15[11:10];
  wire [1:0]    maskDestinationResult_lo_123 = sourceDataVec_15[13:12];
  wire [1:0]    maskDestinationResult_hi_123 = sourceDataVec_15[15:14];
  wire [1:0]    maskDestinationResult_lo_124 = sourceDataVec_15[17:16];
  wire [1:0]    maskDestinationResult_hi_124 = sourceDataVec_15[19:18];
  wire [1:0]    maskDestinationResult_lo_125 = sourceDataVec_15[21:20];
  wire [1:0]    maskDestinationResult_hi_125 = sourceDataVec_15[23:22];
  wire [1:0]    maskDestinationResult_lo_126 = sourceDataVec_15[25:24];
  wire [1:0]    maskDestinationResult_hi_126 = sourceDataVec_15[27:26];
  wire [1:0]    maskDestinationResult_lo_127 = sourceDataVec_15[29:28];
  wire [1:0]    maskDestinationResult_hi_127 = sourceDataVec_15[31:30];
  wire [1:0]    maskDestinationResult_lo_128 = sourceDataVec_16[1:0];
  wire [1:0]    maskDestinationResult_hi_128 = sourceDataVec_16[3:2];
  wire [1:0]    maskDestinationResult_lo_129 = sourceDataVec_16[5:4];
  wire [1:0]    maskDestinationResult_hi_129 = sourceDataVec_16[7:6];
  wire [1:0]    maskDestinationResult_lo_130 = sourceDataVec_16[9:8];
  wire [1:0]    maskDestinationResult_hi_130 = sourceDataVec_16[11:10];
  wire [1:0]    maskDestinationResult_lo_131 = sourceDataVec_16[13:12];
  wire [1:0]    maskDestinationResult_hi_131 = sourceDataVec_16[15:14];
  wire [1:0]    maskDestinationResult_lo_132 = sourceDataVec_16[17:16];
  wire [1:0]    maskDestinationResult_hi_132 = sourceDataVec_16[19:18];
  wire [1:0]    maskDestinationResult_lo_133 = sourceDataVec_16[21:20];
  wire [1:0]    maskDestinationResult_hi_133 = sourceDataVec_16[23:22];
  wire [1:0]    maskDestinationResult_lo_134 = sourceDataVec_16[25:24];
  wire [1:0]    maskDestinationResult_hi_134 = sourceDataVec_16[27:26];
  wire [1:0]    maskDestinationResult_lo_135 = sourceDataVec_16[29:28];
  wire [1:0]    maskDestinationResult_hi_135 = sourceDataVec_16[31:30];
  wire [1:0]    maskDestinationResult_lo_136 = sourceDataVec_17[1:0];
  wire [1:0]    maskDestinationResult_hi_136 = sourceDataVec_17[3:2];
  wire [1:0]    maskDestinationResult_lo_137 = sourceDataVec_17[5:4];
  wire [1:0]    maskDestinationResult_hi_137 = sourceDataVec_17[7:6];
  wire [1:0]    maskDestinationResult_lo_138 = sourceDataVec_17[9:8];
  wire [1:0]    maskDestinationResult_hi_138 = sourceDataVec_17[11:10];
  wire [1:0]    maskDestinationResult_lo_139 = sourceDataVec_17[13:12];
  wire [1:0]    maskDestinationResult_hi_139 = sourceDataVec_17[15:14];
  wire [1:0]    maskDestinationResult_lo_140 = sourceDataVec_17[17:16];
  wire [1:0]    maskDestinationResult_hi_140 = sourceDataVec_17[19:18];
  wire [1:0]    maskDestinationResult_lo_141 = sourceDataVec_17[21:20];
  wire [1:0]    maskDestinationResult_hi_141 = sourceDataVec_17[23:22];
  wire [1:0]    maskDestinationResult_lo_142 = sourceDataVec_17[25:24];
  wire [1:0]    maskDestinationResult_hi_142 = sourceDataVec_17[27:26];
  wire [1:0]    maskDestinationResult_lo_143 = sourceDataVec_17[29:28];
  wire [1:0]    maskDestinationResult_hi_143 = sourceDataVec_17[31:30];
  wire [1:0]    maskDestinationResult_lo_144 = sourceDataVec_18[1:0];
  wire [1:0]    maskDestinationResult_hi_144 = sourceDataVec_18[3:2];
  wire [1:0]    maskDestinationResult_lo_145 = sourceDataVec_18[5:4];
  wire [1:0]    maskDestinationResult_hi_145 = sourceDataVec_18[7:6];
  wire [1:0]    maskDestinationResult_lo_146 = sourceDataVec_18[9:8];
  wire [1:0]    maskDestinationResult_hi_146 = sourceDataVec_18[11:10];
  wire [1:0]    maskDestinationResult_lo_147 = sourceDataVec_18[13:12];
  wire [1:0]    maskDestinationResult_hi_147 = sourceDataVec_18[15:14];
  wire [1:0]    maskDestinationResult_lo_148 = sourceDataVec_18[17:16];
  wire [1:0]    maskDestinationResult_hi_148 = sourceDataVec_18[19:18];
  wire [1:0]    maskDestinationResult_lo_149 = sourceDataVec_18[21:20];
  wire [1:0]    maskDestinationResult_hi_149 = sourceDataVec_18[23:22];
  wire [1:0]    maskDestinationResult_lo_150 = sourceDataVec_18[25:24];
  wire [1:0]    maskDestinationResult_hi_150 = sourceDataVec_18[27:26];
  wire [1:0]    maskDestinationResult_lo_151 = sourceDataVec_18[29:28];
  wire [1:0]    maskDestinationResult_hi_151 = sourceDataVec_18[31:30];
  wire [1:0]    maskDestinationResult_lo_152 = sourceDataVec_19[1:0];
  wire [1:0]    maskDestinationResult_hi_152 = sourceDataVec_19[3:2];
  wire [1:0]    maskDestinationResult_lo_153 = sourceDataVec_19[5:4];
  wire [1:0]    maskDestinationResult_hi_153 = sourceDataVec_19[7:6];
  wire [1:0]    maskDestinationResult_lo_154 = sourceDataVec_19[9:8];
  wire [1:0]    maskDestinationResult_hi_154 = sourceDataVec_19[11:10];
  wire [1:0]    maskDestinationResult_lo_155 = sourceDataVec_19[13:12];
  wire [1:0]    maskDestinationResult_hi_155 = sourceDataVec_19[15:14];
  wire [1:0]    maskDestinationResult_lo_156 = sourceDataVec_19[17:16];
  wire [1:0]    maskDestinationResult_hi_156 = sourceDataVec_19[19:18];
  wire [1:0]    maskDestinationResult_lo_157 = sourceDataVec_19[21:20];
  wire [1:0]    maskDestinationResult_hi_157 = sourceDataVec_19[23:22];
  wire [1:0]    maskDestinationResult_lo_158 = sourceDataVec_19[25:24];
  wire [1:0]    maskDestinationResult_hi_158 = sourceDataVec_19[27:26];
  wire [1:0]    maskDestinationResult_lo_159 = sourceDataVec_19[29:28];
  wire [1:0]    maskDestinationResult_hi_159 = sourceDataVec_19[31:30];
  wire [1:0]    maskDestinationResult_lo_160 = sourceDataVec_20[1:0];
  wire [1:0]    maskDestinationResult_hi_160 = sourceDataVec_20[3:2];
  wire [1:0]    maskDestinationResult_lo_161 = sourceDataVec_20[5:4];
  wire [1:0]    maskDestinationResult_hi_161 = sourceDataVec_20[7:6];
  wire [1:0]    maskDestinationResult_lo_162 = sourceDataVec_20[9:8];
  wire [1:0]    maskDestinationResult_hi_162 = sourceDataVec_20[11:10];
  wire [1:0]    maskDestinationResult_lo_163 = sourceDataVec_20[13:12];
  wire [1:0]    maskDestinationResult_hi_163 = sourceDataVec_20[15:14];
  wire [1:0]    maskDestinationResult_lo_164 = sourceDataVec_20[17:16];
  wire [1:0]    maskDestinationResult_hi_164 = sourceDataVec_20[19:18];
  wire [1:0]    maskDestinationResult_lo_165 = sourceDataVec_20[21:20];
  wire [1:0]    maskDestinationResult_hi_165 = sourceDataVec_20[23:22];
  wire [1:0]    maskDestinationResult_lo_166 = sourceDataVec_20[25:24];
  wire [1:0]    maskDestinationResult_hi_166 = sourceDataVec_20[27:26];
  wire [1:0]    maskDestinationResult_lo_167 = sourceDataVec_20[29:28];
  wire [1:0]    maskDestinationResult_hi_167 = sourceDataVec_20[31:30];
  wire [1:0]    maskDestinationResult_lo_168 = sourceDataVec_21[1:0];
  wire [1:0]    maskDestinationResult_hi_168 = sourceDataVec_21[3:2];
  wire [1:0]    maskDestinationResult_lo_169 = sourceDataVec_21[5:4];
  wire [1:0]    maskDestinationResult_hi_169 = sourceDataVec_21[7:6];
  wire [1:0]    maskDestinationResult_lo_170 = sourceDataVec_21[9:8];
  wire [1:0]    maskDestinationResult_hi_170 = sourceDataVec_21[11:10];
  wire [1:0]    maskDestinationResult_lo_171 = sourceDataVec_21[13:12];
  wire [1:0]    maskDestinationResult_hi_171 = sourceDataVec_21[15:14];
  wire [1:0]    maskDestinationResult_lo_172 = sourceDataVec_21[17:16];
  wire [1:0]    maskDestinationResult_hi_172 = sourceDataVec_21[19:18];
  wire [1:0]    maskDestinationResult_lo_173 = sourceDataVec_21[21:20];
  wire [1:0]    maskDestinationResult_hi_173 = sourceDataVec_21[23:22];
  wire [1:0]    maskDestinationResult_lo_174 = sourceDataVec_21[25:24];
  wire [1:0]    maskDestinationResult_hi_174 = sourceDataVec_21[27:26];
  wire [1:0]    maskDestinationResult_lo_175 = sourceDataVec_21[29:28];
  wire [1:0]    maskDestinationResult_hi_175 = sourceDataVec_21[31:30];
  wire [1:0]    maskDestinationResult_lo_176 = sourceDataVec_22[1:0];
  wire [1:0]    maskDestinationResult_hi_176 = sourceDataVec_22[3:2];
  wire [1:0]    maskDestinationResult_lo_177 = sourceDataVec_22[5:4];
  wire [1:0]    maskDestinationResult_hi_177 = sourceDataVec_22[7:6];
  wire [1:0]    maskDestinationResult_lo_178 = sourceDataVec_22[9:8];
  wire [1:0]    maskDestinationResult_hi_178 = sourceDataVec_22[11:10];
  wire [1:0]    maskDestinationResult_lo_179 = sourceDataVec_22[13:12];
  wire [1:0]    maskDestinationResult_hi_179 = sourceDataVec_22[15:14];
  wire [1:0]    maskDestinationResult_lo_180 = sourceDataVec_22[17:16];
  wire [1:0]    maskDestinationResult_hi_180 = sourceDataVec_22[19:18];
  wire [1:0]    maskDestinationResult_lo_181 = sourceDataVec_22[21:20];
  wire [1:0]    maskDestinationResult_hi_181 = sourceDataVec_22[23:22];
  wire [1:0]    maskDestinationResult_lo_182 = sourceDataVec_22[25:24];
  wire [1:0]    maskDestinationResult_hi_182 = sourceDataVec_22[27:26];
  wire [1:0]    maskDestinationResult_lo_183 = sourceDataVec_22[29:28];
  wire [1:0]    maskDestinationResult_hi_183 = sourceDataVec_22[31:30];
  wire [1:0]    maskDestinationResult_lo_184 = sourceDataVec_23[1:0];
  wire [1:0]    maskDestinationResult_hi_184 = sourceDataVec_23[3:2];
  wire [1:0]    maskDestinationResult_lo_185 = sourceDataVec_23[5:4];
  wire [1:0]    maskDestinationResult_hi_185 = sourceDataVec_23[7:6];
  wire [1:0]    maskDestinationResult_lo_186 = sourceDataVec_23[9:8];
  wire [1:0]    maskDestinationResult_hi_186 = sourceDataVec_23[11:10];
  wire [1:0]    maskDestinationResult_lo_187 = sourceDataVec_23[13:12];
  wire [1:0]    maskDestinationResult_hi_187 = sourceDataVec_23[15:14];
  wire [1:0]    maskDestinationResult_lo_188 = sourceDataVec_23[17:16];
  wire [1:0]    maskDestinationResult_hi_188 = sourceDataVec_23[19:18];
  wire [1:0]    maskDestinationResult_lo_189 = sourceDataVec_23[21:20];
  wire [1:0]    maskDestinationResult_hi_189 = sourceDataVec_23[23:22];
  wire [1:0]    maskDestinationResult_lo_190 = sourceDataVec_23[25:24];
  wire [1:0]    maskDestinationResult_hi_190 = sourceDataVec_23[27:26];
  wire [1:0]    maskDestinationResult_lo_191 = sourceDataVec_23[29:28];
  wire [1:0]    maskDestinationResult_hi_191 = sourceDataVec_23[31:30];
  wire [1:0]    maskDestinationResult_lo_192 = sourceDataVec_24[1:0];
  wire [1:0]    maskDestinationResult_hi_192 = sourceDataVec_24[3:2];
  wire [1:0]    maskDestinationResult_lo_193 = sourceDataVec_24[5:4];
  wire [1:0]    maskDestinationResult_hi_193 = sourceDataVec_24[7:6];
  wire [1:0]    maskDestinationResult_lo_194 = sourceDataVec_24[9:8];
  wire [1:0]    maskDestinationResult_hi_194 = sourceDataVec_24[11:10];
  wire [1:0]    maskDestinationResult_lo_195 = sourceDataVec_24[13:12];
  wire [1:0]    maskDestinationResult_hi_195 = sourceDataVec_24[15:14];
  wire [1:0]    maskDestinationResult_lo_196 = sourceDataVec_24[17:16];
  wire [1:0]    maskDestinationResult_hi_196 = sourceDataVec_24[19:18];
  wire [1:0]    maskDestinationResult_lo_197 = sourceDataVec_24[21:20];
  wire [1:0]    maskDestinationResult_hi_197 = sourceDataVec_24[23:22];
  wire [1:0]    maskDestinationResult_lo_198 = sourceDataVec_24[25:24];
  wire [1:0]    maskDestinationResult_hi_198 = sourceDataVec_24[27:26];
  wire [1:0]    maskDestinationResult_lo_199 = sourceDataVec_24[29:28];
  wire [1:0]    maskDestinationResult_hi_199 = sourceDataVec_24[31:30];
  wire [1:0]    maskDestinationResult_lo_200 = sourceDataVec_25[1:0];
  wire [1:0]    maskDestinationResult_hi_200 = sourceDataVec_25[3:2];
  wire [1:0]    maskDestinationResult_lo_201 = sourceDataVec_25[5:4];
  wire [1:0]    maskDestinationResult_hi_201 = sourceDataVec_25[7:6];
  wire [1:0]    maskDestinationResult_lo_202 = sourceDataVec_25[9:8];
  wire [1:0]    maskDestinationResult_hi_202 = sourceDataVec_25[11:10];
  wire [1:0]    maskDestinationResult_lo_203 = sourceDataVec_25[13:12];
  wire [1:0]    maskDestinationResult_hi_203 = sourceDataVec_25[15:14];
  wire [1:0]    maskDestinationResult_lo_204 = sourceDataVec_25[17:16];
  wire [1:0]    maskDestinationResult_hi_204 = sourceDataVec_25[19:18];
  wire [1:0]    maskDestinationResult_lo_205 = sourceDataVec_25[21:20];
  wire [1:0]    maskDestinationResult_hi_205 = sourceDataVec_25[23:22];
  wire [1:0]    maskDestinationResult_lo_206 = sourceDataVec_25[25:24];
  wire [1:0]    maskDestinationResult_hi_206 = sourceDataVec_25[27:26];
  wire [1:0]    maskDestinationResult_lo_207 = sourceDataVec_25[29:28];
  wire [1:0]    maskDestinationResult_hi_207 = sourceDataVec_25[31:30];
  wire [1:0]    maskDestinationResult_lo_208 = sourceDataVec_26[1:0];
  wire [1:0]    maskDestinationResult_hi_208 = sourceDataVec_26[3:2];
  wire [1:0]    maskDestinationResult_lo_209 = sourceDataVec_26[5:4];
  wire [1:0]    maskDestinationResult_hi_209 = sourceDataVec_26[7:6];
  wire [1:0]    maskDestinationResult_lo_210 = sourceDataVec_26[9:8];
  wire [1:0]    maskDestinationResult_hi_210 = sourceDataVec_26[11:10];
  wire [1:0]    maskDestinationResult_lo_211 = sourceDataVec_26[13:12];
  wire [1:0]    maskDestinationResult_hi_211 = sourceDataVec_26[15:14];
  wire [1:0]    maskDestinationResult_lo_212 = sourceDataVec_26[17:16];
  wire [1:0]    maskDestinationResult_hi_212 = sourceDataVec_26[19:18];
  wire [1:0]    maskDestinationResult_lo_213 = sourceDataVec_26[21:20];
  wire [1:0]    maskDestinationResult_hi_213 = sourceDataVec_26[23:22];
  wire [1:0]    maskDestinationResult_lo_214 = sourceDataVec_26[25:24];
  wire [1:0]    maskDestinationResult_hi_214 = sourceDataVec_26[27:26];
  wire [1:0]    maskDestinationResult_lo_215 = sourceDataVec_26[29:28];
  wire [1:0]    maskDestinationResult_hi_215 = sourceDataVec_26[31:30];
  wire [1:0]    maskDestinationResult_lo_216 = sourceDataVec_27[1:0];
  wire [1:0]    maskDestinationResult_hi_216 = sourceDataVec_27[3:2];
  wire [1:0]    maskDestinationResult_lo_217 = sourceDataVec_27[5:4];
  wire [1:0]    maskDestinationResult_hi_217 = sourceDataVec_27[7:6];
  wire [1:0]    maskDestinationResult_lo_218 = sourceDataVec_27[9:8];
  wire [1:0]    maskDestinationResult_hi_218 = sourceDataVec_27[11:10];
  wire [1:0]    maskDestinationResult_lo_219 = sourceDataVec_27[13:12];
  wire [1:0]    maskDestinationResult_hi_219 = sourceDataVec_27[15:14];
  wire [1:0]    maskDestinationResult_lo_220 = sourceDataVec_27[17:16];
  wire [1:0]    maskDestinationResult_hi_220 = sourceDataVec_27[19:18];
  wire [1:0]    maskDestinationResult_lo_221 = sourceDataVec_27[21:20];
  wire [1:0]    maskDestinationResult_hi_221 = sourceDataVec_27[23:22];
  wire [1:0]    maskDestinationResult_lo_222 = sourceDataVec_27[25:24];
  wire [1:0]    maskDestinationResult_hi_222 = sourceDataVec_27[27:26];
  wire [1:0]    maskDestinationResult_lo_223 = sourceDataVec_27[29:28];
  wire [1:0]    maskDestinationResult_hi_223 = sourceDataVec_27[31:30];
  wire [1:0]    maskDestinationResult_lo_224 = sourceDataVec_28[1:0];
  wire [1:0]    maskDestinationResult_hi_224 = sourceDataVec_28[3:2];
  wire [1:0]    maskDestinationResult_lo_225 = sourceDataVec_28[5:4];
  wire [1:0]    maskDestinationResult_hi_225 = sourceDataVec_28[7:6];
  wire [1:0]    maskDestinationResult_lo_226 = sourceDataVec_28[9:8];
  wire [1:0]    maskDestinationResult_hi_226 = sourceDataVec_28[11:10];
  wire [1:0]    maskDestinationResult_lo_227 = sourceDataVec_28[13:12];
  wire [1:0]    maskDestinationResult_hi_227 = sourceDataVec_28[15:14];
  wire [1:0]    maskDestinationResult_lo_228 = sourceDataVec_28[17:16];
  wire [1:0]    maskDestinationResult_hi_228 = sourceDataVec_28[19:18];
  wire [1:0]    maskDestinationResult_lo_229 = sourceDataVec_28[21:20];
  wire [1:0]    maskDestinationResult_hi_229 = sourceDataVec_28[23:22];
  wire [1:0]    maskDestinationResult_lo_230 = sourceDataVec_28[25:24];
  wire [1:0]    maskDestinationResult_hi_230 = sourceDataVec_28[27:26];
  wire [1:0]    maskDestinationResult_lo_231 = sourceDataVec_28[29:28];
  wire [1:0]    maskDestinationResult_hi_231 = sourceDataVec_28[31:30];
  wire [1:0]    maskDestinationResult_lo_232 = sourceDataVec_29[1:0];
  wire [1:0]    maskDestinationResult_hi_232 = sourceDataVec_29[3:2];
  wire [1:0]    maskDestinationResult_lo_233 = sourceDataVec_29[5:4];
  wire [1:0]    maskDestinationResult_hi_233 = sourceDataVec_29[7:6];
  wire [1:0]    maskDestinationResult_lo_234 = sourceDataVec_29[9:8];
  wire [1:0]    maskDestinationResult_hi_234 = sourceDataVec_29[11:10];
  wire [1:0]    maskDestinationResult_lo_235 = sourceDataVec_29[13:12];
  wire [1:0]    maskDestinationResult_hi_235 = sourceDataVec_29[15:14];
  wire [1:0]    maskDestinationResult_lo_236 = sourceDataVec_29[17:16];
  wire [1:0]    maskDestinationResult_hi_236 = sourceDataVec_29[19:18];
  wire [1:0]    maskDestinationResult_lo_237 = sourceDataVec_29[21:20];
  wire [1:0]    maskDestinationResult_hi_237 = sourceDataVec_29[23:22];
  wire [1:0]    maskDestinationResult_lo_238 = sourceDataVec_29[25:24];
  wire [1:0]    maskDestinationResult_hi_238 = sourceDataVec_29[27:26];
  wire [1:0]    maskDestinationResult_lo_239 = sourceDataVec_29[29:28];
  wire [1:0]    maskDestinationResult_hi_239 = sourceDataVec_29[31:30];
  wire [1:0]    maskDestinationResult_lo_240 = sourceDataVec_30[1:0];
  wire [1:0]    maskDestinationResult_hi_240 = sourceDataVec_30[3:2];
  wire [1:0]    maskDestinationResult_lo_241 = sourceDataVec_30[5:4];
  wire [1:0]    maskDestinationResult_hi_241 = sourceDataVec_30[7:6];
  wire [1:0]    maskDestinationResult_lo_242 = sourceDataVec_30[9:8];
  wire [1:0]    maskDestinationResult_hi_242 = sourceDataVec_30[11:10];
  wire [1:0]    maskDestinationResult_lo_243 = sourceDataVec_30[13:12];
  wire [1:0]    maskDestinationResult_hi_243 = sourceDataVec_30[15:14];
  wire [1:0]    maskDestinationResult_lo_244 = sourceDataVec_30[17:16];
  wire [1:0]    maskDestinationResult_hi_244 = sourceDataVec_30[19:18];
  wire [1:0]    maskDestinationResult_lo_245 = sourceDataVec_30[21:20];
  wire [1:0]    maskDestinationResult_hi_245 = sourceDataVec_30[23:22];
  wire [1:0]    maskDestinationResult_lo_246 = sourceDataVec_30[25:24];
  wire [1:0]    maskDestinationResult_hi_246 = sourceDataVec_30[27:26];
  wire [1:0]    maskDestinationResult_lo_247 = sourceDataVec_30[29:28];
  wire [1:0]    maskDestinationResult_hi_247 = sourceDataVec_30[31:30];
  wire [1:0]    maskDestinationResult_lo_248 = sourceDataVec_31[1:0];
  wire [1:0]    maskDestinationResult_hi_248 = sourceDataVec_31[3:2];
  wire [1:0]    maskDestinationResult_lo_249 = sourceDataVec_31[5:4];
  wire [1:0]    maskDestinationResult_hi_249 = sourceDataVec_31[7:6];
  wire [1:0]    maskDestinationResult_lo_250 = sourceDataVec_31[9:8];
  wire [1:0]    maskDestinationResult_hi_250 = sourceDataVec_31[11:10];
  wire [1:0]    maskDestinationResult_lo_251 = sourceDataVec_31[13:12];
  wire [1:0]    maskDestinationResult_hi_251 = sourceDataVec_31[15:14];
  wire [1:0]    maskDestinationResult_lo_252 = sourceDataVec_31[17:16];
  wire [1:0]    maskDestinationResult_hi_252 = sourceDataVec_31[19:18];
  wire [1:0]    maskDestinationResult_lo_253 = sourceDataVec_31[21:20];
  wire [1:0]    maskDestinationResult_hi_253 = sourceDataVec_31[23:22];
  wire [1:0]    maskDestinationResult_lo_254 = sourceDataVec_31[25:24];
  wire [1:0]    maskDestinationResult_hi_254 = sourceDataVec_31[27:26];
  wire [1:0]    maskDestinationResult_lo_255 = sourceDataVec_31[29:28];
  wire [1:0]    maskDestinationResult_hi_255 = sourceDataVec_31[31:30];
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo = {maskDestinationResult_hi_8, maskDestinationResult_lo_8, maskDestinationResult_hi, maskDestinationResult_lo};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi = {maskDestinationResult_hi_24, maskDestinationResult_lo_24, maskDestinationResult_hi_16, maskDestinationResult_lo_16};
  wire [15:0]   maskDestinationResult_lo_lo_lo = {maskDestinationResult_lo_lo_lo_hi, maskDestinationResult_lo_lo_lo_lo};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo = {maskDestinationResult_hi_40, maskDestinationResult_lo_40, maskDestinationResult_hi_32, maskDestinationResult_lo_32};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi = {maskDestinationResult_hi_56, maskDestinationResult_lo_56, maskDestinationResult_hi_48, maskDestinationResult_lo_48};
  wire [15:0]   maskDestinationResult_lo_lo_hi = {maskDestinationResult_lo_lo_hi_hi, maskDestinationResult_lo_lo_hi_lo};
  wire [31:0]   maskDestinationResult_lo_lo = {maskDestinationResult_lo_lo_hi, maskDestinationResult_lo_lo_lo};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo = {maskDestinationResult_hi_72, maskDestinationResult_lo_72, maskDestinationResult_hi_64, maskDestinationResult_lo_64};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi = {maskDestinationResult_hi_88, maskDestinationResult_lo_88, maskDestinationResult_hi_80, maskDestinationResult_lo_80};
  wire [15:0]   maskDestinationResult_lo_hi_lo = {maskDestinationResult_lo_hi_lo_hi, maskDestinationResult_lo_hi_lo_lo};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo = {maskDestinationResult_hi_104, maskDestinationResult_lo_104, maskDestinationResult_hi_96, maskDestinationResult_lo_96};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi = {maskDestinationResult_hi_120, maskDestinationResult_lo_120, maskDestinationResult_hi_112, maskDestinationResult_lo_112};
  wire [15:0]   maskDestinationResult_lo_hi_hi = {maskDestinationResult_lo_hi_hi_hi, maskDestinationResult_lo_hi_hi_lo};
  wire [31:0]   maskDestinationResult_lo_hi = {maskDestinationResult_lo_hi_hi, maskDestinationResult_lo_hi_lo};
  wire [63:0]   maskDestinationResult_lo_256 = {maskDestinationResult_lo_hi, maskDestinationResult_lo_lo};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo = {maskDestinationResult_hi_136, maskDestinationResult_lo_136, maskDestinationResult_hi_128, maskDestinationResult_lo_128};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi = {maskDestinationResult_hi_152, maskDestinationResult_lo_152, maskDestinationResult_hi_144, maskDestinationResult_lo_144};
  wire [15:0]   maskDestinationResult_hi_lo_lo = {maskDestinationResult_hi_lo_lo_hi, maskDestinationResult_hi_lo_lo_lo};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo = {maskDestinationResult_hi_168, maskDestinationResult_lo_168, maskDestinationResult_hi_160, maskDestinationResult_lo_160};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi = {maskDestinationResult_hi_184, maskDestinationResult_lo_184, maskDestinationResult_hi_176, maskDestinationResult_lo_176};
  wire [15:0]   maskDestinationResult_hi_lo_hi = {maskDestinationResult_hi_lo_hi_hi, maskDestinationResult_hi_lo_hi_lo};
  wire [31:0]   maskDestinationResult_hi_lo = {maskDestinationResult_hi_lo_hi, maskDestinationResult_hi_lo_lo};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo = {maskDestinationResult_hi_200, maskDestinationResult_lo_200, maskDestinationResult_hi_192, maskDestinationResult_lo_192};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi = {maskDestinationResult_hi_216, maskDestinationResult_lo_216, maskDestinationResult_hi_208, maskDestinationResult_lo_208};
  wire [15:0]   maskDestinationResult_hi_hi_lo = {maskDestinationResult_hi_hi_lo_hi, maskDestinationResult_hi_hi_lo_lo};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo = {maskDestinationResult_hi_232, maskDestinationResult_lo_232, maskDestinationResult_hi_224, maskDestinationResult_lo_224};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi = {maskDestinationResult_hi_248, maskDestinationResult_lo_248, maskDestinationResult_hi_240, maskDestinationResult_lo_240};
  wire [15:0]   maskDestinationResult_hi_hi_hi = {maskDestinationResult_hi_hi_hi_hi, maskDestinationResult_hi_hi_hi_lo};
  wire [31:0]   maskDestinationResult_hi_hi = {maskDestinationResult_hi_hi_hi, maskDestinationResult_hi_hi_lo};
  wire [63:0]   maskDestinationResult_hi_256 = {maskDestinationResult_hi_hi, maskDestinationResult_hi_lo};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_1 = {maskDestinationResult_hi_9, maskDestinationResult_lo_9, maskDestinationResult_hi_1, maskDestinationResult_lo_1};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_1 = {maskDestinationResult_hi_25, maskDestinationResult_lo_25, maskDestinationResult_hi_17, maskDestinationResult_lo_17};
  wire [15:0]   maskDestinationResult_lo_lo_lo_1 = {maskDestinationResult_lo_lo_lo_hi_1, maskDestinationResult_lo_lo_lo_lo_1};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_1 = {maskDestinationResult_hi_41, maskDestinationResult_lo_41, maskDestinationResult_hi_33, maskDestinationResult_lo_33};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_1 = {maskDestinationResult_hi_57, maskDestinationResult_lo_57, maskDestinationResult_hi_49, maskDestinationResult_lo_49};
  wire [15:0]   maskDestinationResult_lo_lo_hi_1 = {maskDestinationResult_lo_lo_hi_hi_1, maskDestinationResult_lo_lo_hi_lo_1};
  wire [31:0]   maskDestinationResult_lo_lo_1 = {maskDestinationResult_lo_lo_hi_1, maskDestinationResult_lo_lo_lo_1};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_1 = {maskDestinationResult_hi_73, maskDestinationResult_lo_73, maskDestinationResult_hi_65, maskDestinationResult_lo_65};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_1 = {maskDestinationResult_hi_89, maskDestinationResult_lo_89, maskDestinationResult_hi_81, maskDestinationResult_lo_81};
  wire [15:0]   maskDestinationResult_lo_hi_lo_1 = {maskDestinationResult_lo_hi_lo_hi_1, maskDestinationResult_lo_hi_lo_lo_1};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_1 = {maskDestinationResult_hi_105, maskDestinationResult_lo_105, maskDestinationResult_hi_97, maskDestinationResult_lo_97};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_1 = {maskDestinationResult_hi_121, maskDestinationResult_lo_121, maskDestinationResult_hi_113, maskDestinationResult_lo_113};
  wire [15:0]   maskDestinationResult_lo_hi_hi_1 = {maskDestinationResult_lo_hi_hi_hi_1, maskDestinationResult_lo_hi_hi_lo_1};
  wire [31:0]   maskDestinationResult_lo_hi_1 = {maskDestinationResult_lo_hi_hi_1, maskDestinationResult_lo_hi_lo_1};
  wire [63:0]   maskDestinationResult_lo_257 = {maskDestinationResult_lo_hi_1, maskDestinationResult_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_1 = {maskDestinationResult_hi_137, maskDestinationResult_lo_137, maskDestinationResult_hi_129, maskDestinationResult_lo_129};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_1 = {maskDestinationResult_hi_153, maskDestinationResult_lo_153, maskDestinationResult_hi_145, maskDestinationResult_lo_145};
  wire [15:0]   maskDestinationResult_hi_lo_lo_1 = {maskDestinationResult_hi_lo_lo_hi_1, maskDestinationResult_hi_lo_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_1 = {maskDestinationResult_hi_169, maskDestinationResult_lo_169, maskDestinationResult_hi_161, maskDestinationResult_lo_161};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_1 = {maskDestinationResult_hi_185, maskDestinationResult_lo_185, maskDestinationResult_hi_177, maskDestinationResult_lo_177};
  wire [15:0]   maskDestinationResult_hi_lo_hi_1 = {maskDestinationResult_hi_lo_hi_hi_1, maskDestinationResult_hi_lo_hi_lo_1};
  wire [31:0]   maskDestinationResult_hi_lo_1 = {maskDestinationResult_hi_lo_hi_1, maskDestinationResult_hi_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_1 = {maskDestinationResult_hi_201, maskDestinationResult_lo_201, maskDestinationResult_hi_193, maskDestinationResult_lo_193};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_1 = {maskDestinationResult_hi_217, maskDestinationResult_lo_217, maskDestinationResult_hi_209, maskDestinationResult_lo_209};
  wire [15:0]   maskDestinationResult_hi_hi_lo_1 = {maskDestinationResult_hi_hi_lo_hi_1, maskDestinationResult_hi_hi_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_1 = {maskDestinationResult_hi_233, maskDestinationResult_lo_233, maskDestinationResult_hi_225, maskDestinationResult_lo_225};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_1 = {maskDestinationResult_hi_249, maskDestinationResult_lo_249, maskDestinationResult_hi_241, maskDestinationResult_lo_241};
  wire [15:0]   maskDestinationResult_hi_hi_hi_1 = {maskDestinationResult_hi_hi_hi_hi_1, maskDestinationResult_hi_hi_hi_lo_1};
  wire [31:0]   maskDestinationResult_hi_hi_1 = {maskDestinationResult_hi_hi_hi_1, maskDestinationResult_hi_hi_lo_1};
  wire [63:0]   maskDestinationResult_hi_257 = {maskDestinationResult_hi_hi_1, maskDestinationResult_hi_lo_1};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_2 = {maskDestinationResult_hi_10, maskDestinationResult_lo_10, maskDestinationResult_hi_2, maskDestinationResult_lo_2};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_2 = {maskDestinationResult_hi_26, maskDestinationResult_lo_26, maskDestinationResult_hi_18, maskDestinationResult_lo_18};
  wire [15:0]   maskDestinationResult_lo_lo_lo_2 = {maskDestinationResult_lo_lo_lo_hi_2, maskDestinationResult_lo_lo_lo_lo_2};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_2 = {maskDestinationResult_hi_42, maskDestinationResult_lo_42, maskDestinationResult_hi_34, maskDestinationResult_lo_34};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_2 = {maskDestinationResult_hi_58, maskDestinationResult_lo_58, maskDestinationResult_hi_50, maskDestinationResult_lo_50};
  wire [15:0]   maskDestinationResult_lo_lo_hi_2 = {maskDestinationResult_lo_lo_hi_hi_2, maskDestinationResult_lo_lo_hi_lo_2};
  wire [31:0]   maskDestinationResult_lo_lo_2 = {maskDestinationResult_lo_lo_hi_2, maskDestinationResult_lo_lo_lo_2};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_2 = {maskDestinationResult_hi_74, maskDestinationResult_lo_74, maskDestinationResult_hi_66, maskDestinationResult_lo_66};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_2 = {maskDestinationResult_hi_90, maskDestinationResult_lo_90, maskDestinationResult_hi_82, maskDestinationResult_lo_82};
  wire [15:0]   maskDestinationResult_lo_hi_lo_2 = {maskDestinationResult_lo_hi_lo_hi_2, maskDestinationResult_lo_hi_lo_lo_2};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_2 = {maskDestinationResult_hi_106, maskDestinationResult_lo_106, maskDestinationResult_hi_98, maskDestinationResult_lo_98};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_2 = {maskDestinationResult_hi_122, maskDestinationResult_lo_122, maskDestinationResult_hi_114, maskDestinationResult_lo_114};
  wire [15:0]   maskDestinationResult_lo_hi_hi_2 = {maskDestinationResult_lo_hi_hi_hi_2, maskDestinationResult_lo_hi_hi_lo_2};
  wire [31:0]   maskDestinationResult_lo_hi_2 = {maskDestinationResult_lo_hi_hi_2, maskDestinationResult_lo_hi_lo_2};
  wire [63:0]   maskDestinationResult_lo_258 = {maskDestinationResult_lo_hi_2, maskDestinationResult_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_2 = {maskDestinationResult_hi_138, maskDestinationResult_lo_138, maskDestinationResult_hi_130, maskDestinationResult_lo_130};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_2 = {maskDestinationResult_hi_154, maskDestinationResult_lo_154, maskDestinationResult_hi_146, maskDestinationResult_lo_146};
  wire [15:0]   maskDestinationResult_hi_lo_lo_2 = {maskDestinationResult_hi_lo_lo_hi_2, maskDestinationResult_hi_lo_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_2 = {maskDestinationResult_hi_170, maskDestinationResult_lo_170, maskDestinationResult_hi_162, maskDestinationResult_lo_162};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_2 = {maskDestinationResult_hi_186, maskDestinationResult_lo_186, maskDestinationResult_hi_178, maskDestinationResult_lo_178};
  wire [15:0]   maskDestinationResult_hi_lo_hi_2 = {maskDestinationResult_hi_lo_hi_hi_2, maskDestinationResult_hi_lo_hi_lo_2};
  wire [31:0]   maskDestinationResult_hi_lo_2 = {maskDestinationResult_hi_lo_hi_2, maskDestinationResult_hi_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_2 = {maskDestinationResult_hi_202, maskDestinationResult_lo_202, maskDestinationResult_hi_194, maskDestinationResult_lo_194};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_2 = {maskDestinationResult_hi_218, maskDestinationResult_lo_218, maskDestinationResult_hi_210, maskDestinationResult_lo_210};
  wire [15:0]   maskDestinationResult_hi_hi_lo_2 = {maskDestinationResult_hi_hi_lo_hi_2, maskDestinationResult_hi_hi_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_2 = {maskDestinationResult_hi_234, maskDestinationResult_lo_234, maskDestinationResult_hi_226, maskDestinationResult_lo_226};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_2 = {maskDestinationResult_hi_250, maskDestinationResult_lo_250, maskDestinationResult_hi_242, maskDestinationResult_lo_242};
  wire [15:0]   maskDestinationResult_hi_hi_hi_2 = {maskDestinationResult_hi_hi_hi_hi_2, maskDestinationResult_hi_hi_hi_lo_2};
  wire [31:0]   maskDestinationResult_hi_hi_2 = {maskDestinationResult_hi_hi_hi_2, maskDestinationResult_hi_hi_lo_2};
  wire [63:0]   maskDestinationResult_hi_258 = {maskDestinationResult_hi_hi_2, maskDestinationResult_hi_lo_2};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_3 = {maskDestinationResult_hi_11, maskDestinationResult_lo_11, maskDestinationResult_hi_3, maskDestinationResult_lo_3};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_3 = {maskDestinationResult_hi_27, maskDestinationResult_lo_27, maskDestinationResult_hi_19, maskDestinationResult_lo_19};
  wire [15:0]   maskDestinationResult_lo_lo_lo_3 = {maskDestinationResult_lo_lo_lo_hi_3, maskDestinationResult_lo_lo_lo_lo_3};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_3 = {maskDestinationResult_hi_43, maskDestinationResult_lo_43, maskDestinationResult_hi_35, maskDestinationResult_lo_35};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_3 = {maskDestinationResult_hi_59, maskDestinationResult_lo_59, maskDestinationResult_hi_51, maskDestinationResult_lo_51};
  wire [15:0]   maskDestinationResult_lo_lo_hi_3 = {maskDestinationResult_lo_lo_hi_hi_3, maskDestinationResult_lo_lo_hi_lo_3};
  wire [31:0]   maskDestinationResult_lo_lo_3 = {maskDestinationResult_lo_lo_hi_3, maskDestinationResult_lo_lo_lo_3};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_3 = {maskDestinationResult_hi_75, maskDestinationResult_lo_75, maskDestinationResult_hi_67, maskDestinationResult_lo_67};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_3 = {maskDestinationResult_hi_91, maskDestinationResult_lo_91, maskDestinationResult_hi_83, maskDestinationResult_lo_83};
  wire [15:0]   maskDestinationResult_lo_hi_lo_3 = {maskDestinationResult_lo_hi_lo_hi_3, maskDestinationResult_lo_hi_lo_lo_3};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_3 = {maskDestinationResult_hi_107, maskDestinationResult_lo_107, maskDestinationResult_hi_99, maskDestinationResult_lo_99};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_3 = {maskDestinationResult_hi_123, maskDestinationResult_lo_123, maskDestinationResult_hi_115, maskDestinationResult_lo_115};
  wire [15:0]   maskDestinationResult_lo_hi_hi_3 = {maskDestinationResult_lo_hi_hi_hi_3, maskDestinationResult_lo_hi_hi_lo_3};
  wire [31:0]   maskDestinationResult_lo_hi_3 = {maskDestinationResult_lo_hi_hi_3, maskDestinationResult_lo_hi_lo_3};
  wire [63:0]   maskDestinationResult_lo_259 = {maskDestinationResult_lo_hi_3, maskDestinationResult_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_3 = {maskDestinationResult_hi_139, maskDestinationResult_lo_139, maskDestinationResult_hi_131, maskDestinationResult_lo_131};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_3 = {maskDestinationResult_hi_155, maskDestinationResult_lo_155, maskDestinationResult_hi_147, maskDestinationResult_lo_147};
  wire [15:0]   maskDestinationResult_hi_lo_lo_3 = {maskDestinationResult_hi_lo_lo_hi_3, maskDestinationResult_hi_lo_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_3 = {maskDestinationResult_hi_171, maskDestinationResult_lo_171, maskDestinationResult_hi_163, maskDestinationResult_lo_163};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_3 = {maskDestinationResult_hi_187, maskDestinationResult_lo_187, maskDestinationResult_hi_179, maskDestinationResult_lo_179};
  wire [15:0]   maskDestinationResult_hi_lo_hi_3 = {maskDestinationResult_hi_lo_hi_hi_3, maskDestinationResult_hi_lo_hi_lo_3};
  wire [31:0]   maskDestinationResult_hi_lo_3 = {maskDestinationResult_hi_lo_hi_3, maskDestinationResult_hi_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_3 = {maskDestinationResult_hi_203, maskDestinationResult_lo_203, maskDestinationResult_hi_195, maskDestinationResult_lo_195};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_3 = {maskDestinationResult_hi_219, maskDestinationResult_lo_219, maskDestinationResult_hi_211, maskDestinationResult_lo_211};
  wire [15:0]   maskDestinationResult_hi_hi_lo_3 = {maskDestinationResult_hi_hi_lo_hi_3, maskDestinationResult_hi_hi_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_3 = {maskDestinationResult_hi_235, maskDestinationResult_lo_235, maskDestinationResult_hi_227, maskDestinationResult_lo_227};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_3 = {maskDestinationResult_hi_251, maskDestinationResult_lo_251, maskDestinationResult_hi_243, maskDestinationResult_lo_243};
  wire [15:0]   maskDestinationResult_hi_hi_hi_3 = {maskDestinationResult_hi_hi_hi_hi_3, maskDestinationResult_hi_hi_hi_lo_3};
  wire [31:0]   maskDestinationResult_hi_hi_3 = {maskDestinationResult_hi_hi_hi_3, maskDestinationResult_hi_hi_lo_3};
  wire [63:0]   maskDestinationResult_hi_259 = {maskDestinationResult_hi_hi_3, maskDestinationResult_hi_lo_3};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_4 = {maskDestinationResult_hi_12, maskDestinationResult_lo_12, maskDestinationResult_hi_4, maskDestinationResult_lo_4};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_4 = {maskDestinationResult_hi_28, maskDestinationResult_lo_28, maskDestinationResult_hi_20, maskDestinationResult_lo_20};
  wire [15:0]   maskDestinationResult_lo_lo_lo_4 = {maskDestinationResult_lo_lo_lo_hi_4, maskDestinationResult_lo_lo_lo_lo_4};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_4 = {maskDestinationResult_hi_44, maskDestinationResult_lo_44, maskDestinationResult_hi_36, maskDestinationResult_lo_36};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_4 = {maskDestinationResult_hi_60, maskDestinationResult_lo_60, maskDestinationResult_hi_52, maskDestinationResult_lo_52};
  wire [15:0]   maskDestinationResult_lo_lo_hi_4 = {maskDestinationResult_lo_lo_hi_hi_4, maskDestinationResult_lo_lo_hi_lo_4};
  wire [31:0]   maskDestinationResult_lo_lo_4 = {maskDestinationResult_lo_lo_hi_4, maskDestinationResult_lo_lo_lo_4};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_4 = {maskDestinationResult_hi_76, maskDestinationResult_lo_76, maskDestinationResult_hi_68, maskDestinationResult_lo_68};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_4 = {maskDestinationResult_hi_92, maskDestinationResult_lo_92, maskDestinationResult_hi_84, maskDestinationResult_lo_84};
  wire [15:0]   maskDestinationResult_lo_hi_lo_4 = {maskDestinationResult_lo_hi_lo_hi_4, maskDestinationResult_lo_hi_lo_lo_4};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_4 = {maskDestinationResult_hi_108, maskDestinationResult_lo_108, maskDestinationResult_hi_100, maskDestinationResult_lo_100};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_4 = {maskDestinationResult_hi_124, maskDestinationResult_lo_124, maskDestinationResult_hi_116, maskDestinationResult_lo_116};
  wire [15:0]   maskDestinationResult_lo_hi_hi_4 = {maskDestinationResult_lo_hi_hi_hi_4, maskDestinationResult_lo_hi_hi_lo_4};
  wire [31:0]   maskDestinationResult_lo_hi_4 = {maskDestinationResult_lo_hi_hi_4, maskDestinationResult_lo_hi_lo_4};
  wire [63:0]   maskDestinationResult_lo_260 = {maskDestinationResult_lo_hi_4, maskDestinationResult_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_4 = {maskDestinationResult_hi_140, maskDestinationResult_lo_140, maskDestinationResult_hi_132, maskDestinationResult_lo_132};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_4 = {maskDestinationResult_hi_156, maskDestinationResult_lo_156, maskDestinationResult_hi_148, maskDestinationResult_lo_148};
  wire [15:0]   maskDestinationResult_hi_lo_lo_4 = {maskDestinationResult_hi_lo_lo_hi_4, maskDestinationResult_hi_lo_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_4 = {maskDestinationResult_hi_172, maskDestinationResult_lo_172, maskDestinationResult_hi_164, maskDestinationResult_lo_164};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_4 = {maskDestinationResult_hi_188, maskDestinationResult_lo_188, maskDestinationResult_hi_180, maskDestinationResult_lo_180};
  wire [15:0]   maskDestinationResult_hi_lo_hi_4 = {maskDestinationResult_hi_lo_hi_hi_4, maskDestinationResult_hi_lo_hi_lo_4};
  wire [31:0]   maskDestinationResult_hi_lo_4 = {maskDestinationResult_hi_lo_hi_4, maskDestinationResult_hi_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_4 = {maskDestinationResult_hi_204, maskDestinationResult_lo_204, maskDestinationResult_hi_196, maskDestinationResult_lo_196};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_4 = {maskDestinationResult_hi_220, maskDestinationResult_lo_220, maskDestinationResult_hi_212, maskDestinationResult_lo_212};
  wire [15:0]   maskDestinationResult_hi_hi_lo_4 = {maskDestinationResult_hi_hi_lo_hi_4, maskDestinationResult_hi_hi_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_4 = {maskDestinationResult_hi_236, maskDestinationResult_lo_236, maskDestinationResult_hi_228, maskDestinationResult_lo_228};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_4 = {maskDestinationResult_hi_252, maskDestinationResult_lo_252, maskDestinationResult_hi_244, maskDestinationResult_lo_244};
  wire [15:0]   maskDestinationResult_hi_hi_hi_4 = {maskDestinationResult_hi_hi_hi_hi_4, maskDestinationResult_hi_hi_hi_lo_4};
  wire [31:0]   maskDestinationResult_hi_hi_4 = {maskDestinationResult_hi_hi_hi_4, maskDestinationResult_hi_hi_lo_4};
  wire [63:0]   maskDestinationResult_hi_260 = {maskDestinationResult_hi_hi_4, maskDestinationResult_hi_lo_4};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_5 = {maskDestinationResult_hi_13, maskDestinationResult_lo_13, maskDestinationResult_hi_5, maskDestinationResult_lo_5};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_5 = {maskDestinationResult_hi_29, maskDestinationResult_lo_29, maskDestinationResult_hi_21, maskDestinationResult_lo_21};
  wire [15:0]   maskDestinationResult_lo_lo_lo_5 = {maskDestinationResult_lo_lo_lo_hi_5, maskDestinationResult_lo_lo_lo_lo_5};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_5 = {maskDestinationResult_hi_45, maskDestinationResult_lo_45, maskDestinationResult_hi_37, maskDestinationResult_lo_37};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_5 = {maskDestinationResult_hi_61, maskDestinationResult_lo_61, maskDestinationResult_hi_53, maskDestinationResult_lo_53};
  wire [15:0]   maskDestinationResult_lo_lo_hi_5 = {maskDestinationResult_lo_lo_hi_hi_5, maskDestinationResult_lo_lo_hi_lo_5};
  wire [31:0]   maskDestinationResult_lo_lo_5 = {maskDestinationResult_lo_lo_hi_5, maskDestinationResult_lo_lo_lo_5};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_5 = {maskDestinationResult_hi_77, maskDestinationResult_lo_77, maskDestinationResult_hi_69, maskDestinationResult_lo_69};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_5 = {maskDestinationResult_hi_93, maskDestinationResult_lo_93, maskDestinationResult_hi_85, maskDestinationResult_lo_85};
  wire [15:0]   maskDestinationResult_lo_hi_lo_5 = {maskDestinationResult_lo_hi_lo_hi_5, maskDestinationResult_lo_hi_lo_lo_5};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_5 = {maskDestinationResult_hi_109, maskDestinationResult_lo_109, maskDestinationResult_hi_101, maskDestinationResult_lo_101};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_5 = {maskDestinationResult_hi_125, maskDestinationResult_lo_125, maskDestinationResult_hi_117, maskDestinationResult_lo_117};
  wire [15:0]   maskDestinationResult_lo_hi_hi_5 = {maskDestinationResult_lo_hi_hi_hi_5, maskDestinationResult_lo_hi_hi_lo_5};
  wire [31:0]   maskDestinationResult_lo_hi_5 = {maskDestinationResult_lo_hi_hi_5, maskDestinationResult_lo_hi_lo_5};
  wire [63:0]   maskDestinationResult_lo_261 = {maskDestinationResult_lo_hi_5, maskDestinationResult_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_5 = {maskDestinationResult_hi_141, maskDestinationResult_lo_141, maskDestinationResult_hi_133, maskDestinationResult_lo_133};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_5 = {maskDestinationResult_hi_157, maskDestinationResult_lo_157, maskDestinationResult_hi_149, maskDestinationResult_lo_149};
  wire [15:0]   maskDestinationResult_hi_lo_lo_5 = {maskDestinationResult_hi_lo_lo_hi_5, maskDestinationResult_hi_lo_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_5 = {maskDestinationResult_hi_173, maskDestinationResult_lo_173, maskDestinationResult_hi_165, maskDestinationResult_lo_165};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_5 = {maskDestinationResult_hi_189, maskDestinationResult_lo_189, maskDestinationResult_hi_181, maskDestinationResult_lo_181};
  wire [15:0]   maskDestinationResult_hi_lo_hi_5 = {maskDestinationResult_hi_lo_hi_hi_5, maskDestinationResult_hi_lo_hi_lo_5};
  wire [31:0]   maskDestinationResult_hi_lo_5 = {maskDestinationResult_hi_lo_hi_5, maskDestinationResult_hi_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_5 = {maskDestinationResult_hi_205, maskDestinationResult_lo_205, maskDestinationResult_hi_197, maskDestinationResult_lo_197};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_5 = {maskDestinationResult_hi_221, maskDestinationResult_lo_221, maskDestinationResult_hi_213, maskDestinationResult_lo_213};
  wire [15:0]   maskDestinationResult_hi_hi_lo_5 = {maskDestinationResult_hi_hi_lo_hi_5, maskDestinationResult_hi_hi_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_5 = {maskDestinationResult_hi_237, maskDestinationResult_lo_237, maskDestinationResult_hi_229, maskDestinationResult_lo_229};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_5 = {maskDestinationResult_hi_253, maskDestinationResult_lo_253, maskDestinationResult_hi_245, maskDestinationResult_lo_245};
  wire [15:0]   maskDestinationResult_hi_hi_hi_5 = {maskDestinationResult_hi_hi_hi_hi_5, maskDestinationResult_hi_hi_hi_lo_5};
  wire [31:0]   maskDestinationResult_hi_hi_5 = {maskDestinationResult_hi_hi_hi_5, maskDestinationResult_hi_hi_lo_5};
  wire [63:0]   maskDestinationResult_hi_261 = {maskDestinationResult_hi_hi_5, maskDestinationResult_hi_lo_5};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_6 = {maskDestinationResult_hi_14, maskDestinationResult_lo_14, maskDestinationResult_hi_6, maskDestinationResult_lo_6};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_6 = {maskDestinationResult_hi_30, maskDestinationResult_lo_30, maskDestinationResult_hi_22, maskDestinationResult_lo_22};
  wire [15:0]   maskDestinationResult_lo_lo_lo_6 = {maskDestinationResult_lo_lo_lo_hi_6, maskDestinationResult_lo_lo_lo_lo_6};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_6 = {maskDestinationResult_hi_46, maskDestinationResult_lo_46, maskDestinationResult_hi_38, maskDestinationResult_lo_38};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_6 = {maskDestinationResult_hi_62, maskDestinationResult_lo_62, maskDestinationResult_hi_54, maskDestinationResult_lo_54};
  wire [15:0]   maskDestinationResult_lo_lo_hi_6 = {maskDestinationResult_lo_lo_hi_hi_6, maskDestinationResult_lo_lo_hi_lo_6};
  wire [31:0]   maskDestinationResult_lo_lo_6 = {maskDestinationResult_lo_lo_hi_6, maskDestinationResult_lo_lo_lo_6};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_6 = {maskDestinationResult_hi_78, maskDestinationResult_lo_78, maskDestinationResult_hi_70, maskDestinationResult_lo_70};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_6 = {maskDestinationResult_hi_94, maskDestinationResult_lo_94, maskDestinationResult_hi_86, maskDestinationResult_lo_86};
  wire [15:0]   maskDestinationResult_lo_hi_lo_6 = {maskDestinationResult_lo_hi_lo_hi_6, maskDestinationResult_lo_hi_lo_lo_6};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_6 = {maskDestinationResult_hi_110, maskDestinationResult_lo_110, maskDestinationResult_hi_102, maskDestinationResult_lo_102};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_6 = {maskDestinationResult_hi_126, maskDestinationResult_lo_126, maskDestinationResult_hi_118, maskDestinationResult_lo_118};
  wire [15:0]   maskDestinationResult_lo_hi_hi_6 = {maskDestinationResult_lo_hi_hi_hi_6, maskDestinationResult_lo_hi_hi_lo_6};
  wire [31:0]   maskDestinationResult_lo_hi_6 = {maskDestinationResult_lo_hi_hi_6, maskDestinationResult_lo_hi_lo_6};
  wire [63:0]   maskDestinationResult_lo_262 = {maskDestinationResult_lo_hi_6, maskDestinationResult_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_6 = {maskDestinationResult_hi_142, maskDestinationResult_lo_142, maskDestinationResult_hi_134, maskDestinationResult_lo_134};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_6 = {maskDestinationResult_hi_158, maskDestinationResult_lo_158, maskDestinationResult_hi_150, maskDestinationResult_lo_150};
  wire [15:0]   maskDestinationResult_hi_lo_lo_6 = {maskDestinationResult_hi_lo_lo_hi_6, maskDestinationResult_hi_lo_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_6 = {maskDestinationResult_hi_174, maskDestinationResult_lo_174, maskDestinationResult_hi_166, maskDestinationResult_lo_166};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_6 = {maskDestinationResult_hi_190, maskDestinationResult_lo_190, maskDestinationResult_hi_182, maskDestinationResult_lo_182};
  wire [15:0]   maskDestinationResult_hi_lo_hi_6 = {maskDestinationResult_hi_lo_hi_hi_6, maskDestinationResult_hi_lo_hi_lo_6};
  wire [31:0]   maskDestinationResult_hi_lo_6 = {maskDestinationResult_hi_lo_hi_6, maskDestinationResult_hi_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_6 = {maskDestinationResult_hi_206, maskDestinationResult_lo_206, maskDestinationResult_hi_198, maskDestinationResult_lo_198};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_6 = {maskDestinationResult_hi_222, maskDestinationResult_lo_222, maskDestinationResult_hi_214, maskDestinationResult_lo_214};
  wire [15:0]   maskDestinationResult_hi_hi_lo_6 = {maskDestinationResult_hi_hi_lo_hi_6, maskDestinationResult_hi_hi_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_6 = {maskDestinationResult_hi_238, maskDestinationResult_lo_238, maskDestinationResult_hi_230, maskDestinationResult_lo_230};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_6 = {maskDestinationResult_hi_254, maskDestinationResult_lo_254, maskDestinationResult_hi_246, maskDestinationResult_lo_246};
  wire [15:0]   maskDestinationResult_hi_hi_hi_6 = {maskDestinationResult_hi_hi_hi_hi_6, maskDestinationResult_hi_hi_hi_lo_6};
  wire [31:0]   maskDestinationResult_hi_hi_6 = {maskDestinationResult_hi_hi_hi_6, maskDestinationResult_hi_hi_lo_6};
  wire [63:0]   maskDestinationResult_hi_262 = {maskDestinationResult_hi_hi_6, maskDestinationResult_hi_lo_6};
  wire [7:0]    maskDestinationResult_lo_lo_lo_lo_7 = {maskDestinationResult_hi_15, maskDestinationResult_lo_15, maskDestinationResult_hi_7, maskDestinationResult_lo_7};
  wire [7:0]    maskDestinationResult_lo_lo_lo_hi_7 = {maskDestinationResult_hi_31, maskDestinationResult_lo_31, maskDestinationResult_hi_23, maskDestinationResult_lo_23};
  wire [15:0]   maskDestinationResult_lo_lo_lo_7 = {maskDestinationResult_lo_lo_lo_hi_7, maskDestinationResult_lo_lo_lo_lo_7};
  wire [7:0]    maskDestinationResult_lo_lo_hi_lo_7 = {maskDestinationResult_hi_47, maskDestinationResult_lo_47, maskDestinationResult_hi_39, maskDestinationResult_lo_39};
  wire [7:0]    maskDestinationResult_lo_lo_hi_hi_7 = {maskDestinationResult_hi_63, maskDestinationResult_lo_63, maskDestinationResult_hi_55, maskDestinationResult_lo_55};
  wire [15:0]   maskDestinationResult_lo_lo_hi_7 = {maskDestinationResult_lo_lo_hi_hi_7, maskDestinationResult_lo_lo_hi_lo_7};
  wire [31:0]   maskDestinationResult_lo_lo_7 = {maskDestinationResult_lo_lo_hi_7, maskDestinationResult_lo_lo_lo_7};
  wire [7:0]    maskDestinationResult_lo_hi_lo_lo_7 = {maskDestinationResult_hi_79, maskDestinationResult_lo_79, maskDestinationResult_hi_71, maskDestinationResult_lo_71};
  wire [7:0]    maskDestinationResult_lo_hi_lo_hi_7 = {maskDestinationResult_hi_95, maskDestinationResult_lo_95, maskDestinationResult_hi_87, maskDestinationResult_lo_87};
  wire [15:0]   maskDestinationResult_lo_hi_lo_7 = {maskDestinationResult_lo_hi_lo_hi_7, maskDestinationResult_lo_hi_lo_lo_7};
  wire [7:0]    maskDestinationResult_lo_hi_hi_lo_7 = {maskDestinationResult_hi_111, maskDestinationResult_lo_111, maskDestinationResult_hi_103, maskDestinationResult_lo_103};
  wire [7:0]    maskDestinationResult_lo_hi_hi_hi_7 = {maskDestinationResult_hi_127, maskDestinationResult_lo_127, maskDestinationResult_hi_119, maskDestinationResult_lo_119};
  wire [15:0]   maskDestinationResult_lo_hi_hi_7 = {maskDestinationResult_lo_hi_hi_hi_7, maskDestinationResult_lo_hi_hi_lo_7};
  wire [31:0]   maskDestinationResult_lo_hi_7 = {maskDestinationResult_lo_hi_hi_7, maskDestinationResult_lo_hi_lo_7};
  wire [63:0]   maskDestinationResult_lo_263 = {maskDestinationResult_lo_hi_7, maskDestinationResult_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_lo_lo_lo_7 = {maskDestinationResult_hi_143, maskDestinationResult_lo_143, maskDestinationResult_hi_135, maskDestinationResult_lo_135};
  wire [7:0]    maskDestinationResult_hi_lo_lo_hi_7 = {maskDestinationResult_hi_159, maskDestinationResult_lo_159, maskDestinationResult_hi_151, maskDestinationResult_lo_151};
  wire [15:0]   maskDestinationResult_hi_lo_lo_7 = {maskDestinationResult_hi_lo_lo_hi_7, maskDestinationResult_hi_lo_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_lo_hi_lo_7 = {maskDestinationResult_hi_175, maskDestinationResult_lo_175, maskDestinationResult_hi_167, maskDestinationResult_lo_167};
  wire [7:0]    maskDestinationResult_hi_lo_hi_hi_7 = {maskDestinationResult_hi_191, maskDestinationResult_lo_191, maskDestinationResult_hi_183, maskDestinationResult_lo_183};
  wire [15:0]   maskDestinationResult_hi_lo_hi_7 = {maskDestinationResult_hi_lo_hi_hi_7, maskDestinationResult_hi_lo_hi_lo_7};
  wire [31:0]   maskDestinationResult_hi_lo_7 = {maskDestinationResult_hi_lo_hi_7, maskDestinationResult_hi_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_hi_lo_lo_7 = {maskDestinationResult_hi_207, maskDestinationResult_lo_207, maskDestinationResult_hi_199, maskDestinationResult_lo_199};
  wire [7:0]    maskDestinationResult_hi_hi_lo_hi_7 = {maskDestinationResult_hi_223, maskDestinationResult_lo_223, maskDestinationResult_hi_215, maskDestinationResult_lo_215};
  wire [15:0]   maskDestinationResult_hi_hi_lo_7 = {maskDestinationResult_hi_hi_lo_hi_7, maskDestinationResult_hi_hi_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_hi_hi_lo_7 = {maskDestinationResult_hi_239, maskDestinationResult_lo_239, maskDestinationResult_hi_231, maskDestinationResult_lo_231};
  wire [7:0]    maskDestinationResult_hi_hi_hi_hi_7 = {maskDestinationResult_hi_255, maskDestinationResult_lo_255, maskDestinationResult_hi_247, maskDestinationResult_lo_247};
  wire [15:0]   maskDestinationResult_hi_hi_hi_7 = {maskDestinationResult_hi_hi_hi_hi_7, maskDestinationResult_hi_hi_hi_lo_7};
  wire [31:0]   maskDestinationResult_hi_hi_7 = {maskDestinationResult_hi_hi_hi_7, maskDestinationResult_hi_hi_lo_7};
  wire [63:0]   maskDestinationResult_hi_263 = {maskDestinationResult_hi_hi_7, maskDestinationResult_hi_lo_7};
  wire [255:0]  maskDestinationResult_lo_lo_8 = {maskDestinationResult_hi_257, maskDestinationResult_lo_257, maskDestinationResult_hi_256, maskDestinationResult_lo_256};
  wire [255:0]  maskDestinationResult_lo_hi_8 = {maskDestinationResult_hi_259, maskDestinationResult_lo_259, maskDestinationResult_hi_258, maskDestinationResult_lo_258};
  wire [511:0]  maskDestinationResult_lo_264 = {maskDestinationResult_lo_hi_8, maskDestinationResult_lo_lo_8};
  wire [255:0]  maskDestinationResult_hi_lo_8 = {maskDestinationResult_hi_261, maskDestinationResult_lo_261, maskDestinationResult_hi_260, maskDestinationResult_lo_260};
  wire [255:0]  maskDestinationResult_hi_hi_8 = {maskDestinationResult_hi_263, maskDestinationResult_lo_263, maskDestinationResult_hi_262, maskDestinationResult_lo_262};
  wire [511:0]  maskDestinationResult_hi_264 = {maskDestinationResult_hi_hi_8, maskDestinationResult_hi_lo_8};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_8 = {sourceDataVec_1[1:0], sourceDataVec_0[1:0]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_8 = {sourceDataVec_3[1:0], sourceDataVec_2[1:0]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_8 = {maskDestinationResult_lo_lo_lo_hi_8, maskDestinationResult_lo_lo_lo_lo_8};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_8 = {sourceDataVec_5[1:0], sourceDataVec_4[1:0]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_8 = {sourceDataVec_7[1:0], sourceDataVec_6[1:0]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_8 = {maskDestinationResult_lo_lo_hi_hi_8, maskDestinationResult_lo_lo_hi_lo_8};
  wire [15:0]   maskDestinationResult_lo_lo_9 = {maskDestinationResult_lo_lo_hi_8, maskDestinationResult_lo_lo_lo_8};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_8 = {sourceDataVec_9[1:0], sourceDataVec_8[1:0]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_8 = {sourceDataVec_11[1:0], sourceDataVec_10[1:0]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_8 = {maskDestinationResult_lo_hi_lo_hi_8, maskDestinationResult_lo_hi_lo_lo_8};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_8 = {sourceDataVec_13[1:0], sourceDataVec_12[1:0]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_8 = {sourceDataVec_15[1:0], sourceDataVec_14[1:0]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_8 = {maskDestinationResult_lo_hi_hi_hi_8, maskDestinationResult_lo_hi_hi_lo_8};
  wire [15:0]   maskDestinationResult_lo_hi_9 = {maskDestinationResult_lo_hi_hi_8, maskDestinationResult_lo_hi_lo_8};
  wire [31:0]   maskDestinationResult_lo_265 = {maskDestinationResult_lo_hi_9, maskDestinationResult_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_8 = {sourceDataVec_17[1:0], sourceDataVec_16[1:0]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_8 = {sourceDataVec_19[1:0], sourceDataVec_18[1:0]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_8 = {maskDestinationResult_hi_lo_lo_hi_8, maskDestinationResult_hi_lo_lo_lo_8};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_8 = {sourceDataVec_21[1:0], sourceDataVec_20[1:0]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_8 = {sourceDataVec_23[1:0], sourceDataVec_22[1:0]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_8 = {maskDestinationResult_hi_lo_hi_hi_8, maskDestinationResult_hi_lo_hi_lo_8};
  wire [15:0]   maskDestinationResult_hi_lo_9 = {maskDestinationResult_hi_lo_hi_8, maskDestinationResult_hi_lo_lo_8};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_8 = {sourceDataVec_25[1:0], sourceDataVec_24[1:0]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_8 = {sourceDataVec_27[1:0], sourceDataVec_26[1:0]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_8 = {maskDestinationResult_hi_hi_lo_hi_8, maskDestinationResult_hi_hi_lo_lo_8};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_8 = {sourceDataVec_29[1:0], sourceDataVec_28[1:0]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_8 = {sourceDataVec_31[1:0], sourceDataVec_30[1:0]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_8 = {maskDestinationResult_hi_hi_hi_hi_8, maskDestinationResult_hi_hi_hi_lo_8};
  wire [15:0]   maskDestinationResult_hi_hi_9 = {maskDestinationResult_hi_hi_hi_8, maskDestinationResult_hi_hi_lo_8};
  wire [31:0]   maskDestinationResult_hi_265 = {maskDestinationResult_hi_hi_9, maskDestinationResult_hi_lo_9};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_9 = {sourceDataVec_1[3:2], sourceDataVec_0[3:2]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_9 = {sourceDataVec_3[3:2], sourceDataVec_2[3:2]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_9 = {maskDestinationResult_lo_lo_lo_hi_9, maskDestinationResult_lo_lo_lo_lo_9};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_9 = {sourceDataVec_5[3:2], sourceDataVec_4[3:2]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_9 = {sourceDataVec_7[3:2], sourceDataVec_6[3:2]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_9 = {maskDestinationResult_lo_lo_hi_hi_9, maskDestinationResult_lo_lo_hi_lo_9};
  wire [15:0]   maskDestinationResult_lo_lo_10 = {maskDestinationResult_lo_lo_hi_9, maskDestinationResult_lo_lo_lo_9};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_9 = {sourceDataVec_9[3:2], sourceDataVec_8[3:2]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_9 = {sourceDataVec_11[3:2], sourceDataVec_10[3:2]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_9 = {maskDestinationResult_lo_hi_lo_hi_9, maskDestinationResult_lo_hi_lo_lo_9};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_9 = {sourceDataVec_13[3:2], sourceDataVec_12[3:2]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_9 = {sourceDataVec_15[3:2], sourceDataVec_14[3:2]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_9 = {maskDestinationResult_lo_hi_hi_hi_9, maskDestinationResult_lo_hi_hi_lo_9};
  wire [15:0]   maskDestinationResult_lo_hi_10 = {maskDestinationResult_lo_hi_hi_9, maskDestinationResult_lo_hi_lo_9};
  wire [31:0]   maskDestinationResult_lo_266 = {maskDestinationResult_lo_hi_10, maskDestinationResult_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_9 = {sourceDataVec_17[3:2], sourceDataVec_16[3:2]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_9 = {sourceDataVec_19[3:2], sourceDataVec_18[3:2]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_9 = {maskDestinationResult_hi_lo_lo_hi_9, maskDestinationResult_hi_lo_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_9 = {sourceDataVec_21[3:2], sourceDataVec_20[3:2]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_9 = {sourceDataVec_23[3:2], sourceDataVec_22[3:2]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_9 = {maskDestinationResult_hi_lo_hi_hi_9, maskDestinationResult_hi_lo_hi_lo_9};
  wire [15:0]   maskDestinationResult_hi_lo_10 = {maskDestinationResult_hi_lo_hi_9, maskDestinationResult_hi_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_9 = {sourceDataVec_25[3:2], sourceDataVec_24[3:2]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_9 = {sourceDataVec_27[3:2], sourceDataVec_26[3:2]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_9 = {maskDestinationResult_hi_hi_lo_hi_9, maskDestinationResult_hi_hi_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_9 = {sourceDataVec_29[3:2], sourceDataVec_28[3:2]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_9 = {sourceDataVec_31[3:2], sourceDataVec_30[3:2]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_9 = {maskDestinationResult_hi_hi_hi_hi_9, maskDestinationResult_hi_hi_hi_lo_9};
  wire [15:0]   maskDestinationResult_hi_hi_10 = {maskDestinationResult_hi_hi_hi_9, maskDestinationResult_hi_hi_lo_9};
  wire [31:0]   maskDestinationResult_hi_266 = {maskDestinationResult_hi_hi_10, maskDestinationResult_hi_lo_10};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_10 = {sourceDataVec_1[5:4], sourceDataVec_0[5:4]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_10 = {sourceDataVec_3[5:4], sourceDataVec_2[5:4]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_10 = {maskDestinationResult_lo_lo_lo_hi_10, maskDestinationResult_lo_lo_lo_lo_10};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_10 = {sourceDataVec_5[5:4], sourceDataVec_4[5:4]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_10 = {sourceDataVec_7[5:4], sourceDataVec_6[5:4]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_10 = {maskDestinationResult_lo_lo_hi_hi_10, maskDestinationResult_lo_lo_hi_lo_10};
  wire [15:0]   maskDestinationResult_lo_lo_11 = {maskDestinationResult_lo_lo_hi_10, maskDestinationResult_lo_lo_lo_10};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_10 = {sourceDataVec_9[5:4], sourceDataVec_8[5:4]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_10 = {sourceDataVec_11[5:4], sourceDataVec_10[5:4]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_10 = {maskDestinationResult_lo_hi_lo_hi_10, maskDestinationResult_lo_hi_lo_lo_10};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_10 = {sourceDataVec_13[5:4], sourceDataVec_12[5:4]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_10 = {sourceDataVec_15[5:4], sourceDataVec_14[5:4]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_10 = {maskDestinationResult_lo_hi_hi_hi_10, maskDestinationResult_lo_hi_hi_lo_10};
  wire [15:0]   maskDestinationResult_lo_hi_11 = {maskDestinationResult_lo_hi_hi_10, maskDestinationResult_lo_hi_lo_10};
  wire [31:0]   maskDestinationResult_lo_267 = {maskDestinationResult_lo_hi_11, maskDestinationResult_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_10 = {sourceDataVec_17[5:4], sourceDataVec_16[5:4]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_10 = {sourceDataVec_19[5:4], sourceDataVec_18[5:4]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_10 = {maskDestinationResult_hi_lo_lo_hi_10, maskDestinationResult_hi_lo_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_10 = {sourceDataVec_21[5:4], sourceDataVec_20[5:4]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_10 = {sourceDataVec_23[5:4], sourceDataVec_22[5:4]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_10 = {maskDestinationResult_hi_lo_hi_hi_10, maskDestinationResult_hi_lo_hi_lo_10};
  wire [15:0]   maskDestinationResult_hi_lo_11 = {maskDestinationResult_hi_lo_hi_10, maskDestinationResult_hi_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_10 = {sourceDataVec_25[5:4], sourceDataVec_24[5:4]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_10 = {sourceDataVec_27[5:4], sourceDataVec_26[5:4]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_10 = {maskDestinationResult_hi_hi_lo_hi_10, maskDestinationResult_hi_hi_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_10 = {sourceDataVec_29[5:4], sourceDataVec_28[5:4]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_10 = {sourceDataVec_31[5:4], sourceDataVec_30[5:4]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_10 = {maskDestinationResult_hi_hi_hi_hi_10, maskDestinationResult_hi_hi_hi_lo_10};
  wire [15:0]   maskDestinationResult_hi_hi_11 = {maskDestinationResult_hi_hi_hi_10, maskDestinationResult_hi_hi_lo_10};
  wire [31:0]   maskDestinationResult_hi_267 = {maskDestinationResult_hi_hi_11, maskDestinationResult_hi_lo_11};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_11 = {sourceDataVec_1[7:6], sourceDataVec_0[7:6]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_11 = {sourceDataVec_3[7:6], sourceDataVec_2[7:6]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_11 = {maskDestinationResult_lo_lo_lo_hi_11, maskDestinationResult_lo_lo_lo_lo_11};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_11 = {sourceDataVec_5[7:6], sourceDataVec_4[7:6]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_11 = {sourceDataVec_7[7:6], sourceDataVec_6[7:6]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_11 = {maskDestinationResult_lo_lo_hi_hi_11, maskDestinationResult_lo_lo_hi_lo_11};
  wire [15:0]   maskDestinationResult_lo_lo_12 = {maskDestinationResult_lo_lo_hi_11, maskDestinationResult_lo_lo_lo_11};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_11 = {sourceDataVec_9[7:6], sourceDataVec_8[7:6]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_11 = {sourceDataVec_11[7:6], sourceDataVec_10[7:6]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_11 = {maskDestinationResult_lo_hi_lo_hi_11, maskDestinationResult_lo_hi_lo_lo_11};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_11 = {sourceDataVec_13[7:6], sourceDataVec_12[7:6]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_11 = {sourceDataVec_15[7:6], sourceDataVec_14[7:6]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_11 = {maskDestinationResult_lo_hi_hi_hi_11, maskDestinationResult_lo_hi_hi_lo_11};
  wire [15:0]   maskDestinationResult_lo_hi_12 = {maskDestinationResult_lo_hi_hi_11, maskDestinationResult_lo_hi_lo_11};
  wire [31:0]   maskDestinationResult_lo_268 = {maskDestinationResult_lo_hi_12, maskDestinationResult_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_11 = {sourceDataVec_17[7:6], sourceDataVec_16[7:6]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_11 = {sourceDataVec_19[7:6], sourceDataVec_18[7:6]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_11 = {maskDestinationResult_hi_lo_lo_hi_11, maskDestinationResult_hi_lo_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_11 = {sourceDataVec_21[7:6], sourceDataVec_20[7:6]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_11 = {sourceDataVec_23[7:6], sourceDataVec_22[7:6]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_11 = {maskDestinationResult_hi_lo_hi_hi_11, maskDestinationResult_hi_lo_hi_lo_11};
  wire [15:0]   maskDestinationResult_hi_lo_12 = {maskDestinationResult_hi_lo_hi_11, maskDestinationResult_hi_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_11 = {sourceDataVec_25[7:6], sourceDataVec_24[7:6]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_11 = {sourceDataVec_27[7:6], sourceDataVec_26[7:6]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_11 = {maskDestinationResult_hi_hi_lo_hi_11, maskDestinationResult_hi_hi_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_11 = {sourceDataVec_29[7:6], sourceDataVec_28[7:6]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_11 = {sourceDataVec_31[7:6], sourceDataVec_30[7:6]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_11 = {maskDestinationResult_hi_hi_hi_hi_11, maskDestinationResult_hi_hi_hi_lo_11};
  wire [15:0]   maskDestinationResult_hi_hi_12 = {maskDestinationResult_hi_hi_hi_11, maskDestinationResult_hi_hi_lo_11};
  wire [31:0]   maskDestinationResult_hi_268 = {maskDestinationResult_hi_hi_12, maskDestinationResult_hi_lo_12};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_12 = {sourceDataVec_1[9:8], sourceDataVec_0[9:8]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_12 = {sourceDataVec_3[9:8], sourceDataVec_2[9:8]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_12 = {maskDestinationResult_lo_lo_lo_hi_12, maskDestinationResult_lo_lo_lo_lo_12};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_12 = {sourceDataVec_5[9:8], sourceDataVec_4[9:8]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_12 = {sourceDataVec_7[9:8], sourceDataVec_6[9:8]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_12 = {maskDestinationResult_lo_lo_hi_hi_12, maskDestinationResult_lo_lo_hi_lo_12};
  wire [15:0]   maskDestinationResult_lo_lo_13 = {maskDestinationResult_lo_lo_hi_12, maskDestinationResult_lo_lo_lo_12};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_12 = {sourceDataVec_9[9:8], sourceDataVec_8[9:8]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_12 = {sourceDataVec_11[9:8], sourceDataVec_10[9:8]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_12 = {maskDestinationResult_lo_hi_lo_hi_12, maskDestinationResult_lo_hi_lo_lo_12};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_12 = {sourceDataVec_13[9:8], sourceDataVec_12[9:8]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_12 = {sourceDataVec_15[9:8], sourceDataVec_14[9:8]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_12 = {maskDestinationResult_lo_hi_hi_hi_12, maskDestinationResult_lo_hi_hi_lo_12};
  wire [15:0]   maskDestinationResult_lo_hi_13 = {maskDestinationResult_lo_hi_hi_12, maskDestinationResult_lo_hi_lo_12};
  wire [31:0]   maskDestinationResult_lo_269 = {maskDestinationResult_lo_hi_13, maskDestinationResult_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_12 = {sourceDataVec_17[9:8], sourceDataVec_16[9:8]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_12 = {sourceDataVec_19[9:8], sourceDataVec_18[9:8]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_12 = {maskDestinationResult_hi_lo_lo_hi_12, maskDestinationResult_hi_lo_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_12 = {sourceDataVec_21[9:8], sourceDataVec_20[9:8]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_12 = {sourceDataVec_23[9:8], sourceDataVec_22[9:8]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_12 = {maskDestinationResult_hi_lo_hi_hi_12, maskDestinationResult_hi_lo_hi_lo_12};
  wire [15:0]   maskDestinationResult_hi_lo_13 = {maskDestinationResult_hi_lo_hi_12, maskDestinationResult_hi_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_12 = {sourceDataVec_25[9:8], sourceDataVec_24[9:8]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_12 = {sourceDataVec_27[9:8], sourceDataVec_26[9:8]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_12 = {maskDestinationResult_hi_hi_lo_hi_12, maskDestinationResult_hi_hi_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_12 = {sourceDataVec_29[9:8], sourceDataVec_28[9:8]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_12 = {sourceDataVec_31[9:8], sourceDataVec_30[9:8]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_12 = {maskDestinationResult_hi_hi_hi_hi_12, maskDestinationResult_hi_hi_hi_lo_12};
  wire [15:0]   maskDestinationResult_hi_hi_13 = {maskDestinationResult_hi_hi_hi_12, maskDestinationResult_hi_hi_lo_12};
  wire [31:0]   maskDestinationResult_hi_269 = {maskDestinationResult_hi_hi_13, maskDestinationResult_hi_lo_13};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_13 = {sourceDataVec_1[11:10], sourceDataVec_0[11:10]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_13 = {sourceDataVec_3[11:10], sourceDataVec_2[11:10]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_13 = {maskDestinationResult_lo_lo_lo_hi_13, maskDestinationResult_lo_lo_lo_lo_13};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_13 = {sourceDataVec_5[11:10], sourceDataVec_4[11:10]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_13 = {sourceDataVec_7[11:10], sourceDataVec_6[11:10]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_13 = {maskDestinationResult_lo_lo_hi_hi_13, maskDestinationResult_lo_lo_hi_lo_13};
  wire [15:0]   maskDestinationResult_lo_lo_14 = {maskDestinationResult_lo_lo_hi_13, maskDestinationResult_lo_lo_lo_13};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_13 = {sourceDataVec_9[11:10], sourceDataVec_8[11:10]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_13 = {sourceDataVec_11[11:10], sourceDataVec_10[11:10]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_13 = {maskDestinationResult_lo_hi_lo_hi_13, maskDestinationResult_lo_hi_lo_lo_13};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_13 = {sourceDataVec_13[11:10], sourceDataVec_12[11:10]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_13 = {sourceDataVec_15[11:10], sourceDataVec_14[11:10]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_13 = {maskDestinationResult_lo_hi_hi_hi_13, maskDestinationResult_lo_hi_hi_lo_13};
  wire [15:0]   maskDestinationResult_lo_hi_14 = {maskDestinationResult_lo_hi_hi_13, maskDestinationResult_lo_hi_lo_13};
  wire [31:0]   maskDestinationResult_lo_270 = {maskDestinationResult_lo_hi_14, maskDestinationResult_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_13 = {sourceDataVec_17[11:10], sourceDataVec_16[11:10]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_13 = {sourceDataVec_19[11:10], sourceDataVec_18[11:10]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_13 = {maskDestinationResult_hi_lo_lo_hi_13, maskDestinationResult_hi_lo_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_13 = {sourceDataVec_21[11:10], sourceDataVec_20[11:10]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_13 = {sourceDataVec_23[11:10], sourceDataVec_22[11:10]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_13 = {maskDestinationResult_hi_lo_hi_hi_13, maskDestinationResult_hi_lo_hi_lo_13};
  wire [15:0]   maskDestinationResult_hi_lo_14 = {maskDestinationResult_hi_lo_hi_13, maskDestinationResult_hi_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_13 = {sourceDataVec_25[11:10], sourceDataVec_24[11:10]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_13 = {sourceDataVec_27[11:10], sourceDataVec_26[11:10]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_13 = {maskDestinationResult_hi_hi_lo_hi_13, maskDestinationResult_hi_hi_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_13 = {sourceDataVec_29[11:10], sourceDataVec_28[11:10]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_13 = {sourceDataVec_31[11:10], sourceDataVec_30[11:10]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_13 = {maskDestinationResult_hi_hi_hi_hi_13, maskDestinationResult_hi_hi_hi_lo_13};
  wire [15:0]   maskDestinationResult_hi_hi_14 = {maskDestinationResult_hi_hi_hi_13, maskDestinationResult_hi_hi_lo_13};
  wire [31:0]   maskDestinationResult_hi_270 = {maskDestinationResult_hi_hi_14, maskDestinationResult_hi_lo_14};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_14 = {sourceDataVec_1[13:12], sourceDataVec_0[13:12]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_14 = {sourceDataVec_3[13:12], sourceDataVec_2[13:12]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_14 = {maskDestinationResult_lo_lo_lo_hi_14, maskDestinationResult_lo_lo_lo_lo_14};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_14 = {sourceDataVec_5[13:12], sourceDataVec_4[13:12]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_14 = {sourceDataVec_7[13:12], sourceDataVec_6[13:12]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_14 = {maskDestinationResult_lo_lo_hi_hi_14, maskDestinationResult_lo_lo_hi_lo_14};
  wire [15:0]   maskDestinationResult_lo_lo_15 = {maskDestinationResult_lo_lo_hi_14, maskDestinationResult_lo_lo_lo_14};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_14 = {sourceDataVec_9[13:12], sourceDataVec_8[13:12]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_14 = {sourceDataVec_11[13:12], sourceDataVec_10[13:12]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_14 = {maskDestinationResult_lo_hi_lo_hi_14, maskDestinationResult_lo_hi_lo_lo_14};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_14 = {sourceDataVec_13[13:12], sourceDataVec_12[13:12]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_14 = {sourceDataVec_15[13:12], sourceDataVec_14[13:12]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_14 = {maskDestinationResult_lo_hi_hi_hi_14, maskDestinationResult_lo_hi_hi_lo_14};
  wire [15:0]   maskDestinationResult_lo_hi_15 = {maskDestinationResult_lo_hi_hi_14, maskDestinationResult_lo_hi_lo_14};
  wire [31:0]   maskDestinationResult_lo_271 = {maskDestinationResult_lo_hi_15, maskDestinationResult_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_14 = {sourceDataVec_17[13:12], sourceDataVec_16[13:12]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_14 = {sourceDataVec_19[13:12], sourceDataVec_18[13:12]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_14 = {maskDestinationResult_hi_lo_lo_hi_14, maskDestinationResult_hi_lo_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_14 = {sourceDataVec_21[13:12], sourceDataVec_20[13:12]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_14 = {sourceDataVec_23[13:12], sourceDataVec_22[13:12]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_14 = {maskDestinationResult_hi_lo_hi_hi_14, maskDestinationResult_hi_lo_hi_lo_14};
  wire [15:0]   maskDestinationResult_hi_lo_15 = {maskDestinationResult_hi_lo_hi_14, maskDestinationResult_hi_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_14 = {sourceDataVec_25[13:12], sourceDataVec_24[13:12]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_14 = {sourceDataVec_27[13:12], sourceDataVec_26[13:12]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_14 = {maskDestinationResult_hi_hi_lo_hi_14, maskDestinationResult_hi_hi_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_14 = {sourceDataVec_29[13:12], sourceDataVec_28[13:12]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_14 = {sourceDataVec_31[13:12], sourceDataVec_30[13:12]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_14 = {maskDestinationResult_hi_hi_hi_hi_14, maskDestinationResult_hi_hi_hi_lo_14};
  wire [15:0]   maskDestinationResult_hi_hi_15 = {maskDestinationResult_hi_hi_hi_14, maskDestinationResult_hi_hi_lo_14};
  wire [31:0]   maskDestinationResult_hi_271 = {maskDestinationResult_hi_hi_15, maskDestinationResult_hi_lo_15};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_15 = {sourceDataVec_1[15:14], sourceDataVec_0[15:14]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_15 = {sourceDataVec_3[15:14], sourceDataVec_2[15:14]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_15 = {maskDestinationResult_lo_lo_lo_hi_15, maskDestinationResult_lo_lo_lo_lo_15};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_15 = {sourceDataVec_5[15:14], sourceDataVec_4[15:14]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_15 = {sourceDataVec_7[15:14], sourceDataVec_6[15:14]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_15 = {maskDestinationResult_lo_lo_hi_hi_15, maskDestinationResult_lo_lo_hi_lo_15};
  wire [15:0]   maskDestinationResult_lo_lo_16 = {maskDestinationResult_lo_lo_hi_15, maskDestinationResult_lo_lo_lo_15};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_15 = {sourceDataVec_9[15:14], sourceDataVec_8[15:14]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_15 = {sourceDataVec_11[15:14], sourceDataVec_10[15:14]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_15 = {maskDestinationResult_lo_hi_lo_hi_15, maskDestinationResult_lo_hi_lo_lo_15};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_15 = {sourceDataVec_13[15:14], sourceDataVec_12[15:14]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_15 = {sourceDataVec_15[15:14], sourceDataVec_14[15:14]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_15 = {maskDestinationResult_lo_hi_hi_hi_15, maskDestinationResult_lo_hi_hi_lo_15};
  wire [15:0]   maskDestinationResult_lo_hi_16 = {maskDestinationResult_lo_hi_hi_15, maskDestinationResult_lo_hi_lo_15};
  wire [31:0]   maskDestinationResult_lo_272 = {maskDestinationResult_lo_hi_16, maskDestinationResult_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_15 = {sourceDataVec_17[15:14], sourceDataVec_16[15:14]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_15 = {sourceDataVec_19[15:14], sourceDataVec_18[15:14]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_15 = {maskDestinationResult_hi_lo_lo_hi_15, maskDestinationResult_hi_lo_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_15 = {sourceDataVec_21[15:14], sourceDataVec_20[15:14]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_15 = {sourceDataVec_23[15:14], sourceDataVec_22[15:14]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_15 = {maskDestinationResult_hi_lo_hi_hi_15, maskDestinationResult_hi_lo_hi_lo_15};
  wire [15:0]   maskDestinationResult_hi_lo_16 = {maskDestinationResult_hi_lo_hi_15, maskDestinationResult_hi_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_15 = {sourceDataVec_25[15:14], sourceDataVec_24[15:14]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_15 = {sourceDataVec_27[15:14], sourceDataVec_26[15:14]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_15 = {maskDestinationResult_hi_hi_lo_hi_15, maskDestinationResult_hi_hi_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_15 = {sourceDataVec_29[15:14], sourceDataVec_28[15:14]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_15 = {sourceDataVec_31[15:14], sourceDataVec_30[15:14]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_15 = {maskDestinationResult_hi_hi_hi_hi_15, maskDestinationResult_hi_hi_hi_lo_15};
  wire [15:0]   maskDestinationResult_hi_hi_16 = {maskDestinationResult_hi_hi_hi_15, maskDestinationResult_hi_hi_lo_15};
  wire [31:0]   maskDestinationResult_hi_272 = {maskDestinationResult_hi_hi_16, maskDestinationResult_hi_lo_16};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_16 = {sourceDataVec_1[17:16], sourceDataVec_0[17:16]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_16 = {sourceDataVec_3[17:16], sourceDataVec_2[17:16]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_16 = {maskDestinationResult_lo_lo_lo_hi_16, maskDestinationResult_lo_lo_lo_lo_16};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_16 = {sourceDataVec_5[17:16], sourceDataVec_4[17:16]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_16 = {sourceDataVec_7[17:16], sourceDataVec_6[17:16]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_16 = {maskDestinationResult_lo_lo_hi_hi_16, maskDestinationResult_lo_lo_hi_lo_16};
  wire [15:0]   maskDestinationResult_lo_lo_17 = {maskDestinationResult_lo_lo_hi_16, maskDestinationResult_lo_lo_lo_16};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_16 = {sourceDataVec_9[17:16], sourceDataVec_8[17:16]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_16 = {sourceDataVec_11[17:16], sourceDataVec_10[17:16]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_16 = {maskDestinationResult_lo_hi_lo_hi_16, maskDestinationResult_lo_hi_lo_lo_16};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_16 = {sourceDataVec_13[17:16], sourceDataVec_12[17:16]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_16 = {sourceDataVec_15[17:16], sourceDataVec_14[17:16]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_16 = {maskDestinationResult_lo_hi_hi_hi_16, maskDestinationResult_lo_hi_hi_lo_16};
  wire [15:0]   maskDestinationResult_lo_hi_17 = {maskDestinationResult_lo_hi_hi_16, maskDestinationResult_lo_hi_lo_16};
  wire [31:0]   maskDestinationResult_lo_273 = {maskDestinationResult_lo_hi_17, maskDestinationResult_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_16 = {sourceDataVec_17[17:16], sourceDataVec_16[17:16]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_16 = {sourceDataVec_19[17:16], sourceDataVec_18[17:16]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_16 = {maskDestinationResult_hi_lo_lo_hi_16, maskDestinationResult_hi_lo_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_16 = {sourceDataVec_21[17:16], sourceDataVec_20[17:16]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_16 = {sourceDataVec_23[17:16], sourceDataVec_22[17:16]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_16 = {maskDestinationResult_hi_lo_hi_hi_16, maskDestinationResult_hi_lo_hi_lo_16};
  wire [15:0]   maskDestinationResult_hi_lo_17 = {maskDestinationResult_hi_lo_hi_16, maskDestinationResult_hi_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_16 = {sourceDataVec_25[17:16], sourceDataVec_24[17:16]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_16 = {sourceDataVec_27[17:16], sourceDataVec_26[17:16]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_16 = {maskDestinationResult_hi_hi_lo_hi_16, maskDestinationResult_hi_hi_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_16 = {sourceDataVec_29[17:16], sourceDataVec_28[17:16]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_16 = {sourceDataVec_31[17:16], sourceDataVec_30[17:16]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_16 = {maskDestinationResult_hi_hi_hi_hi_16, maskDestinationResult_hi_hi_hi_lo_16};
  wire [15:0]   maskDestinationResult_hi_hi_17 = {maskDestinationResult_hi_hi_hi_16, maskDestinationResult_hi_hi_lo_16};
  wire [31:0]   maskDestinationResult_hi_273 = {maskDestinationResult_hi_hi_17, maskDestinationResult_hi_lo_17};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_17 = {sourceDataVec_1[19:18], sourceDataVec_0[19:18]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_17 = {sourceDataVec_3[19:18], sourceDataVec_2[19:18]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_17 = {maskDestinationResult_lo_lo_lo_hi_17, maskDestinationResult_lo_lo_lo_lo_17};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_17 = {sourceDataVec_5[19:18], sourceDataVec_4[19:18]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_17 = {sourceDataVec_7[19:18], sourceDataVec_6[19:18]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_17 = {maskDestinationResult_lo_lo_hi_hi_17, maskDestinationResult_lo_lo_hi_lo_17};
  wire [15:0]   maskDestinationResult_lo_lo_18 = {maskDestinationResult_lo_lo_hi_17, maskDestinationResult_lo_lo_lo_17};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_17 = {sourceDataVec_9[19:18], sourceDataVec_8[19:18]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_17 = {sourceDataVec_11[19:18], sourceDataVec_10[19:18]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_17 = {maskDestinationResult_lo_hi_lo_hi_17, maskDestinationResult_lo_hi_lo_lo_17};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_17 = {sourceDataVec_13[19:18], sourceDataVec_12[19:18]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_17 = {sourceDataVec_15[19:18], sourceDataVec_14[19:18]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_17 = {maskDestinationResult_lo_hi_hi_hi_17, maskDestinationResult_lo_hi_hi_lo_17};
  wire [15:0]   maskDestinationResult_lo_hi_18 = {maskDestinationResult_lo_hi_hi_17, maskDestinationResult_lo_hi_lo_17};
  wire [31:0]   maskDestinationResult_lo_274 = {maskDestinationResult_lo_hi_18, maskDestinationResult_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_17 = {sourceDataVec_17[19:18], sourceDataVec_16[19:18]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_17 = {sourceDataVec_19[19:18], sourceDataVec_18[19:18]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_17 = {maskDestinationResult_hi_lo_lo_hi_17, maskDestinationResult_hi_lo_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_17 = {sourceDataVec_21[19:18], sourceDataVec_20[19:18]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_17 = {sourceDataVec_23[19:18], sourceDataVec_22[19:18]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_17 = {maskDestinationResult_hi_lo_hi_hi_17, maskDestinationResult_hi_lo_hi_lo_17};
  wire [15:0]   maskDestinationResult_hi_lo_18 = {maskDestinationResult_hi_lo_hi_17, maskDestinationResult_hi_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_17 = {sourceDataVec_25[19:18], sourceDataVec_24[19:18]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_17 = {sourceDataVec_27[19:18], sourceDataVec_26[19:18]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_17 = {maskDestinationResult_hi_hi_lo_hi_17, maskDestinationResult_hi_hi_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_17 = {sourceDataVec_29[19:18], sourceDataVec_28[19:18]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_17 = {sourceDataVec_31[19:18], sourceDataVec_30[19:18]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_17 = {maskDestinationResult_hi_hi_hi_hi_17, maskDestinationResult_hi_hi_hi_lo_17};
  wire [15:0]   maskDestinationResult_hi_hi_18 = {maskDestinationResult_hi_hi_hi_17, maskDestinationResult_hi_hi_lo_17};
  wire [31:0]   maskDestinationResult_hi_274 = {maskDestinationResult_hi_hi_18, maskDestinationResult_hi_lo_18};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_18 = {sourceDataVec_1[21:20], sourceDataVec_0[21:20]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_18 = {sourceDataVec_3[21:20], sourceDataVec_2[21:20]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_18 = {maskDestinationResult_lo_lo_lo_hi_18, maskDestinationResult_lo_lo_lo_lo_18};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_18 = {sourceDataVec_5[21:20], sourceDataVec_4[21:20]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_18 = {sourceDataVec_7[21:20], sourceDataVec_6[21:20]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_18 = {maskDestinationResult_lo_lo_hi_hi_18, maskDestinationResult_lo_lo_hi_lo_18};
  wire [15:0]   maskDestinationResult_lo_lo_19 = {maskDestinationResult_lo_lo_hi_18, maskDestinationResult_lo_lo_lo_18};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_18 = {sourceDataVec_9[21:20], sourceDataVec_8[21:20]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_18 = {sourceDataVec_11[21:20], sourceDataVec_10[21:20]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_18 = {maskDestinationResult_lo_hi_lo_hi_18, maskDestinationResult_lo_hi_lo_lo_18};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_18 = {sourceDataVec_13[21:20], sourceDataVec_12[21:20]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_18 = {sourceDataVec_15[21:20], sourceDataVec_14[21:20]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_18 = {maskDestinationResult_lo_hi_hi_hi_18, maskDestinationResult_lo_hi_hi_lo_18};
  wire [15:0]   maskDestinationResult_lo_hi_19 = {maskDestinationResult_lo_hi_hi_18, maskDestinationResult_lo_hi_lo_18};
  wire [31:0]   maskDestinationResult_lo_275 = {maskDestinationResult_lo_hi_19, maskDestinationResult_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_18 = {sourceDataVec_17[21:20], sourceDataVec_16[21:20]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_18 = {sourceDataVec_19[21:20], sourceDataVec_18[21:20]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_18 = {maskDestinationResult_hi_lo_lo_hi_18, maskDestinationResult_hi_lo_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_18 = {sourceDataVec_21[21:20], sourceDataVec_20[21:20]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_18 = {sourceDataVec_23[21:20], sourceDataVec_22[21:20]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_18 = {maskDestinationResult_hi_lo_hi_hi_18, maskDestinationResult_hi_lo_hi_lo_18};
  wire [15:0]   maskDestinationResult_hi_lo_19 = {maskDestinationResult_hi_lo_hi_18, maskDestinationResult_hi_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_18 = {sourceDataVec_25[21:20], sourceDataVec_24[21:20]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_18 = {sourceDataVec_27[21:20], sourceDataVec_26[21:20]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_18 = {maskDestinationResult_hi_hi_lo_hi_18, maskDestinationResult_hi_hi_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_18 = {sourceDataVec_29[21:20], sourceDataVec_28[21:20]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_18 = {sourceDataVec_31[21:20], sourceDataVec_30[21:20]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_18 = {maskDestinationResult_hi_hi_hi_hi_18, maskDestinationResult_hi_hi_hi_lo_18};
  wire [15:0]   maskDestinationResult_hi_hi_19 = {maskDestinationResult_hi_hi_hi_18, maskDestinationResult_hi_hi_lo_18};
  wire [31:0]   maskDestinationResult_hi_275 = {maskDestinationResult_hi_hi_19, maskDestinationResult_hi_lo_19};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_19 = {sourceDataVec_1[23:22], sourceDataVec_0[23:22]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_19 = {sourceDataVec_3[23:22], sourceDataVec_2[23:22]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_19 = {maskDestinationResult_lo_lo_lo_hi_19, maskDestinationResult_lo_lo_lo_lo_19};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_19 = {sourceDataVec_5[23:22], sourceDataVec_4[23:22]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_19 = {sourceDataVec_7[23:22], sourceDataVec_6[23:22]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_19 = {maskDestinationResult_lo_lo_hi_hi_19, maskDestinationResult_lo_lo_hi_lo_19};
  wire [15:0]   maskDestinationResult_lo_lo_20 = {maskDestinationResult_lo_lo_hi_19, maskDestinationResult_lo_lo_lo_19};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_19 = {sourceDataVec_9[23:22], sourceDataVec_8[23:22]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_19 = {sourceDataVec_11[23:22], sourceDataVec_10[23:22]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_19 = {maskDestinationResult_lo_hi_lo_hi_19, maskDestinationResult_lo_hi_lo_lo_19};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_19 = {sourceDataVec_13[23:22], sourceDataVec_12[23:22]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_19 = {sourceDataVec_15[23:22], sourceDataVec_14[23:22]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_19 = {maskDestinationResult_lo_hi_hi_hi_19, maskDestinationResult_lo_hi_hi_lo_19};
  wire [15:0]   maskDestinationResult_lo_hi_20 = {maskDestinationResult_lo_hi_hi_19, maskDestinationResult_lo_hi_lo_19};
  wire [31:0]   maskDestinationResult_lo_276 = {maskDestinationResult_lo_hi_20, maskDestinationResult_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_19 = {sourceDataVec_17[23:22], sourceDataVec_16[23:22]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_19 = {sourceDataVec_19[23:22], sourceDataVec_18[23:22]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_19 = {maskDestinationResult_hi_lo_lo_hi_19, maskDestinationResult_hi_lo_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_19 = {sourceDataVec_21[23:22], sourceDataVec_20[23:22]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_19 = {sourceDataVec_23[23:22], sourceDataVec_22[23:22]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_19 = {maskDestinationResult_hi_lo_hi_hi_19, maskDestinationResult_hi_lo_hi_lo_19};
  wire [15:0]   maskDestinationResult_hi_lo_20 = {maskDestinationResult_hi_lo_hi_19, maskDestinationResult_hi_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_19 = {sourceDataVec_25[23:22], sourceDataVec_24[23:22]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_19 = {sourceDataVec_27[23:22], sourceDataVec_26[23:22]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_19 = {maskDestinationResult_hi_hi_lo_hi_19, maskDestinationResult_hi_hi_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_19 = {sourceDataVec_29[23:22], sourceDataVec_28[23:22]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_19 = {sourceDataVec_31[23:22], sourceDataVec_30[23:22]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_19 = {maskDestinationResult_hi_hi_hi_hi_19, maskDestinationResult_hi_hi_hi_lo_19};
  wire [15:0]   maskDestinationResult_hi_hi_20 = {maskDestinationResult_hi_hi_hi_19, maskDestinationResult_hi_hi_lo_19};
  wire [31:0]   maskDestinationResult_hi_276 = {maskDestinationResult_hi_hi_20, maskDestinationResult_hi_lo_20};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_20 = {sourceDataVec_1[25:24], sourceDataVec_0[25:24]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_20 = {sourceDataVec_3[25:24], sourceDataVec_2[25:24]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_20 = {maskDestinationResult_lo_lo_lo_hi_20, maskDestinationResult_lo_lo_lo_lo_20};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_20 = {sourceDataVec_5[25:24], sourceDataVec_4[25:24]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_20 = {sourceDataVec_7[25:24], sourceDataVec_6[25:24]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_20 = {maskDestinationResult_lo_lo_hi_hi_20, maskDestinationResult_lo_lo_hi_lo_20};
  wire [15:0]   maskDestinationResult_lo_lo_21 = {maskDestinationResult_lo_lo_hi_20, maskDestinationResult_lo_lo_lo_20};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_20 = {sourceDataVec_9[25:24], sourceDataVec_8[25:24]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_20 = {sourceDataVec_11[25:24], sourceDataVec_10[25:24]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_20 = {maskDestinationResult_lo_hi_lo_hi_20, maskDestinationResult_lo_hi_lo_lo_20};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_20 = {sourceDataVec_13[25:24], sourceDataVec_12[25:24]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_20 = {sourceDataVec_15[25:24], sourceDataVec_14[25:24]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_20 = {maskDestinationResult_lo_hi_hi_hi_20, maskDestinationResult_lo_hi_hi_lo_20};
  wire [15:0]   maskDestinationResult_lo_hi_21 = {maskDestinationResult_lo_hi_hi_20, maskDestinationResult_lo_hi_lo_20};
  wire [31:0]   maskDestinationResult_lo_277 = {maskDestinationResult_lo_hi_21, maskDestinationResult_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_20 = {sourceDataVec_17[25:24], sourceDataVec_16[25:24]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_20 = {sourceDataVec_19[25:24], sourceDataVec_18[25:24]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_20 = {maskDestinationResult_hi_lo_lo_hi_20, maskDestinationResult_hi_lo_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_20 = {sourceDataVec_21[25:24], sourceDataVec_20[25:24]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_20 = {sourceDataVec_23[25:24], sourceDataVec_22[25:24]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_20 = {maskDestinationResult_hi_lo_hi_hi_20, maskDestinationResult_hi_lo_hi_lo_20};
  wire [15:0]   maskDestinationResult_hi_lo_21 = {maskDestinationResult_hi_lo_hi_20, maskDestinationResult_hi_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_20 = {sourceDataVec_25[25:24], sourceDataVec_24[25:24]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_20 = {sourceDataVec_27[25:24], sourceDataVec_26[25:24]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_20 = {maskDestinationResult_hi_hi_lo_hi_20, maskDestinationResult_hi_hi_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_20 = {sourceDataVec_29[25:24], sourceDataVec_28[25:24]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_20 = {sourceDataVec_31[25:24], sourceDataVec_30[25:24]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_20 = {maskDestinationResult_hi_hi_hi_hi_20, maskDestinationResult_hi_hi_hi_lo_20};
  wire [15:0]   maskDestinationResult_hi_hi_21 = {maskDestinationResult_hi_hi_hi_20, maskDestinationResult_hi_hi_lo_20};
  wire [31:0]   maskDestinationResult_hi_277 = {maskDestinationResult_hi_hi_21, maskDestinationResult_hi_lo_21};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_21 = {sourceDataVec_1[27:26], sourceDataVec_0[27:26]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_21 = {sourceDataVec_3[27:26], sourceDataVec_2[27:26]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_21 = {maskDestinationResult_lo_lo_lo_hi_21, maskDestinationResult_lo_lo_lo_lo_21};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_21 = {sourceDataVec_5[27:26], sourceDataVec_4[27:26]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_21 = {sourceDataVec_7[27:26], sourceDataVec_6[27:26]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_21 = {maskDestinationResult_lo_lo_hi_hi_21, maskDestinationResult_lo_lo_hi_lo_21};
  wire [15:0]   maskDestinationResult_lo_lo_22 = {maskDestinationResult_lo_lo_hi_21, maskDestinationResult_lo_lo_lo_21};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_21 = {sourceDataVec_9[27:26], sourceDataVec_8[27:26]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_21 = {sourceDataVec_11[27:26], sourceDataVec_10[27:26]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_21 = {maskDestinationResult_lo_hi_lo_hi_21, maskDestinationResult_lo_hi_lo_lo_21};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_21 = {sourceDataVec_13[27:26], sourceDataVec_12[27:26]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_21 = {sourceDataVec_15[27:26], sourceDataVec_14[27:26]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_21 = {maskDestinationResult_lo_hi_hi_hi_21, maskDestinationResult_lo_hi_hi_lo_21};
  wire [15:0]   maskDestinationResult_lo_hi_22 = {maskDestinationResult_lo_hi_hi_21, maskDestinationResult_lo_hi_lo_21};
  wire [31:0]   maskDestinationResult_lo_278 = {maskDestinationResult_lo_hi_22, maskDestinationResult_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_21 = {sourceDataVec_17[27:26], sourceDataVec_16[27:26]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_21 = {sourceDataVec_19[27:26], sourceDataVec_18[27:26]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_21 = {maskDestinationResult_hi_lo_lo_hi_21, maskDestinationResult_hi_lo_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_21 = {sourceDataVec_21[27:26], sourceDataVec_20[27:26]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_21 = {sourceDataVec_23[27:26], sourceDataVec_22[27:26]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_21 = {maskDestinationResult_hi_lo_hi_hi_21, maskDestinationResult_hi_lo_hi_lo_21};
  wire [15:0]   maskDestinationResult_hi_lo_22 = {maskDestinationResult_hi_lo_hi_21, maskDestinationResult_hi_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_21 = {sourceDataVec_25[27:26], sourceDataVec_24[27:26]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_21 = {sourceDataVec_27[27:26], sourceDataVec_26[27:26]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_21 = {maskDestinationResult_hi_hi_lo_hi_21, maskDestinationResult_hi_hi_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_21 = {sourceDataVec_29[27:26], sourceDataVec_28[27:26]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_21 = {sourceDataVec_31[27:26], sourceDataVec_30[27:26]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_21 = {maskDestinationResult_hi_hi_hi_hi_21, maskDestinationResult_hi_hi_hi_lo_21};
  wire [15:0]   maskDestinationResult_hi_hi_22 = {maskDestinationResult_hi_hi_hi_21, maskDestinationResult_hi_hi_lo_21};
  wire [31:0]   maskDestinationResult_hi_278 = {maskDestinationResult_hi_hi_22, maskDestinationResult_hi_lo_22};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_22 = {sourceDataVec_1[29:28], sourceDataVec_0[29:28]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_22 = {sourceDataVec_3[29:28], sourceDataVec_2[29:28]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_22 = {maskDestinationResult_lo_lo_lo_hi_22, maskDestinationResult_lo_lo_lo_lo_22};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_22 = {sourceDataVec_5[29:28], sourceDataVec_4[29:28]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_22 = {sourceDataVec_7[29:28], sourceDataVec_6[29:28]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_22 = {maskDestinationResult_lo_lo_hi_hi_22, maskDestinationResult_lo_lo_hi_lo_22};
  wire [15:0]   maskDestinationResult_lo_lo_23 = {maskDestinationResult_lo_lo_hi_22, maskDestinationResult_lo_lo_lo_22};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_22 = {sourceDataVec_9[29:28], sourceDataVec_8[29:28]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_22 = {sourceDataVec_11[29:28], sourceDataVec_10[29:28]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_22 = {maskDestinationResult_lo_hi_lo_hi_22, maskDestinationResult_lo_hi_lo_lo_22};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_22 = {sourceDataVec_13[29:28], sourceDataVec_12[29:28]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_22 = {sourceDataVec_15[29:28], sourceDataVec_14[29:28]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_22 = {maskDestinationResult_lo_hi_hi_hi_22, maskDestinationResult_lo_hi_hi_lo_22};
  wire [15:0]   maskDestinationResult_lo_hi_23 = {maskDestinationResult_lo_hi_hi_22, maskDestinationResult_lo_hi_lo_22};
  wire [31:0]   maskDestinationResult_lo_279 = {maskDestinationResult_lo_hi_23, maskDestinationResult_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_22 = {sourceDataVec_17[29:28], sourceDataVec_16[29:28]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_22 = {sourceDataVec_19[29:28], sourceDataVec_18[29:28]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_22 = {maskDestinationResult_hi_lo_lo_hi_22, maskDestinationResult_hi_lo_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_22 = {sourceDataVec_21[29:28], sourceDataVec_20[29:28]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_22 = {sourceDataVec_23[29:28], sourceDataVec_22[29:28]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_22 = {maskDestinationResult_hi_lo_hi_hi_22, maskDestinationResult_hi_lo_hi_lo_22};
  wire [15:0]   maskDestinationResult_hi_lo_23 = {maskDestinationResult_hi_lo_hi_22, maskDestinationResult_hi_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_22 = {sourceDataVec_25[29:28], sourceDataVec_24[29:28]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_22 = {sourceDataVec_27[29:28], sourceDataVec_26[29:28]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_22 = {maskDestinationResult_hi_hi_lo_hi_22, maskDestinationResult_hi_hi_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_22 = {sourceDataVec_29[29:28], sourceDataVec_28[29:28]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_22 = {sourceDataVec_31[29:28], sourceDataVec_30[29:28]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_22 = {maskDestinationResult_hi_hi_hi_hi_22, maskDestinationResult_hi_hi_hi_lo_22};
  wire [15:0]   maskDestinationResult_hi_hi_23 = {maskDestinationResult_hi_hi_hi_22, maskDestinationResult_hi_hi_lo_22};
  wire [31:0]   maskDestinationResult_hi_279 = {maskDestinationResult_hi_hi_23, maskDestinationResult_hi_lo_23};
  wire [3:0]    maskDestinationResult_lo_lo_lo_lo_23 = {sourceDataVec_1[31:30], sourceDataVec_0[31:30]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_hi_23 = {sourceDataVec_3[31:30], sourceDataVec_2[31:30]};
  wire [7:0]    maskDestinationResult_lo_lo_lo_23 = {maskDestinationResult_lo_lo_lo_hi_23, maskDestinationResult_lo_lo_lo_lo_23};
  wire [3:0]    maskDestinationResult_lo_lo_hi_lo_23 = {sourceDataVec_5[31:30], sourceDataVec_4[31:30]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_hi_23 = {sourceDataVec_7[31:30], sourceDataVec_6[31:30]};
  wire [7:0]    maskDestinationResult_lo_lo_hi_23 = {maskDestinationResult_lo_lo_hi_hi_23, maskDestinationResult_lo_lo_hi_lo_23};
  wire [15:0]   maskDestinationResult_lo_lo_24 = {maskDestinationResult_lo_lo_hi_23, maskDestinationResult_lo_lo_lo_23};
  wire [3:0]    maskDestinationResult_lo_hi_lo_lo_23 = {sourceDataVec_9[31:30], sourceDataVec_8[31:30]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_hi_23 = {sourceDataVec_11[31:30], sourceDataVec_10[31:30]};
  wire [7:0]    maskDestinationResult_lo_hi_lo_23 = {maskDestinationResult_lo_hi_lo_hi_23, maskDestinationResult_lo_hi_lo_lo_23};
  wire [3:0]    maskDestinationResult_lo_hi_hi_lo_23 = {sourceDataVec_13[31:30], sourceDataVec_12[31:30]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_hi_23 = {sourceDataVec_15[31:30], sourceDataVec_14[31:30]};
  wire [7:0]    maskDestinationResult_lo_hi_hi_23 = {maskDestinationResult_lo_hi_hi_hi_23, maskDestinationResult_lo_hi_hi_lo_23};
  wire [15:0]   maskDestinationResult_lo_hi_24 = {maskDestinationResult_lo_hi_hi_23, maskDestinationResult_lo_hi_lo_23};
  wire [31:0]   maskDestinationResult_lo_280 = {maskDestinationResult_lo_hi_24, maskDestinationResult_lo_lo_24};
  wire [3:0]    maskDestinationResult_hi_lo_lo_lo_23 = {sourceDataVec_17[31:30], sourceDataVec_16[31:30]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_hi_23 = {sourceDataVec_19[31:30], sourceDataVec_18[31:30]};
  wire [7:0]    maskDestinationResult_hi_lo_lo_23 = {maskDestinationResult_hi_lo_lo_hi_23, maskDestinationResult_hi_lo_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_lo_hi_lo_23 = {sourceDataVec_21[31:30], sourceDataVec_20[31:30]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_hi_23 = {sourceDataVec_23[31:30], sourceDataVec_22[31:30]};
  wire [7:0]    maskDestinationResult_hi_lo_hi_23 = {maskDestinationResult_hi_lo_hi_hi_23, maskDestinationResult_hi_lo_hi_lo_23};
  wire [15:0]   maskDestinationResult_hi_lo_24 = {maskDestinationResult_hi_lo_hi_23, maskDestinationResult_hi_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_hi_lo_lo_23 = {sourceDataVec_25[31:30], sourceDataVec_24[31:30]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_hi_23 = {sourceDataVec_27[31:30], sourceDataVec_26[31:30]};
  wire [7:0]    maskDestinationResult_hi_hi_lo_23 = {maskDestinationResult_hi_hi_lo_hi_23, maskDestinationResult_hi_hi_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_hi_hi_lo_23 = {sourceDataVec_29[31:30], sourceDataVec_28[31:30]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_hi_23 = {sourceDataVec_31[31:30], sourceDataVec_30[31:30]};
  wire [7:0]    maskDestinationResult_hi_hi_hi_23 = {maskDestinationResult_hi_hi_hi_hi_23, maskDestinationResult_hi_hi_hi_lo_23};
  wire [15:0]   maskDestinationResult_hi_hi_24 = {maskDestinationResult_hi_hi_hi_23, maskDestinationResult_hi_hi_lo_23};
  wire [31:0]   maskDestinationResult_hi_280 = {maskDestinationResult_hi_hi_24, maskDestinationResult_hi_lo_24};
  wire [127:0]  maskDestinationResult_lo_lo_lo_24 = {maskDestinationResult_hi_266, maskDestinationResult_lo_266, maskDestinationResult_hi_265, maskDestinationResult_lo_265};
  wire [127:0]  maskDestinationResult_lo_lo_hi_24 = {maskDestinationResult_hi_268, maskDestinationResult_lo_268, maskDestinationResult_hi_267, maskDestinationResult_lo_267};
  wire [255:0]  maskDestinationResult_lo_lo_25 = {maskDestinationResult_lo_lo_hi_24, maskDestinationResult_lo_lo_lo_24};
  wire [127:0]  maskDestinationResult_lo_hi_lo_24 = {maskDestinationResult_hi_270, maskDestinationResult_lo_270, maskDestinationResult_hi_269, maskDestinationResult_lo_269};
  wire [127:0]  maskDestinationResult_lo_hi_hi_24 = {maskDestinationResult_hi_272, maskDestinationResult_lo_272, maskDestinationResult_hi_271, maskDestinationResult_lo_271};
  wire [255:0]  maskDestinationResult_lo_hi_25 = {maskDestinationResult_lo_hi_hi_24, maskDestinationResult_lo_hi_lo_24};
  wire [511:0]  maskDestinationResult_lo_281 = {maskDestinationResult_lo_hi_25, maskDestinationResult_lo_lo_25};
  wire [127:0]  maskDestinationResult_hi_lo_lo_24 = {maskDestinationResult_hi_274, maskDestinationResult_lo_274, maskDestinationResult_hi_273, maskDestinationResult_lo_273};
  wire [127:0]  maskDestinationResult_hi_lo_hi_24 = {maskDestinationResult_hi_276, maskDestinationResult_lo_276, maskDestinationResult_hi_275, maskDestinationResult_lo_275};
  wire [255:0]  maskDestinationResult_hi_lo_25 = {maskDestinationResult_hi_lo_hi_24, maskDestinationResult_hi_lo_lo_24};
  wire [127:0]  maskDestinationResult_hi_hi_lo_24 = {maskDestinationResult_hi_278, maskDestinationResult_lo_278, maskDestinationResult_hi_277, maskDestinationResult_lo_277};
  wire [127:0]  maskDestinationResult_hi_hi_hi_24 = {maskDestinationResult_hi_280, maskDestinationResult_lo_280, maskDestinationResult_hi_279, maskDestinationResult_lo_279};
  wire [255:0]  maskDestinationResult_hi_hi_25 = {maskDestinationResult_hi_hi_hi_24, maskDestinationResult_hi_hi_lo_24};
  wire [511:0]  maskDestinationResult_hi_281 = {maskDestinationResult_hi_hi_25, maskDestinationResult_hi_lo_25};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_24 = {sourceDataVec_1[0], sourceDataVec_0[0]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_24 = {sourceDataVec_3[0], sourceDataVec_2[0]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_25 = {maskDestinationResult_lo_lo_lo_hi_24, maskDestinationResult_lo_lo_lo_lo_24};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_24 = {sourceDataVec_5[0], sourceDataVec_4[0]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_24 = {sourceDataVec_7[0], sourceDataVec_6[0]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_25 = {maskDestinationResult_lo_lo_hi_hi_24, maskDestinationResult_lo_lo_hi_lo_24};
  wire [7:0]    maskDestinationResult_lo_lo_26 = {maskDestinationResult_lo_lo_hi_25, maskDestinationResult_lo_lo_lo_25};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_24 = {sourceDataVec_9[0], sourceDataVec_8[0]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_24 = {sourceDataVec_11[0], sourceDataVec_10[0]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_25 = {maskDestinationResult_lo_hi_lo_hi_24, maskDestinationResult_lo_hi_lo_lo_24};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_24 = {sourceDataVec_13[0], sourceDataVec_12[0]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_24 = {sourceDataVec_15[0], sourceDataVec_14[0]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_25 = {maskDestinationResult_lo_hi_hi_hi_24, maskDestinationResult_lo_hi_hi_lo_24};
  wire [7:0]    maskDestinationResult_lo_hi_26 = {maskDestinationResult_lo_hi_hi_25, maskDestinationResult_lo_hi_lo_25};
  wire [15:0]   maskDestinationResult_lo_282 = {maskDestinationResult_lo_hi_26, maskDestinationResult_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_24 = {sourceDataVec_17[0], sourceDataVec_16[0]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_24 = {sourceDataVec_19[0], sourceDataVec_18[0]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_25 = {maskDestinationResult_hi_lo_lo_hi_24, maskDestinationResult_hi_lo_lo_lo_24};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_24 = {sourceDataVec_21[0], sourceDataVec_20[0]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_24 = {sourceDataVec_23[0], sourceDataVec_22[0]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_25 = {maskDestinationResult_hi_lo_hi_hi_24, maskDestinationResult_hi_lo_hi_lo_24};
  wire [7:0]    maskDestinationResult_hi_lo_26 = {maskDestinationResult_hi_lo_hi_25, maskDestinationResult_hi_lo_lo_25};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_24 = {sourceDataVec_25[0], sourceDataVec_24[0]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_24 = {sourceDataVec_27[0], sourceDataVec_26[0]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_25 = {maskDestinationResult_hi_hi_lo_hi_24, maskDestinationResult_hi_hi_lo_lo_24};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_24 = {sourceDataVec_29[0], sourceDataVec_28[0]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_24 = {sourceDataVec_31[0], sourceDataVec_30[0]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_25 = {maskDestinationResult_hi_hi_hi_hi_24, maskDestinationResult_hi_hi_hi_lo_24};
  wire [7:0]    maskDestinationResult_hi_hi_26 = {maskDestinationResult_hi_hi_hi_25, maskDestinationResult_hi_hi_lo_25};
  wire [15:0]   maskDestinationResult_hi_282 = {maskDestinationResult_hi_hi_26, maskDestinationResult_hi_lo_26};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_25 = {sourceDataVec_1[1], sourceDataVec_0[1]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_25 = {sourceDataVec_3[1], sourceDataVec_2[1]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_26 = {maskDestinationResult_lo_lo_lo_hi_25, maskDestinationResult_lo_lo_lo_lo_25};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_25 = {sourceDataVec_5[1], sourceDataVec_4[1]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_25 = {sourceDataVec_7[1], sourceDataVec_6[1]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_26 = {maskDestinationResult_lo_lo_hi_hi_25, maskDestinationResult_lo_lo_hi_lo_25};
  wire [7:0]    maskDestinationResult_lo_lo_27 = {maskDestinationResult_lo_lo_hi_26, maskDestinationResult_lo_lo_lo_26};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_25 = {sourceDataVec_9[1], sourceDataVec_8[1]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_25 = {sourceDataVec_11[1], sourceDataVec_10[1]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_26 = {maskDestinationResult_lo_hi_lo_hi_25, maskDestinationResult_lo_hi_lo_lo_25};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_25 = {sourceDataVec_13[1], sourceDataVec_12[1]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_25 = {sourceDataVec_15[1], sourceDataVec_14[1]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_26 = {maskDestinationResult_lo_hi_hi_hi_25, maskDestinationResult_lo_hi_hi_lo_25};
  wire [7:0]    maskDestinationResult_lo_hi_27 = {maskDestinationResult_lo_hi_hi_26, maskDestinationResult_lo_hi_lo_26};
  wire [15:0]   maskDestinationResult_lo_283 = {maskDestinationResult_lo_hi_27, maskDestinationResult_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_25 = {sourceDataVec_17[1], sourceDataVec_16[1]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_25 = {sourceDataVec_19[1], sourceDataVec_18[1]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_26 = {maskDestinationResult_hi_lo_lo_hi_25, maskDestinationResult_hi_lo_lo_lo_25};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_25 = {sourceDataVec_21[1], sourceDataVec_20[1]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_25 = {sourceDataVec_23[1], sourceDataVec_22[1]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_26 = {maskDestinationResult_hi_lo_hi_hi_25, maskDestinationResult_hi_lo_hi_lo_25};
  wire [7:0]    maskDestinationResult_hi_lo_27 = {maskDestinationResult_hi_lo_hi_26, maskDestinationResult_hi_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_25 = {sourceDataVec_25[1], sourceDataVec_24[1]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_25 = {sourceDataVec_27[1], sourceDataVec_26[1]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_26 = {maskDestinationResult_hi_hi_lo_hi_25, maskDestinationResult_hi_hi_lo_lo_25};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_25 = {sourceDataVec_29[1], sourceDataVec_28[1]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_25 = {sourceDataVec_31[1], sourceDataVec_30[1]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_26 = {maskDestinationResult_hi_hi_hi_hi_25, maskDestinationResult_hi_hi_hi_lo_25};
  wire [7:0]    maskDestinationResult_hi_hi_27 = {maskDestinationResult_hi_hi_hi_26, maskDestinationResult_hi_hi_lo_26};
  wire [15:0]   maskDestinationResult_hi_283 = {maskDestinationResult_hi_hi_27, maskDestinationResult_hi_lo_27};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_26 = {sourceDataVec_1[2], sourceDataVec_0[2]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_26 = {sourceDataVec_3[2], sourceDataVec_2[2]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_27 = {maskDestinationResult_lo_lo_lo_hi_26, maskDestinationResult_lo_lo_lo_lo_26};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_26 = {sourceDataVec_5[2], sourceDataVec_4[2]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_26 = {sourceDataVec_7[2], sourceDataVec_6[2]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_27 = {maskDestinationResult_lo_lo_hi_hi_26, maskDestinationResult_lo_lo_hi_lo_26};
  wire [7:0]    maskDestinationResult_lo_lo_28 = {maskDestinationResult_lo_lo_hi_27, maskDestinationResult_lo_lo_lo_27};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_26 = {sourceDataVec_9[2], sourceDataVec_8[2]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_26 = {sourceDataVec_11[2], sourceDataVec_10[2]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_27 = {maskDestinationResult_lo_hi_lo_hi_26, maskDestinationResult_lo_hi_lo_lo_26};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_26 = {sourceDataVec_13[2], sourceDataVec_12[2]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_26 = {sourceDataVec_15[2], sourceDataVec_14[2]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_27 = {maskDestinationResult_lo_hi_hi_hi_26, maskDestinationResult_lo_hi_hi_lo_26};
  wire [7:0]    maskDestinationResult_lo_hi_28 = {maskDestinationResult_lo_hi_hi_27, maskDestinationResult_lo_hi_lo_27};
  wire [15:0]   maskDestinationResult_lo_284 = {maskDestinationResult_lo_hi_28, maskDestinationResult_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_26 = {sourceDataVec_17[2], sourceDataVec_16[2]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_26 = {sourceDataVec_19[2], sourceDataVec_18[2]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_27 = {maskDestinationResult_hi_lo_lo_hi_26, maskDestinationResult_hi_lo_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_26 = {sourceDataVec_21[2], sourceDataVec_20[2]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_26 = {sourceDataVec_23[2], sourceDataVec_22[2]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_27 = {maskDestinationResult_hi_lo_hi_hi_26, maskDestinationResult_hi_lo_hi_lo_26};
  wire [7:0]    maskDestinationResult_hi_lo_28 = {maskDestinationResult_hi_lo_hi_27, maskDestinationResult_hi_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_26 = {sourceDataVec_25[2], sourceDataVec_24[2]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_26 = {sourceDataVec_27[2], sourceDataVec_26[2]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_27 = {maskDestinationResult_hi_hi_lo_hi_26, maskDestinationResult_hi_hi_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_26 = {sourceDataVec_29[2], sourceDataVec_28[2]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_26 = {sourceDataVec_31[2], sourceDataVec_30[2]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_27 = {maskDestinationResult_hi_hi_hi_hi_26, maskDestinationResult_hi_hi_hi_lo_26};
  wire [7:0]    maskDestinationResult_hi_hi_28 = {maskDestinationResult_hi_hi_hi_27, maskDestinationResult_hi_hi_lo_27};
  wire [15:0]   maskDestinationResult_hi_284 = {maskDestinationResult_hi_hi_28, maskDestinationResult_hi_lo_28};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_27 = {sourceDataVec_1[3], sourceDataVec_0[3]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_27 = {sourceDataVec_3[3], sourceDataVec_2[3]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_28 = {maskDestinationResult_lo_lo_lo_hi_27, maskDestinationResult_lo_lo_lo_lo_27};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_27 = {sourceDataVec_5[3], sourceDataVec_4[3]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_27 = {sourceDataVec_7[3], sourceDataVec_6[3]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_28 = {maskDestinationResult_lo_lo_hi_hi_27, maskDestinationResult_lo_lo_hi_lo_27};
  wire [7:0]    maskDestinationResult_lo_lo_29 = {maskDestinationResult_lo_lo_hi_28, maskDestinationResult_lo_lo_lo_28};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_27 = {sourceDataVec_9[3], sourceDataVec_8[3]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_27 = {sourceDataVec_11[3], sourceDataVec_10[3]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_28 = {maskDestinationResult_lo_hi_lo_hi_27, maskDestinationResult_lo_hi_lo_lo_27};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_27 = {sourceDataVec_13[3], sourceDataVec_12[3]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_27 = {sourceDataVec_15[3], sourceDataVec_14[3]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_28 = {maskDestinationResult_lo_hi_hi_hi_27, maskDestinationResult_lo_hi_hi_lo_27};
  wire [7:0]    maskDestinationResult_lo_hi_29 = {maskDestinationResult_lo_hi_hi_28, maskDestinationResult_lo_hi_lo_28};
  wire [15:0]   maskDestinationResult_lo_285 = {maskDestinationResult_lo_hi_29, maskDestinationResult_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_27 = {sourceDataVec_17[3], sourceDataVec_16[3]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_27 = {sourceDataVec_19[3], sourceDataVec_18[3]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_28 = {maskDestinationResult_hi_lo_lo_hi_27, maskDestinationResult_hi_lo_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_27 = {sourceDataVec_21[3], sourceDataVec_20[3]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_27 = {sourceDataVec_23[3], sourceDataVec_22[3]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_28 = {maskDestinationResult_hi_lo_hi_hi_27, maskDestinationResult_hi_lo_hi_lo_27};
  wire [7:0]    maskDestinationResult_hi_lo_29 = {maskDestinationResult_hi_lo_hi_28, maskDestinationResult_hi_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_27 = {sourceDataVec_25[3], sourceDataVec_24[3]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_27 = {sourceDataVec_27[3], sourceDataVec_26[3]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_28 = {maskDestinationResult_hi_hi_lo_hi_27, maskDestinationResult_hi_hi_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_27 = {sourceDataVec_29[3], sourceDataVec_28[3]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_27 = {sourceDataVec_31[3], sourceDataVec_30[3]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_28 = {maskDestinationResult_hi_hi_hi_hi_27, maskDestinationResult_hi_hi_hi_lo_27};
  wire [7:0]    maskDestinationResult_hi_hi_29 = {maskDestinationResult_hi_hi_hi_28, maskDestinationResult_hi_hi_lo_28};
  wire [15:0]   maskDestinationResult_hi_285 = {maskDestinationResult_hi_hi_29, maskDestinationResult_hi_lo_29};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_28 = {sourceDataVec_1[4], sourceDataVec_0[4]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_28 = {sourceDataVec_3[4], sourceDataVec_2[4]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_29 = {maskDestinationResult_lo_lo_lo_hi_28, maskDestinationResult_lo_lo_lo_lo_28};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_28 = {sourceDataVec_5[4], sourceDataVec_4[4]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_28 = {sourceDataVec_7[4], sourceDataVec_6[4]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_29 = {maskDestinationResult_lo_lo_hi_hi_28, maskDestinationResult_lo_lo_hi_lo_28};
  wire [7:0]    maskDestinationResult_lo_lo_30 = {maskDestinationResult_lo_lo_hi_29, maskDestinationResult_lo_lo_lo_29};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_28 = {sourceDataVec_9[4], sourceDataVec_8[4]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_28 = {sourceDataVec_11[4], sourceDataVec_10[4]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_29 = {maskDestinationResult_lo_hi_lo_hi_28, maskDestinationResult_lo_hi_lo_lo_28};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_28 = {sourceDataVec_13[4], sourceDataVec_12[4]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_28 = {sourceDataVec_15[4], sourceDataVec_14[4]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_29 = {maskDestinationResult_lo_hi_hi_hi_28, maskDestinationResult_lo_hi_hi_lo_28};
  wire [7:0]    maskDestinationResult_lo_hi_30 = {maskDestinationResult_lo_hi_hi_29, maskDestinationResult_lo_hi_lo_29};
  wire [15:0]   maskDestinationResult_lo_286 = {maskDestinationResult_lo_hi_30, maskDestinationResult_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_28 = {sourceDataVec_17[4], sourceDataVec_16[4]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_28 = {sourceDataVec_19[4], sourceDataVec_18[4]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_29 = {maskDestinationResult_hi_lo_lo_hi_28, maskDestinationResult_hi_lo_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_28 = {sourceDataVec_21[4], sourceDataVec_20[4]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_28 = {sourceDataVec_23[4], sourceDataVec_22[4]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_29 = {maskDestinationResult_hi_lo_hi_hi_28, maskDestinationResult_hi_lo_hi_lo_28};
  wire [7:0]    maskDestinationResult_hi_lo_30 = {maskDestinationResult_hi_lo_hi_29, maskDestinationResult_hi_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_28 = {sourceDataVec_25[4], sourceDataVec_24[4]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_28 = {sourceDataVec_27[4], sourceDataVec_26[4]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_29 = {maskDestinationResult_hi_hi_lo_hi_28, maskDestinationResult_hi_hi_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_28 = {sourceDataVec_29[4], sourceDataVec_28[4]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_28 = {sourceDataVec_31[4], sourceDataVec_30[4]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_29 = {maskDestinationResult_hi_hi_hi_hi_28, maskDestinationResult_hi_hi_hi_lo_28};
  wire [7:0]    maskDestinationResult_hi_hi_30 = {maskDestinationResult_hi_hi_hi_29, maskDestinationResult_hi_hi_lo_29};
  wire [15:0]   maskDestinationResult_hi_286 = {maskDestinationResult_hi_hi_30, maskDestinationResult_hi_lo_30};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_29 = {sourceDataVec_1[5], sourceDataVec_0[5]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_29 = {sourceDataVec_3[5], sourceDataVec_2[5]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_30 = {maskDestinationResult_lo_lo_lo_hi_29, maskDestinationResult_lo_lo_lo_lo_29};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_29 = {sourceDataVec_5[5], sourceDataVec_4[5]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_29 = {sourceDataVec_7[5], sourceDataVec_6[5]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_30 = {maskDestinationResult_lo_lo_hi_hi_29, maskDestinationResult_lo_lo_hi_lo_29};
  wire [7:0]    maskDestinationResult_lo_lo_31 = {maskDestinationResult_lo_lo_hi_30, maskDestinationResult_lo_lo_lo_30};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_29 = {sourceDataVec_9[5], sourceDataVec_8[5]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_29 = {sourceDataVec_11[5], sourceDataVec_10[5]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_30 = {maskDestinationResult_lo_hi_lo_hi_29, maskDestinationResult_lo_hi_lo_lo_29};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_29 = {sourceDataVec_13[5], sourceDataVec_12[5]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_29 = {sourceDataVec_15[5], sourceDataVec_14[5]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_30 = {maskDestinationResult_lo_hi_hi_hi_29, maskDestinationResult_lo_hi_hi_lo_29};
  wire [7:0]    maskDestinationResult_lo_hi_31 = {maskDestinationResult_lo_hi_hi_30, maskDestinationResult_lo_hi_lo_30};
  wire [15:0]   maskDestinationResult_lo_287 = {maskDestinationResult_lo_hi_31, maskDestinationResult_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_29 = {sourceDataVec_17[5], sourceDataVec_16[5]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_29 = {sourceDataVec_19[5], sourceDataVec_18[5]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_30 = {maskDestinationResult_hi_lo_lo_hi_29, maskDestinationResult_hi_lo_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_29 = {sourceDataVec_21[5], sourceDataVec_20[5]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_29 = {sourceDataVec_23[5], sourceDataVec_22[5]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_30 = {maskDestinationResult_hi_lo_hi_hi_29, maskDestinationResult_hi_lo_hi_lo_29};
  wire [7:0]    maskDestinationResult_hi_lo_31 = {maskDestinationResult_hi_lo_hi_30, maskDestinationResult_hi_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_29 = {sourceDataVec_25[5], sourceDataVec_24[5]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_29 = {sourceDataVec_27[5], sourceDataVec_26[5]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_30 = {maskDestinationResult_hi_hi_lo_hi_29, maskDestinationResult_hi_hi_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_29 = {sourceDataVec_29[5], sourceDataVec_28[5]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_29 = {sourceDataVec_31[5], sourceDataVec_30[5]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_30 = {maskDestinationResult_hi_hi_hi_hi_29, maskDestinationResult_hi_hi_hi_lo_29};
  wire [7:0]    maskDestinationResult_hi_hi_31 = {maskDestinationResult_hi_hi_hi_30, maskDestinationResult_hi_hi_lo_30};
  wire [15:0]   maskDestinationResult_hi_287 = {maskDestinationResult_hi_hi_31, maskDestinationResult_hi_lo_31};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_30 = {sourceDataVec_1[6], sourceDataVec_0[6]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_30 = {sourceDataVec_3[6], sourceDataVec_2[6]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_31 = {maskDestinationResult_lo_lo_lo_hi_30, maskDestinationResult_lo_lo_lo_lo_30};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_30 = {sourceDataVec_5[6], sourceDataVec_4[6]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_30 = {sourceDataVec_7[6], sourceDataVec_6[6]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_31 = {maskDestinationResult_lo_lo_hi_hi_30, maskDestinationResult_lo_lo_hi_lo_30};
  wire [7:0]    maskDestinationResult_lo_lo_32 = {maskDestinationResult_lo_lo_hi_31, maskDestinationResult_lo_lo_lo_31};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_30 = {sourceDataVec_9[6], sourceDataVec_8[6]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_30 = {sourceDataVec_11[6], sourceDataVec_10[6]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_31 = {maskDestinationResult_lo_hi_lo_hi_30, maskDestinationResult_lo_hi_lo_lo_30};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_30 = {sourceDataVec_13[6], sourceDataVec_12[6]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_30 = {sourceDataVec_15[6], sourceDataVec_14[6]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_31 = {maskDestinationResult_lo_hi_hi_hi_30, maskDestinationResult_lo_hi_hi_lo_30};
  wire [7:0]    maskDestinationResult_lo_hi_32 = {maskDestinationResult_lo_hi_hi_31, maskDestinationResult_lo_hi_lo_31};
  wire [15:0]   maskDestinationResult_lo_288 = {maskDestinationResult_lo_hi_32, maskDestinationResult_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_30 = {sourceDataVec_17[6], sourceDataVec_16[6]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_30 = {sourceDataVec_19[6], sourceDataVec_18[6]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_31 = {maskDestinationResult_hi_lo_lo_hi_30, maskDestinationResult_hi_lo_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_30 = {sourceDataVec_21[6], sourceDataVec_20[6]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_30 = {sourceDataVec_23[6], sourceDataVec_22[6]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_31 = {maskDestinationResult_hi_lo_hi_hi_30, maskDestinationResult_hi_lo_hi_lo_30};
  wire [7:0]    maskDestinationResult_hi_lo_32 = {maskDestinationResult_hi_lo_hi_31, maskDestinationResult_hi_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_30 = {sourceDataVec_25[6], sourceDataVec_24[6]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_30 = {sourceDataVec_27[6], sourceDataVec_26[6]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_31 = {maskDestinationResult_hi_hi_lo_hi_30, maskDestinationResult_hi_hi_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_30 = {sourceDataVec_29[6], sourceDataVec_28[6]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_30 = {sourceDataVec_31[6], sourceDataVec_30[6]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_31 = {maskDestinationResult_hi_hi_hi_hi_30, maskDestinationResult_hi_hi_hi_lo_30};
  wire [7:0]    maskDestinationResult_hi_hi_32 = {maskDestinationResult_hi_hi_hi_31, maskDestinationResult_hi_hi_lo_31};
  wire [15:0]   maskDestinationResult_hi_288 = {maskDestinationResult_hi_hi_32, maskDestinationResult_hi_lo_32};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_31 = {sourceDataVec_1[7], sourceDataVec_0[7]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_31 = {sourceDataVec_3[7], sourceDataVec_2[7]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_32 = {maskDestinationResult_lo_lo_lo_hi_31, maskDestinationResult_lo_lo_lo_lo_31};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_31 = {sourceDataVec_5[7], sourceDataVec_4[7]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_31 = {sourceDataVec_7[7], sourceDataVec_6[7]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_32 = {maskDestinationResult_lo_lo_hi_hi_31, maskDestinationResult_lo_lo_hi_lo_31};
  wire [7:0]    maskDestinationResult_lo_lo_33 = {maskDestinationResult_lo_lo_hi_32, maskDestinationResult_lo_lo_lo_32};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_31 = {sourceDataVec_9[7], sourceDataVec_8[7]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_31 = {sourceDataVec_11[7], sourceDataVec_10[7]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_32 = {maskDestinationResult_lo_hi_lo_hi_31, maskDestinationResult_lo_hi_lo_lo_31};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_31 = {sourceDataVec_13[7], sourceDataVec_12[7]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_31 = {sourceDataVec_15[7], sourceDataVec_14[7]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_32 = {maskDestinationResult_lo_hi_hi_hi_31, maskDestinationResult_lo_hi_hi_lo_31};
  wire [7:0]    maskDestinationResult_lo_hi_33 = {maskDestinationResult_lo_hi_hi_32, maskDestinationResult_lo_hi_lo_32};
  wire [15:0]   maskDestinationResult_lo_289 = {maskDestinationResult_lo_hi_33, maskDestinationResult_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_31 = {sourceDataVec_17[7], sourceDataVec_16[7]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_31 = {sourceDataVec_19[7], sourceDataVec_18[7]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_32 = {maskDestinationResult_hi_lo_lo_hi_31, maskDestinationResult_hi_lo_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_31 = {sourceDataVec_21[7], sourceDataVec_20[7]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_31 = {sourceDataVec_23[7], sourceDataVec_22[7]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_32 = {maskDestinationResult_hi_lo_hi_hi_31, maskDestinationResult_hi_lo_hi_lo_31};
  wire [7:0]    maskDestinationResult_hi_lo_33 = {maskDestinationResult_hi_lo_hi_32, maskDestinationResult_hi_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_31 = {sourceDataVec_25[7], sourceDataVec_24[7]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_31 = {sourceDataVec_27[7], sourceDataVec_26[7]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_32 = {maskDestinationResult_hi_hi_lo_hi_31, maskDestinationResult_hi_hi_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_31 = {sourceDataVec_29[7], sourceDataVec_28[7]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_31 = {sourceDataVec_31[7], sourceDataVec_30[7]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_32 = {maskDestinationResult_hi_hi_hi_hi_31, maskDestinationResult_hi_hi_hi_lo_31};
  wire [7:0]    maskDestinationResult_hi_hi_33 = {maskDestinationResult_hi_hi_hi_32, maskDestinationResult_hi_hi_lo_32};
  wire [15:0]   maskDestinationResult_hi_289 = {maskDestinationResult_hi_hi_33, maskDestinationResult_hi_lo_33};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_32 = {sourceDataVec_1[8], sourceDataVec_0[8]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_32 = {sourceDataVec_3[8], sourceDataVec_2[8]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_33 = {maskDestinationResult_lo_lo_lo_hi_32, maskDestinationResult_lo_lo_lo_lo_32};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_32 = {sourceDataVec_5[8], sourceDataVec_4[8]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_32 = {sourceDataVec_7[8], sourceDataVec_6[8]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_33 = {maskDestinationResult_lo_lo_hi_hi_32, maskDestinationResult_lo_lo_hi_lo_32};
  wire [7:0]    maskDestinationResult_lo_lo_34 = {maskDestinationResult_lo_lo_hi_33, maskDestinationResult_lo_lo_lo_33};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_32 = {sourceDataVec_9[8], sourceDataVec_8[8]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_32 = {sourceDataVec_11[8], sourceDataVec_10[8]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_33 = {maskDestinationResult_lo_hi_lo_hi_32, maskDestinationResult_lo_hi_lo_lo_32};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_32 = {sourceDataVec_13[8], sourceDataVec_12[8]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_32 = {sourceDataVec_15[8], sourceDataVec_14[8]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_33 = {maskDestinationResult_lo_hi_hi_hi_32, maskDestinationResult_lo_hi_hi_lo_32};
  wire [7:0]    maskDestinationResult_lo_hi_34 = {maskDestinationResult_lo_hi_hi_33, maskDestinationResult_lo_hi_lo_33};
  wire [15:0]   maskDestinationResult_lo_290 = {maskDestinationResult_lo_hi_34, maskDestinationResult_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_32 = {sourceDataVec_17[8], sourceDataVec_16[8]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_32 = {sourceDataVec_19[8], sourceDataVec_18[8]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_33 = {maskDestinationResult_hi_lo_lo_hi_32, maskDestinationResult_hi_lo_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_32 = {sourceDataVec_21[8], sourceDataVec_20[8]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_32 = {sourceDataVec_23[8], sourceDataVec_22[8]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_33 = {maskDestinationResult_hi_lo_hi_hi_32, maskDestinationResult_hi_lo_hi_lo_32};
  wire [7:0]    maskDestinationResult_hi_lo_34 = {maskDestinationResult_hi_lo_hi_33, maskDestinationResult_hi_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_32 = {sourceDataVec_25[8], sourceDataVec_24[8]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_32 = {sourceDataVec_27[8], sourceDataVec_26[8]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_33 = {maskDestinationResult_hi_hi_lo_hi_32, maskDestinationResult_hi_hi_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_32 = {sourceDataVec_29[8], sourceDataVec_28[8]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_32 = {sourceDataVec_31[8], sourceDataVec_30[8]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_33 = {maskDestinationResult_hi_hi_hi_hi_32, maskDestinationResult_hi_hi_hi_lo_32};
  wire [7:0]    maskDestinationResult_hi_hi_34 = {maskDestinationResult_hi_hi_hi_33, maskDestinationResult_hi_hi_lo_33};
  wire [15:0]   maskDestinationResult_hi_290 = {maskDestinationResult_hi_hi_34, maskDestinationResult_hi_lo_34};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_33 = {sourceDataVec_1[9], sourceDataVec_0[9]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_33 = {sourceDataVec_3[9], sourceDataVec_2[9]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_34 = {maskDestinationResult_lo_lo_lo_hi_33, maskDestinationResult_lo_lo_lo_lo_33};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_33 = {sourceDataVec_5[9], sourceDataVec_4[9]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_33 = {sourceDataVec_7[9], sourceDataVec_6[9]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_34 = {maskDestinationResult_lo_lo_hi_hi_33, maskDestinationResult_lo_lo_hi_lo_33};
  wire [7:0]    maskDestinationResult_lo_lo_35 = {maskDestinationResult_lo_lo_hi_34, maskDestinationResult_lo_lo_lo_34};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_33 = {sourceDataVec_9[9], sourceDataVec_8[9]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_33 = {sourceDataVec_11[9], sourceDataVec_10[9]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_34 = {maskDestinationResult_lo_hi_lo_hi_33, maskDestinationResult_lo_hi_lo_lo_33};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_33 = {sourceDataVec_13[9], sourceDataVec_12[9]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_33 = {sourceDataVec_15[9], sourceDataVec_14[9]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_34 = {maskDestinationResult_lo_hi_hi_hi_33, maskDestinationResult_lo_hi_hi_lo_33};
  wire [7:0]    maskDestinationResult_lo_hi_35 = {maskDestinationResult_lo_hi_hi_34, maskDestinationResult_lo_hi_lo_34};
  wire [15:0]   maskDestinationResult_lo_291 = {maskDestinationResult_lo_hi_35, maskDestinationResult_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_33 = {sourceDataVec_17[9], sourceDataVec_16[9]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_33 = {sourceDataVec_19[9], sourceDataVec_18[9]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_34 = {maskDestinationResult_hi_lo_lo_hi_33, maskDestinationResult_hi_lo_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_33 = {sourceDataVec_21[9], sourceDataVec_20[9]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_33 = {sourceDataVec_23[9], sourceDataVec_22[9]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_34 = {maskDestinationResult_hi_lo_hi_hi_33, maskDestinationResult_hi_lo_hi_lo_33};
  wire [7:0]    maskDestinationResult_hi_lo_35 = {maskDestinationResult_hi_lo_hi_34, maskDestinationResult_hi_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_33 = {sourceDataVec_25[9], sourceDataVec_24[9]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_33 = {sourceDataVec_27[9], sourceDataVec_26[9]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_34 = {maskDestinationResult_hi_hi_lo_hi_33, maskDestinationResult_hi_hi_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_33 = {sourceDataVec_29[9], sourceDataVec_28[9]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_33 = {sourceDataVec_31[9], sourceDataVec_30[9]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_34 = {maskDestinationResult_hi_hi_hi_hi_33, maskDestinationResult_hi_hi_hi_lo_33};
  wire [7:0]    maskDestinationResult_hi_hi_35 = {maskDestinationResult_hi_hi_hi_34, maskDestinationResult_hi_hi_lo_34};
  wire [15:0]   maskDestinationResult_hi_291 = {maskDestinationResult_hi_hi_35, maskDestinationResult_hi_lo_35};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_34 = {sourceDataVec_1[10], sourceDataVec_0[10]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_34 = {sourceDataVec_3[10], sourceDataVec_2[10]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_35 = {maskDestinationResult_lo_lo_lo_hi_34, maskDestinationResult_lo_lo_lo_lo_34};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_34 = {sourceDataVec_5[10], sourceDataVec_4[10]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_34 = {sourceDataVec_7[10], sourceDataVec_6[10]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_35 = {maskDestinationResult_lo_lo_hi_hi_34, maskDestinationResult_lo_lo_hi_lo_34};
  wire [7:0]    maskDestinationResult_lo_lo_36 = {maskDestinationResult_lo_lo_hi_35, maskDestinationResult_lo_lo_lo_35};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_34 = {sourceDataVec_9[10], sourceDataVec_8[10]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_34 = {sourceDataVec_11[10], sourceDataVec_10[10]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_35 = {maskDestinationResult_lo_hi_lo_hi_34, maskDestinationResult_lo_hi_lo_lo_34};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_34 = {sourceDataVec_13[10], sourceDataVec_12[10]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_34 = {sourceDataVec_15[10], sourceDataVec_14[10]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_35 = {maskDestinationResult_lo_hi_hi_hi_34, maskDestinationResult_lo_hi_hi_lo_34};
  wire [7:0]    maskDestinationResult_lo_hi_36 = {maskDestinationResult_lo_hi_hi_35, maskDestinationResult_lo_hi_lo_35};
  wire [15:0]   maskDestinationResult_lo_292 = {maskDestinationResult_lo_hi_36, maskDestinationResult_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_34 = {sourceDataVec_17[10], sourceDataVec_16[10]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_34 = {sourceDataVec_19[10], sourceDataVec_18[10]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_35 = {maskDestinationResult_hi_lo_lo_hi_34, maskDestinationResult_hi_lo_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_34 = {sourceDataVec_21[10], sourceDataVec_20[10]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_34 = {sourceDataVec_23[10], sourceDataVec_22[10]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_35 = {maskDestinationResult_hi_lo_hi_hi_34, maskDestinationResult_hi_lo_hi_lo_34};
  wire [7:0]    maskDestinationResult_hi_lo_36 = {maskDestinationResult_hi_lo_hi_35, maskDestinationResult_hi_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_34 = {sourceDataVec_25[10], sourceDataVec_24[10]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_34 = {sourceDataVec_27[10], sourceDataVec_26[10]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_35 = {maskDestinationResult_hi_hi_lo_hi_34, maskDestinationResult_hi_hi_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_34 = {sourceDataVec_29[10], sourceDataVec_28[10]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_34 = {sourceDataVec_31[10], sourceDataVec_30[10]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_35 = {maskDestinationResult_hi_hi_hi_hi_34, maskDestinationResult_hi_hi_hi_lo_34};
  wire [7:0]    maskDestinationResult_hi_hi_36 = {maskDestinationResult_hi_hi_hi_35, maskDestinationResult_hi_hi_lo_35};
  wire [15:0]   maskDestinationResult_hi_292 = {maskDestinationResult_hi_hi_36, maskDestinationResult_hi_lo_36};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_35 = {sourceDataVec_1[11], sourceDataVec_0[11]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_35 = {sourceDataVec_3[11], sourceDataVec_2[11]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_36 = {maskDestinationResult_lo_lo_lo_hi_35, maskDestinationResult_lo_lo_lo_lo_35};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_35 = {sourceDataVec_5[11], sourceDataVec_4[11]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_35 = {sourceDataVec_7[11], sourceDataVec_6[11]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_36 = {maskDestinationResult_lo_lo_hi_hi_35, maskDestinationResult_lo_lo_hi_lo_35};
  wire [7:0]    maskDestinationResult_lo_lo_37 = {maskDestinationResult_lo_lo_hi_36, maskDestinationResult_lo_lo_lo_36};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_35 = {sourceDataVec_9[11], sourceDataVec_8[11]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_35 = {sourceDataVec_11[11], sourceDataVec_10[11]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_36 = {maskDestinationResult_lo_hi_lo_hi_35, maskDestinationResult_lo_hi_lo_lo_35};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_35 = {sourceDataVec_13[11], sourceDataVec_12[11]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_35 = {sourceDataVec_15[11], sourceDataVec_14[11]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_36 = {maskDestinationResult_lo_hi_hi_hi_35, maskDestinationResult_lo_hi_hi_lo_35};
  wire [7:0]    maskDestinationResult_lo_hi_37 = {maskDestinationResult_lo_hi_hi_36, maskDestinationResult_lo_hi_lo_36};
  wire [15:0]   maskDestinationResult_lo_293 = {maskDestinationResult_lo_hi_37, maskDestinationResult_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_35 = {sourceDataVec_17[11], sourceDataVec_16[11]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_35 = {sourceDataVec_19[11], sourceDataVec_18[11]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_36 = {maskDestinationResult_hi_lo_lo_hi_35, maskDestinationResult_hi_lo_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_35 = {sourceDataVec_21[11], sourceDataVec_20[11]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_35 = {sourceDataVec_23[11], sourceDataVec_22[11]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_36 = {maskDestinationResult_hi_lo_hi_hi_35, maskDestinationResult_hi_lo_hi_lo_35};
  wire [7:0]    maskDestinationResult_hi_lo_37 = {maskDestinationResult_hi_lo_hi_36, maskDestinationResult_hi_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_35 = {sourceDataVec_25[11], sourceDataVec_24[11]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_35 = {sourceDataVec_27[11], sourceDataVec_26[11]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_36 = {maskDestinationResult_hi_hi_lo_hi_35, maskDestinationResult_hi_hi_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_35 = {sourceDataVec_29[11], sourceDataVec_28[11]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_35 = {sourceDataVec_31[11], sourceDataVec_30[11]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_36 = {maskDestinationResult_hi_hi_hi_hi_35, maskDestinationResult_hi_hi_hi_lo_35};
  wire [7:0]    maskDestinationResult_hi_hi_37 = {maskDestinationResult_hi_hi_hi_36, maskDestinationResult_hi_hi_lo_36};
  wire [15:0]   maskDestinationResult_hi_293 = {maskDestinationResult_hi_hi_37, maskDestinationResult_hi_lo_37};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_36 = {sourceDataVec_1[12], sourceDataVec_0[12]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_36 = {sourceDataVec_3[12], sourceDataVec_2[12]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_37 = {maskDestinationResult_lo_lo_lo_hi_36, maskDestinationResult_lo_lo_lo_lo_36};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_36 = {sourceDataVec_5[12], sourceDataVec_4[12]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_36 = {sourceDataVec_7[12], sourceDataVec_6[12]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_37 = {maskDestinationResult_lo_lo_hi_hi_36, maskDestinationResult_lo_lo_hi_lo_36};
  wire [7:0]    maskDestinationResult_lo_lo_38 = {maskDestinationResult_lo_lo_hi_37, maskDestinationResult_lo_lo_lo_37};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_36 = {sourceDataVec_9[12], sourceDataVec_8[12]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_36 = {sourceDataVec_11[12], sourceDataVec_10[12]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_37 = {maskDestinationResult_lo_hi_lo_hi_36, maskDestinationResult_lo_hi_lo_lo_36};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_36 = {sourceDataVec_13[12], sourceDataVec_12[12]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_36 = {sourceDataVec_15[12], sourceDataVec_14[12]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_37 = {maskDestinationResult_lo_hi_hi_hi_36, maskDestinationResult_lo_hi_hi_lo_36};
  wire [7:0]    maskDestinationResult_lo_hi_38 = {maskDestinationResult_lo_hi_hi_37, maskDestinationResult_lo_hi_lo_37};
  wire [15:0]   maskDestinationResult_lo_294 = {maskDestinationResult_lo_hi_38, maskDestinationResult_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_36 = {sourceDataVec_17[12], sourceDataVec_16[12]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_36 = {sourceDataVec_19[12], sourceDataVec_18[12]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_37 = {maskDestinationResult_hi_lo_lo_hi_36, maskDestinationResult_hi_lo_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_36 = {sourceDataVec_21[12], sourceDataVec_20[12]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_36 = {sourceDataVec_23[12], sourceDataVec_22[12]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_37 = {maskDestinationResult_hi_lo_hi_hi_36, maskDestinationResult_hi_lo_hi_lo_36};
  wire [7:0]    maskDestinationResult_hi_lo_38 = {maskDestinationResult_hi_lo_hi_37, maskDestinationResult_hi_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_36 = {sourceDataVec_25[12], sourceDataVec_24[12]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_36 = {sourceDataVec_27[12], sourceDataVec_26[12]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_37 = {maskDestinationResult_hi_hi_lo_hi_36, maskDestinationResult_hi_hi_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_36 = {sourceDataVec_29[12], sourceDataVec_28[12]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_36 = {sourceDataVec_31[12], sourceDataVec_30[12]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_37 = {maskDestinationResult_hi_hi_hi_hi_36, maskDestinationResult_hi_hi_hi_lo_36};
  wire [7:0]    maskDestinationResult_hi_hi_38 = {maskDestinationResult_hi_hi_hi_37, maskDestinationResult_hi_hi_lo_37};
  wire [15:0]   maskDestinationResult_hi_294 = {maskDestinationResult_hi_hi_38, maskDestinationResult_hi_lo_38};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_37 = {sourceDataVec_1[13], sourceDataVec_0[13]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_37 = {sourceDataVec_3[13], sourceDataVec_2[13]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_38 = {maskDestinationResult_lo_lo_lo_hi_37, maskDestinationResult_lo_lo_lo_lo_37};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_37 = {sourceDataVec_5[13], sourceDataVec_4[13]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_37 = {sourceDataVec_7[13], sourceDataVec_6[13]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_38 = {maskDestinationResult_lo_lo_hi_hi_37, maskDestinationResult_lo_lo_hi_lo_37};
  wire [7:0]    maskDestinationResult_lo_lo_39 = {maskDestinationResult_lo_lo_hi_38, maskDestinationResult_lo_lo_lo_38};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_37 = {sourceDataVec_9[13], sourceDataVec_8[13]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_37 = {sourceDataVec_11[13], sourceDataVec_10[13]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_38 = {maskDestinationResult_lo_hi_lo_hi_37, maskDestinationResult_lo_hi_lo_lo_37};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_37 = {sourceDataVec_13[13], sourceDataVec_12[13]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_37 = {sourceDataVec_15[13], sourceDataVec_14[13]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_38 = {maskDestinationResult_lo_hi_hi_hi_37, maskDestinationResult_lo_hi_hi_lo_37};
  wire [7:0]    maskDestinationResult_lo_hi_39 = {maskDestinationResult_lo_hi_hi_38, maskDestinationResult_lo_hi_lo_38};
  wire [15:0]   maskDestinationResult_lo_295 = {maskDestinationResult_lo_hi_39, maskDestinationResult_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_37 = {sourceDataVec_17[13], sourceDataVec_16[13]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_37 = {sourceDataVec_19[13], sourceDataVec_18[13]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_38 = {maskDestinationResult_hi_lo_lo_hi_37, maskDestinationResult_hi_lo_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_37 = {sourceDataVec_21[13], sourceDataVec_20[13]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_37 = {sourceDataVec_23[13], sourceDataVec_22[13]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_38 = {maskDestinationResult_hi_lo_hi_hi_37, maskDestinationResult_hi_lo_hi_lo_37};
  wire [7:0]    maskDestinationResult_hi_lo_39 = {maskDestinationResult_hi_lo_hi_38, maskDestinationResult_hi_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_37 = {sourceDataVec_25[13], sourceDataVec_24[13]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_37 = {sourceDataVec_27[13], sourceDataVec_26[13]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_38 = {maskDestinationResult_hi_hi_lo_hi_37, maskDestinationResult_hi_hi_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_37 = {sourceDataVec_29[13], sourceDataVec_28[13]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_37 = {sourceDataVec_31[13], sourceDataVec_30[13]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_38 = {maskDestinationResult_hi_hi_hi_hi_37, maskDestinationResult_hi_hi_hi_lo_37};
  wire [7:0]    maskDestinationResult_hi_hi_39 = {maskDestinationResult_hi_hi_hi_38, maskDestinationResult_hi_hi_lo_38};
  wire [15:0]   maskDestinationResult_hi_295 = {maskDestinationResult_hi_hi_39, maskDestinationResult_hi_lo_39};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_38 = {sourceDataVec_1[14], sourceDataVec_0[14]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_38 = {sourceDataVec_3[14], sourceDataVec_2[14]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_39 = {maskDestinationResult_lo_lo_lo_hi_38, maskDestinationResult_lo_lo_lo_lo_38};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_38 = {sourceDataVec_5[14], sourceDataVec_4[14]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_38 = {sourceDataVec_7[14], sourceDataVec_6[14]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_39 = {maskDestinationResult_lo_lo_hi_hi_38, maskDestinationResult_lo_lo_hi_lo_38};
  wire [7:0]    maskDestinationResult_lo_lo_40 = {maskDestinationResult_lo_lo_hi_39, maskDestinationResult_lo_lo_lo_39};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_38 = {sourceDataVec_9[14], sourceDataVec_8[14]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_38 = {sourceDataVec_11[14], sourceDataVec_10[14]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_39 = {maskDestinationResult_lo_hi_lo_hi_38, maskDestinationResult_lo_hi_lo_lo_38};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_38 = {sourceDataVec_13[14], sourceDataVec_12[14]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_38 = {sourceDataVec_15[14], sourceDataVec_14[14]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_39 = {maskDestinationResult_lo_hi_hi_hi_38, maskDestinationResult_lo_hi_hi_lo_38};
  wire [7:0]    maskDestinationResult_lo_hi_40 = {maskDestinationResult_lo_hi_hi_39, maskDestinationResult_lo_hi_lo_39};
  wire [15:0]   maskDestinationResult_lo_296 = {maskDestinationResult_lo_hi_40, maskDestinationResult_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_38 = {sourceDataVec_17[14], sourceDataVec_16[14]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_38 = {sourceDataVec_19[14], sourceDataVec_18[14]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_39 = {maskDestinationResult_hi_lo_lo_hi_38, maskDestinationResult_hi_lo_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_38 = {sourceDataVec_21[14], sourceDataVec_20[14]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_38 = {sourceDataVec_23[14], sourceDataVec_22[14]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_39 = {maskDestinationResult_hi_lo_hi_hi_38, maskDestinationResult_hi_lo_hi_lo_38};
  wire [7:0]    maskDestinationResult_hi_lo_40 = {maskDestinationResult_hi_lo_hi_39, maskDestinationResult_hi_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_38 = {sourceDataVec_25[14], sourceDataVec_24[14]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_38 = {sourceDataVec_27[14], sourceDataVec_26[14]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_39 = {maskDestinationResult_hi_hi_lo_hi_38, maskDestinationResult_hi_hi_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_38 = {sourceDataVec_29[14], sourceDataVec_28[14]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_38 = {sourceDataVec_31[14], sourceDataVec_30[14]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_39 = {maskDestinationResult_hi_hi_hi_hi_38, maskDestinationResult_hi_hi_hi_lo_38};
  wire [7:0]    maskDestinationResult_hi_hi_40 = {maskDestinationResult_hi_hi_hi_39, maskDestinationResult_hi_hi_lo_39};
  wire [15:0]   maskDestinationResult_hi_296 = {maskDestinationResult_hi_hi_40, maskDestinationResult_hi_lo_40};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_39 = {sourceDataVec_1[15], sourceDataVec_0[15]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_39 = {sourceDataVec_3[15], sourceDataVec_2[15]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_40 = {maskDestinationResult_lo_lo_lo_hi_39, maskDestinationResult_lo_lo_lo_lo_39};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_39 = {sourceDataVec_5[15], sourceDataVec_4[15]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_39 = {sourceDataVec_7[15], sourceDataVec_6[15]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_40 = {maskDestinationResult_lo_lo_hi_hi_39, maskDestinationResult_lo_lo_hi_lo_39};
  wire [7:0]    maskDestinationResult_lo_lo_41 = {maskDestinationResult_lo_lo_hi_40, maskDestinationResult_lo_lo_lo_40};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_39 = {sourceDataVec_9[15], sourceDataVec_8[15]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_39 = {sourceDataVec_11[15], sourceDataVec_10[15]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_40 = {maskDestinationResult_lo_hi_lo_hi_39, maskDestinationResult_lo_hi_lo_lo_39};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_39 = {sourceDataVec_13[15], sourceDataVec_12[15]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_39 = {sourceDataVec_15[15], sourceDataVec_14[15]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_40 = {maskDestinationResult_lo_hi_hi_hi_39, maskDestinationResult_lo_hi_hi_lo_39};
  wire [7:0]    maskDestinationResult_lo_hi_41 = {maskDestinationResult_lo_hi_hi_40, maskDestinationResult_lo_hi_lo_40};
  wire [15:0]   maskDestinationResult_lo_297 = {maskDestinationResult_lo_hi_41, maskDestinationResult_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_39 = {sourceDataVec_17[15], sourceDataVec_16[15]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_39 = {sourceDataVec_19[15], sourceDataVec_18[15]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_40 = {maskDestinationResult_hi_lo_lo_hi_39, maskDestinationResult_hi_lo_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_39 = {sourceDataVec_21[15], sourceDataVec_20[15]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_39 = {sourceDataVec_23[15], sourceDataVec_22[15]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_40 = {maskDestinationResult_hi_lo_hi_hi_39, maskDestinationResult_hi_lo_hi_lo_39};
  wire [7:0]    maskDestinationResult_hi_lo_41 = {maskDestinationResult_hi_lo_hi_40, maskDestinationResult_hi_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_39 = {sourceDataVec_25[15], sourceDataVec_24[15]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_39 = {sourceDataVec_27[15], sourceDataVec_26[15]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_40 = {maskDestinationResult_hi_hi_lo_hi_39, maskDestinationResult_hi_hi_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_39 = {sourceDataVec_29[15], sourceDataVec_28[15]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_39 = {sourceDataVec_31[15], sourceDataVec_30[15]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_40 = {maskDestinationResult_hi_hi_hi_hi_39, maskDestinationResult_hi_hi_hi_lo_39};
  wire [7:0]    maskDestinationResult_hi_hi_41 = {maskDestinationResult_hi_hi_hi_40, maskDestinationResult_hi_hi_lo_40};
  wire [15:0]   maskDestinationResult_hi_297 = {maskDestinationResult_hi_hi_41, maskDestinationResult_hi_lo_41};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_40 = {sourceDataVec_1[16], sourceDataVec_0[16]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_40 = {sourceDataVec_3[16], sourceDataVec_2[16]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_41 = {maskDestinationResult_lo_lo_lo_hi_40, maskDestinationResult_lo_lo_lo_lo_40};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_40 = {sourceDataVec_5[16], sourceDataVec_4[16]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_40 = {sourceDataVec_7[16], sourceDataVec_6[16]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_41 = {maskDestinationResult_lo_lo_hi_hi_40, maskDestinationResult_lo_lo_hi_lo_40};
  wire [7:0]    maskDestinationResult_lo_lo_42 = {maskDestinationResult_lo_lo_hi_41, maskDestinationResult_lo_lo_lo_41};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_40 = {sourceDataVec_9[16], sourceDataVec_8[16]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_40 = {sourceDataVec_11[16], sourceDataVec_10[16]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_41 = {maskDestinationResult_lo_hi_lo_hi_40, maskDestinationResult_lo_hi_lo_lo_40};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_40 = {sourceDataVec_13[16], sourceDataVec_12[16]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_40 = {sourceDataVec_15[16], sourceDataVec_14[16]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_41 = {maskDestinationResult_lo_hi_hi_hi_40, maskDestinationResult_lo_hi_hi_lo_40};
  wire [7:0]    maskDestinationResult_lo_hi_42 = {maskDestinationResult_lo_hi_hi_41, maskDestinationResult_lo_hi_lo_41};
  wire [15:0]   maskDestinationResult_lo_298 = {maskDestinationResult_lo_hi_42, maskDestinationResult_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_40 = {sourceDataVec_17[16], sourceDataVec_16[16]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_40 = {sourceDataVec_19[16], sourceDataVec_18[16]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_41 = {maskDestinationResult_hi_lo_lo_hi_40, maskDestinationResult_hi_lo_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_40 = {sourceDataVec_21[16], sourceDataVec_20[16]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_40 = {sourceDataVec_23[16], sourceDataVec_22[16]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_41 = {maskDestinationResult_hi_lo_hi_hi_40, maskDestinationResult_hi_lo_hi_lo_40};
  wire [7:0]    maskDestinationResult_hi_lo_42 = {maskDestinationResult_hi_lo_hi_41, maskDestinationResult_hi_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_40 = {sourceDataVec_25[16], sourceDataVec_24[16]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_40 = {sourceDataVec_27[16], sourceDataVec_26[16]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_41 = {maskDestinationResult_hi_hi_lo_hi_40, maskDestinationResult_hi_hi_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_40 = {sourceDataVec_29[16], sourceDataVec_28[16]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_40 = {sourceDataVec_31[16], sourceDataVec_30[16]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_41 = {maskDestinationResult_hi_hi_hi_hi_40, maskDestinationResult_hi_hi_hi_lo_40};
  wire [7:0]    maskDestinationResult_hi_hi_42 = {maskDestinationResult_hi_hi_hi_41, maskDestinationResult_hi_hi_lo_41};
  wire [15:0]   maskDestinationResult_hi_298 = {maskDestinationResult_hi_hi_42, maskDestinationResult_hi_lo_42};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_41 = {sourceDataVec_1[17], sourceDataVec_0[17]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_41 = {sourceDataVec_3[17], sourceDataVec_2[17]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_42 = {maskDestinationResult_lo_lo_lo_hi_41, maskDestinationResult_lo_lo_lo_lo_41};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_41 = {sourceDataVec_5[17], sourceDataVec_4[17]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_41 = {sourceDataVec_7[17], sourceDataVec_6[17]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_42 = {maskDestinationResult_lo_lo_hi_hi_41, maskDestinationResult_lo_lo_hi_lo_41};
  wire [7:0]    maskDestinationResult_lo_lo_43 = {maskDestinationResult_lo_lo_hi_42, maskDestinationResult_lo_lo_lo_42};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_41 = {sourceDataVec_9[17], sourceDataVec_8[17]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_41 = {sourceDataVec_11[17], sourceDataVec_10[17]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_42 = {maskDestinationResult_lo_hi_lo_hi_41, maskDestinationResult_lo_hi_lo_lo_41};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_41 = {sourceDataVec_13[17], sourceDataVec_12[17]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_41 = {sourceDataVec_15[17], sourceDataVec_14[17]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_42 = {maskDestinationResult_lo_hi_hi_hi_41, maskDestinationResult_lo_hi_hi_lo_41};
  wire [7:0]    maskDestinationResult_lo_hi_43 = {maskDestinationResult_lo_hi_hi_42, maskDestinationResult_lo_hi_lo_42};
  wire [15:0]   maskDestinationResult_lo_299 = {maskDestinationResult_lo_hi_43, maskDestinationResult_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_41 = {sourceDataVec_17[17], sourceDataVec_16[17]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_41 = {sourceDataVec_19[17], sourceDataVec_18[17]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_42 = {maskDestinationResult_hi_lo_lo_hi_41, maskDestinationResult_hi_lo_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_41 = {sourceDataVec_21[17], sourceDataVec_20[17]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_41 = {sourceDataVec_23[17], sourceDataVec_22[17]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_42 = {maskDestinationResult_hi_lo_hi_hi_41, maskDestinationResult_hi_lo_hi_lo_41};
  wire [7:0]    maskDestinationResult_hi_lo_43 = {maskDestinationResult_hi_lo_hi_42, maskDestinationResult_hi_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_41 = {sourceDataVec_25[17], sourceDataVec_24[17]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_41 = {sourceDataVec_27[17], sourceDataVec_26[17]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_42 = {maskDestinationResult_hi_hi_lo_hi_41, maskDestinationResult_hi_hi_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_41 = {sourceDataVec_29[17], sourceDataVec_28[17]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_41 = {sourceDataVec_31[17], sourceDataVec_30[17]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_42 = {maskDestinationResult_hi_hi_hi_hi_41, maskDestinationResult_hi_hi_hi_lo_41};
  wire [7:0]    maskDestinationResult_hi_hi_43 = {maskDestinationResult_hi_hi_hi_42, maskDestinationResult_hi_hi_lo_42};
  wire [15:0]   maskDestinationResult_hi_299 = {maskDestinationResult_hi_hi_43, maskDestinationResult_hi_lo_43};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_42 = {sourceDataVec_1[18], sourceDataVec_0[18]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_42 = {sourceDataVec_3[18], sourceDataVec_2[18]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_43 = {maskDestinationResult_lo_lo_lo_hi_42, maskDestinationResult_lo_lo_lo_lo_42};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_42 = {sourceDataVec_5[18], sourceDataVec_4[18]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_42 = {sourceDataVec_7[18], sourceDataVec_6[18]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_43 = {maskDestinationResult_lo_lo_hi_hi_42, maskDestinationResult_lo_lo_hi_lo_42};
  wire [7:0]    maskDestinationResult_lo_lo_44 = {maskDestinationResult_lo_lo_hi_43, maskDestinationResult_lo_lo_lo_43};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_42 = {sourceDataVec_9[18], sourceDataVec_8[18]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_42 = {sourceDataVec_11[18], sourceDataVec_10[18]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_43 = {maskDestinationResult_lo_hi_lo_hi_42, maskDestinationResult_lo_hi_lo_lo_42};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_42 = {sourceDataVec_13[18], sourceDataVec_12[18]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_42 = {sourceDataVec_15[18], sourceDataVec_14[18]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_43 = {maskDestinationResult_lo_hi_hi_hi_42, maskDestinationResult_lo_hi_hi_lo_42};
  wire [7:0]    maskDestinationResult_lo_hi_44 = {maskDestinationResult_lo_hi_hi_43, maskDestinationResult_lo_hi_lo_43};
  wire [15:0]   maskDestinationResult_lo_300 = {maskDestinationResult_lo_hi_44, maskDestinationResult_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_42 = {sourceDataVec_17[18], sourceDataVec_16[18]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_42 = {sourceDataVec_19[18], sourceDataVec_18[18]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_43 = {maskDestinationResult_hi_lo_lo_hi_42, maskDestinationResult_hi_lo_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_42 = {sourceDataVec_21[18], sourceDataVec_20[18]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_42 = {sourceDataVec_23[18], sourceDataVec_22[18]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_43 = {maskDestinationResult_hi_lo_hi_hi_42, maskDestinationResult_hi_lo_hi_lo_42};
  wire [7:0]    maskDestinationResult_hi_lo_44 = {maskDestinationResult_hi_lo_hi_43, maskDestinationResult_hi_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_42 = {sourceDataVec_25[18], sourceDataVec_24[18]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_42 = {sourceDataVec_27[18], sourceDataVec_26[18]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_43 = {maskDestinationResult_hi_hi_lo_hi_42, maskDestinationResult_hi_hi_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_42 = {sourceDataVec_29[18], sourceDataVec_28[18]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_42 = {sourceDataVec_31[18], sourceDataVec_30[18]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_43 = {maskDestinationResult_hi_hi_hi_hi_42, maskDestinationResult_hi_hi_hi_lo_42};
  wire [7:0]    maskDestinationResult_hi_hi_44 = {maskDestinationResult_hi_hi_hi_43, maskDestinationResult_hi_hi_lo_43};
  wire [15:0]   maskDestinationResult_hi_300 = {maskDestinationResult_hi_hi_44, maskDestinationResult_hi_lo_44};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_43 = {sourceDataVec_1[19], sourceDataVec_0[19]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_43 = {sourceDataVec_3[19], sourceDataVec_2[19]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_44 = {maskDestinationResult_lo_lo_lo_hi_43, maskDestinationResult_lo_lo_lo_lo_43};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_43 = {sourceDataVec_5[19], sourceDataVec_4[19]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_43 = {sourceDataVec_7[19], sourceDataVec_6[19]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_44 = {maskDestinationResult_lo_lo_hi_hi_43, maskDestinationResult_lo_lo_hi_lo_43};
  wire [7:0]    maskDestinationResult_lo_lo_45 = {maskDestinationResult_lo_lo_hi_44, maskDestinationResult_lo_lo_lo_44};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_43 = {sourceDataVec_9[19], sourceDataVec_8[19]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_43 = {sourceDataVec_11[19], sourceDataVec_10[19]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_44 = {maskDestinationResult_lo_hi_lo_hi_43, maskDestinationResult_lo_hi_lo_lo_43};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_43 = {sourceDataVec_13[19], sourceDataVec_12[19]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_43 = {sourceDataVec_15[19], sourceDataVec_14[19]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_44 = {maskDestinationResult_lo_hi_hi_hi_43, maskDestinationResult_lo_hi_hi_lo_43};
  wire [7:0]    maskDestinationResult_lo_hi_45 = {maskDestinationResult_lo_hi_hi_44, maskDestinationResult_lo_hi_lo_44};
  wire [15:0]   maskDestinationResult_lo_301 = {maskDestinationResult_lo_hi_45, maskDestinationResult_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_43 = {sourceDataVec_17[19], sourceDataVec_16[19]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_43 = {sourceDataVec_19[19], sourceDataVec_18[19]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_44 = {maskDestinationResult_hi_lo_lo_hi_43, maskDestinationResult_hi_lo_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_43 = {sourceDataVec_21[19], sourceDataVec_20[19]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_43 = {sourceDataVec_23[19], sourceDataVec_22[19]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_44 = {maskDestinationResult_hi_lo_hi_hi_43, maskDestinationResult_hi_lo_hi_lo_43};
  wire [7:0]    maskDestinationResult_hi_lo_45 = {maskDestinationResult_hi_lo_hi_44, maskDestinationResult_hi_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_43 = {sourceDataVec_25[19], sourceDataVec_24[19]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_43 = {sourceDataVec_27[19], sourceDataVec_26[19]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_44 = {maskDestinationResult_hi_hi_lo_hi_43, maskDestinationResult_hi_hi_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_43 = {sourceDataVec_29[19], sourceDataVec_28[19]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_43 = {sourceDataVec_31[19], sourceDataVec_30[19]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_44 = {maskDestinationResult_hi_hi_hi_hi_43, maskDestinationResult_hi_hi_hi_lo_43};
  wire [7:0]    maskDestinationResult_hi_hi_45 = {maskDestinationResult_hi_hi_hi_44, maskDestinationResult_hi_hi_lo_44};
  wire [15:0]   maskDestinationResult_hi_301 = {maskDestinationResult_hi_hi_45, maskDestinationResult_hi_lo_45};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_44 = {sourceDataVec_1[20], sourceDataVec_0[20]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_44 = {sourceDataVec_3[20], sourceDataVec_2[20]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_45 = {maskDestinationResult_lo_lo_lo_hi_44, maskDestinationResult_lo_lo_lo_lo_44};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_44 = {sourceDataVec_5[20], sourceDataVec_4[20]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_44 = {sourceDataVec_7[20], sourceDataVec_6[20]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_45 = {maskDestinationResult_lo_lo_hi_hi_44, maskDestinationResult_lo_lo_hi_lo_44};
  wire [7:0]    maskDestinationResult_lo_lo_46 = {maskDestinationResult_lo_lo_hi_45, maskDestinationResult_lo_lo_lo_45};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_44 = {sourceDataVec_9[20], sourceDataVec_8[20]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_44 = {sourceDataVec_11[20], sourceDataVec_10[20]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_45 = {maskDestinationResult_lo_hi_lo_hi_44, maskDestinationResult_lo_hi_lo_lo_44};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_44 = {sourceDataVec_13[20], sourceDataVec_12[20]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_44 = {sourceDataVec_15[20], sourceDataVec_14[20]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_45 = {maskDestinationResult_lo_hi_hi_hi_44, maskDestinationResult_lo_hi_hi_lo_44};
  wire [7:0]    maskDestinationResult_lo_hi_46 = {maskDestinationResult_lo_hi_hi_45, maskDestinationResult_lo_hi_lo_45};
  wire [15:0]   maskDestinationResult_lo_302 = {maskDestinationResult_lo_hi_46, maskDestinationResult_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_44 = {sourceDataVec_17[20], sourceDataVec_16[20]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_44 = {sourceDataVec_19[20], sourceDataVec_18[20]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_45 = {maskDestinationResult_hi_lo_lo_hi_44, maskDestinationResult_hi_lo_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_44 = {sourceDataVec_21[20], sourceDataVec_20[20]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_44 = {sourceDataVec_23[20], sourceDataVec_22[20]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_45 = {maskDestinationResult_hi_lo_hi_hi_44, maskDestinationResult_hi_lo_hi_lo_44};
  wire [7:0]    maskDestinationResult_hi_lo_46 = {maskDestinationResult_hi_lo_hi_45, maskDestinationResult_hi_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_44 = {sourceDataVec_25[20], sourceDataVec_24[20]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_44 = {sourceDataVec_27[20], sourceDataVec_26[20]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_45 = {maskDestinationResult_hi_hi_lo_hi_44, maskDestinationResult_hi_hi_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_44 = {sourceDataVec_29[20], sourceDataVec_28[20]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_44 = {sourceDataVec_31[20], sourceDataVec_30[20]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_45 = {maskDestinationResult_hi_hi_hi_hi_44, maskDestinationResult_hi_hi_hi_lo_44};
  wire [7:0]    maskDestinationResult_hi_hi_46 = {maskDestinationResult_hi_hi_hi_45, maskDestinationResult_hi_hi_lo_45};
  wire [15:0]   maskDestinationResult_hi_302 = {maskDestinationResult_hi_hi_46, maskDestinationResult_hi_lo_46};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_45 = {sourceDataVec_1[21], sourceDataVec_0[21]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_45 = {sourceDataVec_3[21], sourceDataVec_2[21]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_46 = {maskDestinationResult_lo_lo_lo_hi_45, maskDestinationResult_lo_lo_lo_lo_45};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_45 = {sourceDataVec_5[21], sourceDataVec_4[21]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_45 = {sourceDataVec_7[21], sourceDataVec_6[21]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_46 = {maskDestinationResult_lo_lo_hi_hi_45, maskDestinationResult_lo_lo_hi_lo_45};
  wire [7:0]    maskDestinationResult_lo_lo_47 = {maskDestinationResult_lo_lo_hi_46, maskDestinationResult_lo_lo_lo_46};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_45 = {sourceDataVec_9[21], sourceDataVec_8[21]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_45 = {sourceDataVec_11[21], sourceDataVec_10[21]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_46 = {maskDestinationResult_lo_hi_lo_hi_45, maskDestinationResult_lo_hi_lo_lo_45};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_45 = {sourceDataVec_13[21], sourceDataVec_12[21]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_45 = {sourceDataVec_15[21], sourceDataVec_14[21]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_46 = {maskDestinationResult_lo_hi_hi_hi_45, maskDestinationResult_lo_hi_hi_lo_45};
  wire [7:0]    maskDestinationResult_lo_hi_47 = {maskDestinationResult_lo_hi_hi_46, maskDestinationResult_lo_hi_lo_46};
  wire [15:0]   maskDestinationResult_lo_303 = {maskDestinationResult_lo_hi_47, maskDestinationResult_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_45 = {sourceDataVec_17[21], sourceDataVec_16[21]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_45 = {sourceDataVec_19[21], sourceDataVec_18[21]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_46 = {maskDestinationResult_hi_lo_lo_hi_45, maskDestinationResult_hi_lo_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_45 = {sourceDataVec_21[21], sourceDataVec_20[21]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_45 = {sourceDataVec_23[21], sourceDataVec_22[21]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_46 = {maskDestinationResult_hi_lo_hi_hi_45, maskDestinationResult_hi_lo_hi_lo_45};
  wire [7:0]    maskDestinationResult_hi_lo_47 = {maskDestinationResult_hi_lo_hi_46, maskDestinationResult_hi_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_45 = {sourceDataVec_25[21], sourceDataVec_24[21]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_45 = {sourceDataVec_27[21], sourceDataVec_26[21]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_46 = {maskDestinationResult_hi_hi_lo_hi_45, maskDestinationResult_hi_hi_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_45 = {sourceDataVec_29[21], sourceDataVec_28[21]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_45 = {sourceDataVec_31[21], sourceDataVec_30[21]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_46 = {maskDestinationResult_hi_hi_hi_hi_45, maskDestinationResult_hi_hi_hi_lo_45};
  wire [7:0]    maskDestinationResult_hi_hi_47 = {maskDestinationResult_hi_hi_hi_46, maskDestinationResult_hi_hi_lo_46};
  wire [15:0]   maskDestinationResult_hi_303 = {maskDestinationResult_hi_hi_47, maskDestinationResult_hi_lo_47};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_46 = {sourceDataVec_1[22], sourceDataVec_0[22]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_46 = {sourceDataVec_3[22], sourceDataVec_2[22]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_47 = {maskDestinationResult_lo_lo_lo_hi_46, maskDestinationResult_lo_lo_lo_lo_46};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_46 = {sourceDataVec_5[22], sourceDataVec_4[22]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_46 = {sourceDataVec_7[22], sourceDataVec_6[22]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_47 = {maskDestinationResult_lo_lo_hi_hi_46, maskDestinationResult_lo_lo_hi_lo_46};
  wire [7:0]    maskDestinationResult_lo_lo_48 = {maskDestinationResult_lo_lo_hi_47, maskDestinationResult_lo_lo_lo_47};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_46 = {sourceDataVec_9[22], sourceDataVec_8[22]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_46 = {sourceDataVec_11[22], sourceDataVec_10[22]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_47 = {maskDestinationResult_lo_hi_lo_hi_46, maskDestinationResult_lo_hi_lo_lo_46};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_46 = {sourceDataVec_13[22], sourceDataVec_12[22]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_46 = {sourceDataVec_15[22], sourceDataVec_14[22]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_47 = {maskDestinationResult_lo_hi_hi_hi_46, maskDestinationResult_lo_hi_hi_lo_46};
  wire [7:0]    maskDestinationResult_lo_hi_48 = {maskDestinationResult_lo_hi_hi_47, maskDestinationResult_lo_hi_lo_47};
  wire [15:0]   maskDestinationResult_lo_304 = {maskDestinationResult_lo_hi_48, maskDestinationResult_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_46 = {sourceDataVec_17[22], sourceDataVec_16[22]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_46 = {sourceDataVec_19[22], sourceDataVec_18[22]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_47 = {maskDestinationResult_hi_lo_lo_hi_46, maskDestinationResult_hi_lo_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_46 = {sourceDataVec_21[22], sourceDataVec_20[22]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_46 = {sourceDataVec_23[22], sourceDataVec_22[22]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_47 = {maskDestinationResult_hi_lo_hi_hi_46, maskDestinationResult_hi_lo_hi_lo_46};
  wire [7:0]    maskDestinationResult_hi_lo_48 = {maskDestinationResult_hi_lo_hi_47, maskDestinationResult_hi_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_46 = {sourceDataVec_25[22], sourceDataVec_24[22]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_46 = {sourceDataVec_27[22], sourceDataVec_26[22]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_47 = {maskDestinationResult_hi_hi_lo_hi_46, maskDestinationResult_hi_hi_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_46 = {sourceDataVec_29[22], sourceDataVec_28[22]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_46 = {sourceDataVec_31[22], sourceDataVec_30[22]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_47 = {maskDestinationResult_hi_hi_hi_hi_46, maskDestinationResult_hi_hi_hi_lo_46};
  wire [7:0]    maskDestinationResult_hi_hi_48 = {maskDestinationResult_hi_hi_hi_47, maskDestinationResult_hi_hi_lo_47};
  wire [15:0]   maskDestinationResult_hi_304 = {maskDestinationResult_hi_hi_48, maskDestinationResult_hi_lo_48};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_47 = {sourceDataVec_1[23], sourceDataVec_0[23]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_47 = {sourceDataVec_3[23], sourceDataVec_2[23]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_48 = {maskDestinationResult_lo_lo_lo_hi_47, maskDestinationResult_lo_lo_lo_lo_47};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_47 = {sourceDataVec_5[23], sourceDataVec_4[23]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_47 = {sourceDataVec_7[23], sourceDataVec_6[23]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_48 = {maskDestinationResult_lo_lo_hi_hi_47, maskDestinationResult_lo_lo_hi_lo_47};
  wire [7:0]    maskDestinationResult_lo_lo_49 = {maskDestinationResult_lo_lo_hi_48, maskDestinationResult_lo_lo_lo_48};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_47 = {sourceDataVec_9[23], sourceDataVec_8[23]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_47 = {sourceDataVec_11[23], sourceDataVec_10[23]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_48 = {maskDestinationResult_lo_hi_lo_hi_47, maskDestinationResult_lo_hi_lo_lo_47};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_47 = {sourceDataVec_13[23], sourceDataVec_12[23]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_47 = {sourceDataVec_15[23], sourceDataVec_14[23]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_48 = {maskDestinationResult_lo_hi_hi_hi_47, maskDestinationResult_lo_hi_hi_lo_47};
  wire [7:0]    maskDestinationResult_lo_hi_49 = {maskDestinationResult_lo_hi_hi_48, maskDestinationResult_lo_hi_lo_48};
  wire [15:0]   maskDestinationResult_lo_305 = {maskDestinationResult_lo_hi_49, maskDestinationResult_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_47 = {sourceDataVec_17[23], sourceDataVec_16[23]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_47 = {sourceDataVec_19[23], sourceDataVec_18[23]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_48 = {maskDestinationResult_hi_lo_lo_hi_47, maskDestinationResult_hi_lo_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_47 = {sourceDataVec_21[23], sourceDataVec_20[23]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_47 = {sourceDataVec_23[23], sourceDataVec_22[23]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_48 = {maskDestinationResult_hi_lo_hi_hi_47, maskDestinationResult_hi_lo_hi_lo_47};
  wire [7:0]    maskDestinationResult_hi_lo_49 = {maskDestinationResult_hi_lo_hi_48, maskDestinationResult_hi_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_47 = {sourceDataVec_25[23], sourceDataVec_24[23]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_47 = {sourceDataVec_27[23], sourceDataVec_26[23]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_48 = {maskDestinationResult_hi_hi_lo_hi_47, maskDestinationResult_hi_hi_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_47 = {sourceDataVec_29[23], sourceDataVec_28[23]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_47 = {sourceDataVec_31[23], sourceDataVec_30[23]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_48 = {maskDestinationResult_hi_hi_hi_hi_47, maskDestinationResult_hi_hi_hi_lo_47};
  wire [7:0]    maskDestinationResult_hi_hi_49 = {maskDestinationResult_hi_hi_hi_48, maskDestinationResult_hi_hi_lo_48};
  wire [15:0]   maskDestinationResult_hi_305 = {maskDestinationResult_hi_hi_49, maskDestinationResult_hi_lo_49};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_48 = {sourceDataVec_1[24], sourceDataVec_0[24]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_48 = {sourceDataVec_3[24], sourceDataVec_2[24]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_49 = {maskDestinationResult_lo_lo_lo_hi_48, maskDestinationResult_lo_lo_lo_lo_48};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_48 = {sourceDataVec_5[24], sourceDataVec_4[24]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_48 = {sourceDataVec_7[24], sourceDataVec_6[24]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_49 = {maskDestinationResult_lo_lo_hi_hi_48, maskDestinationResult_lo_lo_hi_lo_48};
  wire [7:0]    maskDestinationResult_lo_lo_50 = {maskDestinationResult_lo_lo_hi_49, maskDestinationResult_lo_lo_lo_49};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_48 = {sourceDataVec_9[24], sourceDataVec_8[24]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_48 = {sourceDataVec_11[24], sourceDataVec_10[24]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_49 = {maskDestinationResult_lo_hi_lo_hi_48, maskDestinationResult_lo_hi_lo_lo_48};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_48 = {sourceDataVec_13[24], sourceDataVec_12[24]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_48 = {sourceDataVec_15[24], sourceDataVec_14[24]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_49 = {maskDestinationResult_lo_hi_hi_hi_48, maskDestinationResult_lo_hi_hi_lo_48};
  wire [7:0]    maskDestinationResult_lo_hi_50 = {maskDestinationResult_lo_hi_hi_49, maskDestinationResult_lo_hi_lo_49};
  wire [15:0]   maskDestinationResult_lo_306 = {maskDestinationResult_lo_hi_50, maskDestinationResult_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_48 = {sourceDataVec_17[24], sourceDataVec_16[24]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_48 = {sourceDataVec_19[24], sourceDataVec_18[24]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_49 = {maskDestinationResult_hi_lo_lo_hi_48, maskDestinationResult_hi_lo_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_48 = {sourceDataVec_21[24], sourceDataVec_20[24]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_48 = {sourceDataVec_23[24], sourceDataVec_22[24]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_49 = {maskDestinationResult_hi_lo_hi_hi_48, maskDestinationResult_hi_lo_hi_lo_48};
  wire [7:0]    maskDestinationResult_hi_lo_50 = {maskDestinationResult_hi_lo_hi_49, maskDestinationResult_hi_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_48 = {sourceDataVec_25[24], sourceDataVec_24[24]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_48 = {sourceDataVec_27[24], sourceDataVec_26[24]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_49 = {maskDestinationResult_hi_hi_lo_hi_48, maskDestinationResult_hi_hi_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_48 = {sourceDataVec_29[24], sourceDataVec_28[24]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_48 = {sourceDataVec_31[24], sourceDataVec_30[24]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_49 = {maskDestinationResult_hi_hi_hi_hi_48, maskDestinationResult_hi_hi_hi_lo_48};
  wire [7:0]    maskDestinationResult_hi_hi_50 = {maskDestinationResult_hi_hi_hi_49, maskDestinationResult_hi_hi_lo_49};
  wire [15:0]   maskDestinationResult_hi_306 = {maskDestinationResult_hi_hi_50, maskDestinationResult_hi_lo_50};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_49 = {sourceDataVec_1[25], sourceDataVec_0[25]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_49 = {sourceDataVec_3[25], sourceDataVec_2[25]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_50 = {maskDestinationResult_lo_lo_lo_hi_49, maskDestinationResult_lo_lo_lo_lo_49};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_49 = {sourceDataVec_5[25], sourceDataVec_4[25]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_49 = {sourceDataVec_7[25], sourceDataVec_6[25]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_50 = {maskDestinationResult_lo_lo_hi_hi_49, maskDestinationResult_lo_lo_hi_lo_49};
  wire [7:0]    maskDestinationResult_lo_lo_51 = {maskDestinationResult_lo_lo_hi_50, maskDestinationResult_lo_lo_lo_50};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_49 = {sourceDataVec_9[25], sourceDataVec_8[25]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_49 = {sourceDataVec_11[25], sourceDataVec_10[25]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_50 = {maskDestinationResult_lo_hi_lo_hi_49, maskDestinationResult_lo_hi_lo_lo_49};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_49 = {sourceDataVec_13[25], sourceDataVec_12[25]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_49 = {sourceDataVec_15[25], sourceDataVec_14[25]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_50 = {maskDestinationResult_lo_hi_hi_hi_49, maskDestinationResult_lo_hi_hi_lo_49};
  wire [7:0]    maskDestinationResult_lo_hi_51 = {maskDestinationResult_lo_hi_hi_50, maskDestinationResult_lo_hi_lo_50};
  wire [15:0]   maskDestinationResult_lo_307 = {maskDestinationResult_lo_hi_51, maskDestinationResult_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_49 = {sourceDataVec_17[25], sourceDataVec_16[25]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_49 = {sourceDataVec_19[25], sourceDataVec_18[25]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_50 = {maskDestinationResult_hi_lo_lo_hi_49, maskDestinationResult_hi_lo_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_49 = {sourceDataVec_21[25], sourceDataVec_20[25]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_49 = {sourceDataVec_23[25], sourceDataVec_22[25]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_50 = {maskDestinationResult_hi_lo_hi_hi_49, maskDestinationResult_hi_lo_hi_lo_49};
  wire [7:0]    maskDestinationResult_hi_lo_51 = {maskDestinationResult_hi_lo_hi_50, maskDestinationResult_hi_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_49 = {sourceDataVec_25[25], sourceDataVec_24[25]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_49 = {sourceDataVec_27[25], sourceDataVec_26[25]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_50 = {maskDestinationResult_hi_hi_lo_hi_49, maskDestinationResult_hi_hi_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_49 = {sourceDataVec_29[25], sourceDataVec_28[25]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_49 = {sourceDataVec_31[25], sourceDataVec_30[25]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_50 = {maskDestinationResult_hi_hi_hi_hi_49, maskDestinationResult_hi_hi_hi_lo_49};
  wire [7:0]    maskDestinationResult_hi_hi_51 = {maskDestinationResult_hi_hi_hi_50, maskDestinationResult_hi_hi_lo_50};
  wire [15:0]   maskDestinationResult_hi_307 = {maskDestinationResult_hi_hi_51, maskDestinationResult_hi_lo_51};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_50 = {sourceDataVec_1[26], sourceDataVec_0[26]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_50 = {sourceDataVec_3[26], sourceDataVec_2[26]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_51 = {maskDestinationResult_lo_lo_lo_hi_50, maskDestinationResult_lo_lo_lo_lo_50};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_50 = {sourceDataVec_5[26], sourceDataVec_4[26]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_50 = {sourceDataVec_7[26], sourceDataVec_6[26]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_51 = {maskDestinationResult_lo_lo_hi_hi_50, maskDestinationResult_lo_lo_hi_lo_50};
  wire [7:0]    maskDestinationResult_lo_lo_52 = {maskDestinationResult_lo_lo_hi_51, maskDestinationResult_lo_lo_lo_51};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_50 = {sourceDataVec_9[26], sourceDataVec_8[26]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_50 = {sourceDataVec_11[26], sourceDataVec_10[26]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_51 = {maskDestinationResult_lo_hi_lo_hi_50, maskDestinationResult_lo_hi_lo_lo_50};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_50 = {sourceDataVec_13[26], sourceDataVec_12[26]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_50 = {sourceDataVec_15[26], sourceDataVec_14[26]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_51 = {maskDestinationResult_lo_hi_hi_hi_50, maskDestinationResult_lo_hi_hi_lo_50};
  wire [7:0]    maskDestinationResult_lo_hi_52 = {maskDestinationResult_lo_hi_hi_51, maskDestinationResult_lo_hi_lo_51};
  wire [15:0]   maskDestinationResult_lo_308 = {maskDestinationResult_lo_hi_52, maskDestinationResult_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_50 = {sourceDataVec_17[26], sourceDataVec_16[26]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_50 = {sourceDataVec_19[26], sourceDataVec_18[26]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_51 = {maskDestinationResult_hi_lo_lo_hi_50, maskDestinationResult_hi_lo_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_50 = {sourceDataVec_21[26], sourceDataVec_20[26]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_50 = {sourceDataVec_23[26], sourceDataVec_22[26]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_51 = {maskDestinationResult_hi_lo_hi_hi_50, maskDestinationResult_hi_lo_hi_lo_50};
  wire [7:0]    maskDestinationResult_hi_lo_52 = {maskDestinationResult_hi_lo_hi_51, maskDestinationResult_hi_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_50 = {sourceDataVec_25[26], sourceDataVec_24[26]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_50 = {sourceDataVec_27[26], sourceDataVec_26[26]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_51 = {maskDestinationResult_hi_hi_lo_hi_50, maskDestinationResult_hi_hi_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_50 = {sourceDataVec_29[26], sourceDataVec_28[26]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_50 = {sourceDataVec_31[26], sourceDataVec_30[26]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_51 = {maskDestinationResult_hi_hi_hi_hi_50, maskDestinationResult_hi_hi_hi_lo_50};
  wire [7:0]    maskDestinationResult_hi_hi_52 = {maskDestinationResult_hi_hi_hi_51, maskDestinationResult_hi_hi_lo_51};
  wire [15:0]   maskDestinationResult_hi_308 = {maskDestinationResult_hi_hi_52, maskDestinationResult_hi_lo_52};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_51 = {sourceDataVec_1[27], sourceDataVec_0[27]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_51 = {sourceDataVec_3[27], sourceDataVec_2[27]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_52 = {maskDestinationResult_lo_lo_lo_hi_51, maskDestinationResult_lo_lo_lo_lo_51};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_51 = {sourceDataVec_5[27], sourceDataVec_4[27]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_51 = {sourceDataVec_7[27], sourceDataVec_6[27]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_52 = {maskDestinationResult_lo_lo_hi_hi_51, maskDestinationResult_lo_lo_hi_lo_51};
  wire [7:0]    maskDestinationResult_lo_lo_53 = {maskDestinationResult_lo_lo_hi_52, maskDestinationResult_lo_lo_lo_52};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_51 = {sourceDataVec_9[27], sourceDataVec_8[27]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_51 = {sourceDataVec_11[27], sourceDataVec_10[27]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_52 = {maskDestinationResult_lo_hi_lo_hi_51, maskDestinationResult_lo_hi_lo_lo_51};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_51 = {sourceDataVec_13[27], sourceDataVec_12[27]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_51 = {sourceDataVec_15[27], sourceDataVec_14[27]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_52 = {maskDestinationResult_lo_hi_hi_hi_51, maskDestinationResult_lo_hi_hi_lo_51};
  wire [7:0]    maskDestinationResult_lo_hi_53 = {maskDestinationResult_lo_hi_hi_52, maskDestinationResult_lo_hi_lo_52};
  wire [15:0]   maskDestinationResult_lo_309 = {maskDestinationResult_lo_hi_53, maskDestinationResult_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_51 = {sourceDataVec_17[27], sourceDataVec_16[27]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_51 = {sourceDataVec_19[27], sourceDataVec_18[27]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_52 = {maskDestinationResult_hi_lo_lo_hi_51, maskDestinationResult_hi_lo_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_51 = {sourceDataVec_21[27], sourceDataVec_20[27]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_51 = {sourceDataVec_23[27], sourceDataVec_22[27]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_52 = {maskDestinationResult_hi_lo_hi_hi_51, maskDestinationResult_hi_lo_hi_lo_51};
  wire [7:0]    maskDestinationResult_hi_lo_53 = {maskDestinationResult_hi_lo_hi_52, maskDestinationResult_hi_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_51 = {sourceDataVec_25[27], sourceDataVec_24[27]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_51 = {sourceDataVec_27[27], sourceDataVec_26[27]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_52 = {maskDestinationResult_hi_hi_lo_hi_51, maskDestinationResult_hi_hi_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_51 = {sourceDataVec_29[27], sourceDataVec_28[27]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_51 = {sourceDataVec_31[27], sourceDataVec_30[27]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_52 = {maskDestinationResult_hi_hi_hi_hi_51, maskDestinationResult_hi_hi_hi_lo_51};
  wire [7:0]    maskDestinationResult_hi_hi_53 = {maskDestinationResult_hi_hi_hi_52, maskDestinationResult_hi_hi_lo_52};
  wire [15:0]   maskDestinationResult_hi_309 = {maskDestinationResult_hi_hi_53, maskDestinationResult_hi_lo_53};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_52 = {sourceDataVec_1[28], sourceDataVec_0[28]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_52 = {sourceDataVec_3[28], sourceDataVec_2[28]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_53 = {maskDestinationResult_lo_lo_lo_hi_52, maskDestinationResult_lo_lo_lo_lo_52};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_52 = {sourceDataVec_5[28], sourceDataVec_4[28]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_52 = {sourceDataVec_7[28], sourceDataVec_6[28]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_53 = {maskDestinationResult_lo_lo_hi_hi_52, maskDestinationResult_lo_lo_hi_lo_52};
  wire [7:0]    maskDestinationResult_lo_lo_54 = {maskDestinationResult_lo_lo_hi_53, maskDestinationResult_lo_lo_lo_53};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_52 = {sourceDataVec_9[28], sourceDataVec_8[28]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_52 = {sourceDataVec_11[28], sourceDataVec_10[28]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_53 = {maskDestinationResult_lo_hi_lo_hi_52, maskDestinationResult_lo_hi_lo_lo_52};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_52 = {sourceDataVec_13[28], sourceDataVec_12[28]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_52 = {sourceDataVec_15[28], sourceDataVec_14[28]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_53 = {maskDestinationResult_lo_hi_hi_hi_52, maskDestinationResult_lo_hi_hi_lo_52};
  wire [7:0]    maskDestinationResult_lo_hi_54 = {maskDestinationResult_lo_hi_hi_53, maskDestinationResult_lo_hi_lo_53};
  wire [15:0]   maskDestinationResult_lo_310 = {maskDestinationResult_lo_hi_54, maskDestinationResult_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_52 = {sourceDataVec_17[28], sourceDataVec_16[28]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_52 = {sourceDataVec_19[28], sourceDataVec_18[28]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_53 = {maskDestinationResult_hi_lo_lo_hi_52, maskDestinationResult_hi_lo_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_52 = {sourceDataVec_21[28], sourceDataVec_20[28]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_52 = {sourceDataVec_23[28], sourceDataVec_22[28]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_53 = {maskDestinationResult_hi_lo_hi_hi_52, maskDestinationResult_hi_lo_hi_lo_52};
  wire [7:0]    maskDestinationResult_hi_lo_54 = {maskDestinationResult_hi_lo_hi_53, maskDestinationResult_hi_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_52 = {sourceDataVec_25[28], sourceDataVec_24[28]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_52 = {sourceDataVec_27[28], sourceDataVec_26[28]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_53 = {maskDestinationResult_hi_hi_lo_hi_52, maskDestinationResult_hi_hi_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_52 = {sourceDataVec_29[28], sourceDataVec_28[28]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_52 = {sourceDataVec_31[28], sourceDataVec_30[28]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_53 = {maskDestinationResult_hi_hi_hi_hi_52, maskDestinationResult_hi_hi_hi_lo_52};
  wire [7:0]    maskDestinationResult_hi_hi_54 = {maskDestinationResult_hi_hi_hi_53, maskDestinationResult_hi_hi_lo_53};
  wire [15:0]   maskDestinationResult_hi_310 = {maskDestinationResult_hi_hi_54, maskDestinationResult_hi_lo_54};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_53 = {sourceDataVec_1[29], sourceDataVec_0[29]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_53 = {sourceDataVec_3[29], sourceDataVec_2[29]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_54 = {maskDestinationResult_lo_lo_lo_hi_53, maskDestinationResult_lo_lo_lo_lo_53};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_53 = {sourceDataVec_5[29], sourceDataVec_4[29]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_53 = {sourceDataVec_7[29], sourceDataVec_6[29]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_54 = {maskDestinationResult_lo_lo_hi_hi_53, maskDestinationResult_lo_lo_hi_lo_53};
  wire [7:0]    maskDestinationResult_lo_lo_55 = {maskDestinationResult_lo_lo_hi_54, maskDestinationResult_lo_lo_lo_54};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_53 = {sourceDataVec_9[29], sourceDataVec_8[29]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_53 = {sourceDataVec_11[29], sourceDataVec_10[29]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_54 = {maskDestinationResult_lo_hi_lo_hi_53, maskDestinationResult_lo_hi_lo_lo_53};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_53 = {sourceDataVec_13[29], sourceDataVec_12[29]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_53 = {sourceDataVec_15[29], sourceDataVec_14[29]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_54 = {maskDestinationResult_lo_hi_hi_hi_53, maskDestinationResult_lo_hi_hi_lo_53};
  wire [7:0]    maskDestinationResult_lo_hi_55 = {maskDestinationResult_lo_hi_hi_54, maskDestinationResult_lo_hi_lo_54};
  wire [15:0]   maskDestinationResult_lo_311 = {maskDestinationResult_lo_hi_55, maskDestinationResult_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_53 = {sourceDataVec_17[29], sourceDataVec_16[29]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_53 = {sourceDataVec_19[29], sourceDataVec_18[29]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_54 = {maskDestinationResult_hi_lo_lo_hi_53, maskDestinationResult_hi_lo_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_53 = {sourceDataVec_21[29], sourceDataVec_20[29]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_53 = {sourceDataVec_23[29], sourceDataVec_22[29]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_54 = {maskDestinationResult_hi_lo_hi_hi_53, maskDestinationResult_hi_lo_hi_lo_53};
  wire [7:0]    maskDestinationResult_hi_lo_55 = {maskDestinationResult_hi_lo_hi_54, maskDestinationResult_hi_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_53 = {sourceDataVec_25[29], sourceDataVec_24[29]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_53 = {sourceDataVec_27[29], sourceDataVec_26[29]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_54 = {maskDestinationResult_hi_hi_lo_hi_53, maskDestinationResult_hi_hi_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_53 = {sourceDataVec_29[29], sourceDataVec_28[29]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_53 = {sourceDataVec_31[29], sourceDataVec_30[29]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_54 = {maskDestinationResult_hi_hi_hi_hi_53, maskDestinationResult_hi_hi_hi_lo_53};
  wire [7:0]    maskDestinationResult_hi_hi_55 = {maskDestinationResult_hi_hi_hi_54, maskDestinationResult_hi_hi_lo_54};
  wire [15:0]   maskDestinationResult_hi_311 = {maskDestinationResult_hi_hi_55, maskDestinationResult_hi_lo_55};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_54 = {sourceDataVec_1[30], sourceDataVec_0[30]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_54 = {sourceDataVec_3[30], sourceDataVec_2[30]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_55 = {maskDestinationResult_lo_lo_lo_hi_54, maskDestinationResult_lo_lo_lo_lo_54};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_54 = {sourceDataVec_5[30], sourceDataVec_4[30]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_54 = {sourceDataVec_7[30], sourceDataVec_6[30]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_55 = {maskDestinationResult_lo_lo_hi_hi_54, maskDestinationResult_lo_lo_hi_lo_54};
  wire [7:0]    maskDestinationResult_lo_lo_56 = {maskDestinationResult_lo_lo_hi_55, maskDestinationResult_lo_lo_lo_55};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_54 = {sourceDataVec_9[30], sourceDataVec_8[30]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_54 = {sourceDataVec_11[30], sourceDataVec_10[30]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_55 = {maskDestinationResult_lo_hi_lo_hi_54, maskDestinationResult_lo_hi_lo_lo_54};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_54 = {sourceDataVec_13[30], sourceDataVec_12[30]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_54 = {sourceDataVec_15[30], sourceDataVec_14[30]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_55 = {maskDestinationResult_lo_hi_hi_hi_54, maskDestinationResult_lo_hi_hi_lo_54};
  wire [7:0]    maskDestinationResult_lo_hi_56 = {maskDestinationResult_lo_hi_hi_55, maskDestinationResult_lo_hi_lo_55};
  wire [15:0]   maskDestinationResult_lo_312 = {maskDestinationResult_lo_hi_56, maskDestinationResult_lo_lo_56};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_54 = {sourceDataVec_17[30], sourceDataVec_16[30]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_54 = {sourceDataVec_19[30], sourceDataVec_18[30]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_55 = {maskDestinationResult_hi_lo_lo_hi_54, maskDestinationResult_hi_lo_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_54 = {sourceDataVec_21[30], sourceDataVec_20[30]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_54 = {sourceDataVec_23[30], sourceDataVec_22[30]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_55 = {maskDestinationResult_hi_lo_hi_hi_54, maskDestinationResult_hi_lo_hi_lo_54};
  wire [7:0]    maskDestinationResult_hi_lo_56 = {maskDestinationResult_hi_lo_hi_55, maskDestinationResult_hi_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_54 = {sourceDataVec_25[30], sourceDataVec_24[30]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_54 = {sourceDataVec_27[30], sourceDataVec_26[30]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_55 = {maskDestinationResult_hi_hi_lo_hi_54, maskDestinationResult_hi_hi_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_54 = {sourceDataVec_29[30], sourceDataVec_28[30]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_54 = {sourceDataVec_31[30], sourceDataVec_30[30]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_55 = {maskDestinationResult_hi_hi_hi_hi_54, maskDestinationResult_hi_hi_hi_lo_54};
  wire [7:0]    maskDestinationResult_hi_hi_56 = {maskDestinationResult_hi_hi_hi_55, maskDestinationResult_hi_hi_lo_55};
  wire [15:0]   maskDestinationResult_hi_312 = {maskDestinationResult_hi_hi_56, maskDestinationResult_hi_lo_56};
  wire [1:0]    maskDestinationResult_lo_lo_lo_lo_55 = {sourceDataVec_1[31], sourceDataVec_0[31]};
  wire [1:0]    maskDestinationResult_lo_lo_lo_hi_55 = {sourceDataVec_3[31], sourceDataVec_2[31]};
  wire [3:0]    maskDestinationResult_lo_lo_lo_56 = {maskDestinationResult_lo_lo_lo_hi_55, maskDestinationResult_lo_lo_lo_lo_55};
  wire [1:0]    maskDestinationResult_lo_lo_hi_lo_55 = {sourceDataVec_5[31], sourceDataVec_4[31]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_hi_55 = {sourceDataVec_7[31], sourceDataVec_6[31]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_56 = {maskDestinationResult_lo_lo_hi_hi_55, maskDestinationResult_lo_lo_hi_lo_55};
  wire [7:0]    maskDestinationResult_lo_lo_57 = {maskDestinationResult_lo_lo_hi_56, maskDestinationResult_lo_lo_lo_56};
  wire [1:0]    maskDestinationResult_lo_hi_lo_lo_55 = {sourceDataVec_9[31], sourceDataVec_8[31]};
  wire [1:0]    maskDestinationResult_lo_hi_lo_hi_55 = {sourceDataVec_11[31], sourceDataVec_10[31]};
  wire [3:0]    maskDestinationResult_lo_hi_lo_56 = {maskDestinationResult_lo_hi_lo_hi_55, maskDestinationResult_lo_hi_lo_lo_55};
  wire [1:0]    maskDestinationResult_lo_hi_hi_lo_55 = {sourceDataVec_13[31], sourceDataVec_12[31]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_hi_55 = {sourceDataVec_15[31], sourceDataVec_14[31]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_56 = {maskDestinationResult_lo_hi_hi_hi_55, maskDestinationResult_lo_hi_hi_lo_55};
  wire [7:0]    maskDestinationResult_lo_hi_57 = {maskDestinationResult_lo_hi_hi_56, maskDestinationResult_lo_hi_lo_56};
  wire [15:0]   maskDestinationResult_lo_313 = {maskDestinationResult_lo_hi_57, maskDestinationResult_lo_lo_57};
  wire [1:0]    maskDestinationResult_hi_lo_lo_lo_55 = {sourceDataVec_17[31], sourceDataVec_16[31]};
  wire [1:0]    maskDestinationResult_hi_lo_lo_hi_55 = {sourceDataVec_19[31], sourceDataVec_18[31]};
  wire [3:0]    maskDestinationResult_hi_lo_lo_56 = {maskDestinationResult_hi_lo_lo_hi_55, maskDestinationResult_hi_lo_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_lo_hi_lo_55 = {sourceDataVec_21[31], sourceDataVec_20[31]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_hi_55 = {sourceDataVec_23[31], sourceDataVec_22[31]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_56 = {maskDestinationResult_hi_lo_hi_hi_55, maskDestinationResult_hi_lo_hi_lo_55};
  wire [7:0]    maskDestinationResult_hi_lo_57 = {maskDestinationResult_hi_lo_hi_56, maskDestinationResult_hi_lo_lo_56};
  wire [1:0]    maskDestinationResult_hi_hi_lo_lo_55 = {sourceDataVec_25[31], sourceDataVec_24[31]};
  wire [1:0]    maskDestinationResult_hi_hi_lo_hi_55 = {sourceDataVec_27[31], sourceDataVec_26[31]};
  wire [3:0]    maskDestinationResult_hi_hi_lo_56 = {maskDestinationResult_hi_hi_lo_hi_55, maskDestinationResult_hi_hi_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_hi_hi_lo_55 = {sourceDataVec_29[31], sourceDataVec_28[31]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_hi_55 = {sourceDataVec_31[31], sourceDataVec_30[31]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_56 = {maskDestinationResult_hi_hi_hi_hi_55, maskDestinationResult_hi_hi_hi_lo_55};
  wire [7:0]    maskDestinationResult_hi_hi_57 = {maskDestinationResult_hi_hi_hi_56, maskDestinationResult_hi_hi_lo_56};
  wire [15:0]   maskDestinationResult_hi_313 = {maskDestinationResult_hi_hi_57, maskDestinationResult_hi_lo_57};
  wire [63:0]   maskDestinationResult_lo_lo_lo_lo_56 = {maskDestinationResult_hi_283, maskDestinationResult_lo_283, maskDestinationResult_hi_282, maskDestinationResult_lo_282};
  wire [63:0]   maskDestinationResult_lo_lo_lo_hi_56 = {maskDestinationResult_hi_285, maskDestinationResult_lo_285, maskDestinationResult_hi_284, maskDestinationResult_lo_284};
  wire [127:0]  maskDestinationResult_lo_lo_lo_57 = {maskDestinationResult_lo_lo_lo_hi_56, maskDestinationResult_lo_lo_lo_lo_56};
  wire [63:0]   maskDestinationResult_lo_lo_hi_lo_56 = {maskDestinationResult_hi_287, maskDestinationResult_lo_287, maskDestinationResult_hi_286, maskDestinationResult_lo_286};
  wire [63:0]   maskDestinationResult_lo_lo_hi_hi_56 = {maskDestinationResult_hi_289, maskDestinationResult_lo_289, maskDestinationResult_hi_288, maskDestinationResult_lo_288};
  wire [127:0]  maskDestinationResult_lo_lo_hi_57 = {maskDestinationResult_lo_lo_hi_hi_56, maskDestinationResult_lo_lo_hi_lo_56};
  wire [255:0]  maskDestinationResult_lo_lo_58 = {maskDestinationResult_lo_lo_hi_57, maskDestinationResult_lo_lo_lo_57};
  wire [63:0]   maskDestinationResult_lo_hi_lo_lo_56 = {maskDestinationResult_hi_291, maskDestinationResult_lo_291, maskDestinationResult_hi_290, maskDestinationResult_lo_290};
  wire [63:0]   maskDestinationResult_lo_hi_lo_hi_56 = {maskDestinationResult_hi_293, maskDestinationResult_lo_293, maskDestinationResult_hi_292, maskDestinationResult_lo_292};
  wire [127:0]  maskDestinationResult_lo_hi_lo_57 = {maskDestinationResult_lo_hi_lo_hi_56, maskDestinationResult_lo_hi_lo_lo_56};
  wire [63:0]   maskDestinationResult_lo_hi_hi_lo_56 = {maskDestinationResult_hi_295, maskDestinationResult_lo_295, maskDestinationResult_hi_294, maskDestinationResult_lo_294};
  wire [63:0]   maskDestinationResult_lo_hi_hi_hi_56 = {maskDestinationResult_hi_297, maskDestinationResult_lo_297, maskDestinationResult_hi_296, maskDestinationResult_lo_296};
  wire [127:0]  maskDestinationResult_lo_hi_hi_57 = {maskDestinationResult_lo_hi_hi_hi_56, maskDestinationResult_lo_hi_hi_lo_56};
  wire [255:0]  maskDestinationResult_lo_hi_58 = {maskDestinationResult_lo_hi_hi_57, maskDestinationResult_lo_hi_lo_57};
  wire [511:0]  maskDestinationResult_lo_314 = {maskDestinationResult_lo_hi_58, maskDestinationResult_lo_lo_58};
  wire [63:0]   maskDestinationResult_hi_lo_lo_lo_56 = {maskDestinationResult_hi_299, maskDestinationResult_lo_299, maskDestinationResult_hi_298, maskDestinationResult_lo_298};
  wire [63:0]   maskDestinationResult_hi_lo_lo_hi_56 = {maskDestinationResult_hi_301, maskDestinationResult_lo_301, maskDestinationResult_hi_300, maskDestinationResult_lo_300};
  wire [127:0]  maskDestinationResult_hi_lo_lo_57 = {maskDestinationResult_hi_lo_lo_hi_56, maskDestinationResult_hi_lo_lo_lo_56};
  wire [63:0]   maskDestinationResult_hi_lo_hi_lo_56 = {maskDestinationResult_hi_303, maskDestinationResult_lo_303, maskDestinationResult_hi_302, maskDestinationResult_lo_302};
  wire [63:0]   maskDestinationResult_hi_lo_hi_hi_56 = {maskDestinationResult_hi_305, maskDestinationResult_lo_305, maskDestinationResult_hi_304, maskDestinationResult_lo_304};
  wire [127:0]  maskDestinationResult_hi_lo_hi_57 = {maskDestinationResult_hi_lo_hi_hi_56, maskDestinationResult_hi_lo_hi_lo_56};
  wire [255:0]  maskDestinationResult_hi_lo_58 = {maskDestinationResult_hi_lo_hi_57, maskDestinationResult_hi_lo_lo_57};
  wire [63:0]   maskDestinationResult_hi_hi_lo_lo_56 = {maskDestinationResult_hi_307, maskDestinationResult_lo_307, maskDestinationResult_hi_306, maskDestinationResult_lo_306};
  wire [63:0]   maskDestinationResult_hi_hi_lo_hi_56 = {maskDestinationResult_hi_309, maskDestinationResult_lo_309, maskDestinationResult_hi_308, maskDestinationResult_lo_308};
  wire [127:0]  maskDestinationResult_hi_hi_lo_57 = {maskDestinationResult_hi_hi_lo_hi_56, maskDestinationResult_hi_hi_lo_lo_56};
  wire [63:0]   maskDestinationResult_hi_hi_hi_lo_56 = {maskDestinationResult_hi_311, maskDestinationResult_lo_311, maskDestinationResult_hi_310, maskDestinationResult_lo_310};
  wire [63:0]   maskDestinationResult_hi_hi_hi_hi_56 = {maskDestinationResult_hi_313, maskDestinationResult_lo_313, maskDestinationResult_hi_312, maskDestinationResult_lo_312};
  wire [127:0]  maskDestinationResult_hi_hi_hi_57 = {maskDestinationResult_hi_hi_hi_hi_56, maskDestinationResult_hi_hi_hi_lo_56};
  wire [255:0]  maskDestinationResult_hi_hi_58 = {maskDestinationResult_hi_hi_hi_57, maskDestinationResult_hi_hi_lo_57};
  wire [511:0]  maskDestinationResult_hi_314 = {maskDestinationResult_hi_hi_58, maskDestinationResult_hi_lo_58};
  wire [1023:0] maskDestinationResult =
    (eew1H[0] ? {maskDestinationResult_hi_264, maskDestinationResult_lo_264} : 1024'h0) | (eew1H[1] ? {maskDestinationResult_hi_281, maskDestinationResult_lo_281} : 1024'h0)
    | (eew1H[2] ? {maskDestinationResult_hi_314, maskDestinationResult_lo_314} : 1024'h0);
  wire          sign = in_uop[0];
  wire          extendRatio = in_uop[2];
  wire [3:0]    _source2_T_1 = 4'h1 << in_groupCounter[1:0];
  wire [1:0]    _source2_T_18 = 2'h1 << in_groupCounter[0];
  wire [511:0]  source2 =
    extendRatio
      ? {256'h0, (_source2_T_1[0] ? in_source2[255:0] : 256'h0) | (_source2_T_1[1] ? in_source2[511:256] : 256'h0) | (_source2_T_1[2] ? in_source2[767:512] : 256'h0) | (_source2_T_1[3] ? in_source2[1023:768] : 256'h0)}
      : (_source2_T_18[0] ? in_source2[511:0] : 512'h0) | (_source2_T_18[1] ? in_source2[1023:512] : 512'h0);
  wire [1:0]    _extendResult_T_969 = 2'h1 << extendRatio;
  wire [31:0]   extendResult_lo_lo_lo_lo_lo = {{8{source2[15] & sign}}, source2[15:8], {8{source2[7] & sign}}, source2[7:0]};
  wire [31:0]   extendResult_lo_lo_lo_lo_hi = {{8{source2[31] & sign}}, source2[31:24], {8{source2[23] & sign}}, source2[23:16]};
  wire [63:0]   extendResult_lo_lo_lo_lo = {extendResult_lo_lo_lo_lo_hi, extendResult_lo_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_lo_hi_lo = {{8{source2[47] & sign}}, source2[47:40], {8{source2[39] & sign}}, source2[39:32]};
  wire [31:0]   extendResult_lo_lo_lo_hi_hi = {{8{source2[63] & sign}}, source2[63:56], {8{source2[55] & sign}}, source2[55:48]};
  wire [63:0]   extendResult_lo_lo_lo_hi = {extendResult_lo_lo_lo_hi_hi, extendResult_lo_lo_lo_hi_lo};
  wire [127:0]  extendResult_lo_lo_lo = {extendResult_lo_lo_lo_hi, extendResult_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_lo_lo = {{8{source2[79] & sign}}, source2[79:72], {8{source2[71] & sign}}, source2[71:64]};
  wire [31:0]   extendResult_lo_lo_hi_lo_hi = {{8{source2[95] & sign}}, source2[95:88], {8{source2[87] & sign}}, source2[87:80]};
  wire [63:0]   extendResult_lo_lo_hi_lo = {extendResult_lo_lo_hi_lo_hi, extendResult_lo_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_hi_lo = {{8{source2[111] & sign}}, source2[111:104], {8{source2[103] & sign}}, source2[103:96]};
  wire [31:0]   extendResult_lo_lo_hi_hi_hi = {{8{source2[127] & sign}}, source2[127:120], {8{source2[119] & sign}}, source2[119:112]};
  wire [63:0]   extendResult_lo_lo_hi_hi = {extendResult_lo_lo_hi_hi_hi, extendResult_lo_lo_hi_hi_lo};
  wire [127:0]  extendResult_lo_lo_hi = {extendResult_lo_lo_hi_hi, extendResult_lo_lo_hi_lo};
  wire [255:0]  extendResult_lo_lo = {extendResult_lo_lo_hi, extendResult_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_lo_lo = {{8{source2[143] & sign}}, source2[143:136], {8{source2[135] & sign}}, source2[135:128]};
  wire [31:0]   extendResult_lo_hi_lo_lo_hi = {{8{source2[159] & sign}}, source2[159:152], {8{source2[151] & sign}}, source2[151:144]};
  wire [63:0]   extendResult_lo_hi_lo_lo = {extendResult_lo_hi_lo_lo_hi, extendResult_lo_hi_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_hi_lo = {{8{source2[175] & sign}}, source2[175:168], {8{source2[167] & sign}}, source2[167:160]};
  wire [31:0]   extendResult_lo_hi_lo_hi_hi = {{8{source2[191] & sign}}, source2[191:184], {8{source2[183] & sign}}, source2[183:176]};
  wire [63:0]   extendResult_lo_hi_lo_hi = {extendResult_lo_hi_lo_hi_hi, extendResult_lo_hi_lo_hi_lo};
  wire [127:0]  extendResult_lo_hi_lo = {extendResult_lo_hi_lo_hi, extendResult_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_lo_lo = {{8{source2[207] & sign}}, source2[207:200], {8{source2[199] & sign}}, source2[199:192]};
  wire [31:0]   extendResult_lo_hi_hi_lo_hi = {{8{source2[223] & sign}}, source2[223:216], {8{source2[215] & sign}}, source2[215:208]};
  wire [63:0]   extendResult_lo_hi_hi_lo = {extendResult_lo_hi_hi_lo_hi, extendResult_lo_hi_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_hi_lo = {{8{source2[239] & sign}}, source2[239:232], {8{source2[231] & sign}}, source2[231:224]};
  wire [31:0]   extendResult_lo_hi_hi_hi_hi = {{8{source2[255] & sign}}, source2[255:248], {8{source2[247] & sign}}, source2[247:240]};
  wire [63:0]   extendResult_lo_hi_hi_hi = {extendResult_lo_hi_hi_hi_hi, extendResult_lo_hi_hi_hi_lo};
  wire [127:0]  extendResult_lo_hi_hi = {extendResult_lo_hi_hi_hi, extendResult_lo_hi_hi_lo};
  wire [255:0]  extendResult_lo_hi = {extendResult_lo_hi_hi, extendResult_lo_hi_lo};
  wire [511:0]  extendResult_lo = {extendResult_lo_hi, extendResult_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_lo_lo = {{8{source2[271] & sign}}, source2[271:264], {8{source2[263] & sign}}, source2[263:256]};
  wire [31:0]   extendResult_hi_lo_lo_lo_hi = {{8{source2[287] & sign}}, source2[287:280], {8{source2[279] & sign}}, source2[279:272]};
  wire [63:0]   extendResult_hi_lo_lo_lo = {extendResult_hi_lo_lo_lo_hi, extendResult_hi_lo_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_hi_lo = {{8{source2[303] & sign}}, source2[303:296], {8{source2[295] & sign}}, source2[295:288]};
  wire [31:0]   extendResult_hi_lo_lo_hi_hi = {{8{source2[319] & sign}}, source2[319:312], {8{source2[311] & sign}}, source2[311:304]};
  wire [63:0]   extendResult_hi_lo_lo_hi = {extendResult_hi_lo_lo_hi_hi, extendResult_hi_lo_lo_hi_lo};
  wire [127:0]  extendResult_hi_lo_lo = {extendResult_hi_lo_lo_hi, extendResult_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_lo_lo = {{8{source2[335] & sign}}, source2[335:328], {8{source2[327] & sign}}, source2[327:320]};
  wire [31:0]   extendResult_hi_lo_hi_lo_hi = {{8{source2[351] & sign}}, source2[351:344], {8{source2[343] & sign}}, source2[343:336]};
  wire [63:0]   extendResult_hi_lo_hi_lo = {extendResult_hi_lo_hi_lo_hi, extendResult_hi_lo_hi_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_hi_lo = {{8{source2[367] & sign}}, source2[367:360], {8{source2[359] & sign}}, source2[359:352]};
  wire [31:0]   extendResult_hi_lo_hi_hi_hi = {{8{source2[383] & sign}}, source2[383:376], {8{source2[375] & sign}}, source2[375:368]};
  wire [63:0]   extendResult_hi_lo_hi_hi = {extendResult_hi_lo_hi_hi_hi, extendResult_hi_lo_hi_hi_lo};
  wire [127:0]  extendResult_hi_lo_hi = {extendResult_hi_lo_hi_hi, extendResult_hi_lo_hi_lo};
  wire [255:0]  extendResult_hi_lo = {extendResult_hi_lo_hi, extendResult_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_lo_lo = {{8{source2[399] & sign}}, source2[399:392], {8{source2[391] & sign}}, source2[391:384]};
  wire [31:0]   extendResult_hi_hi_lo_lo_hi = {{8{source2[415] & sign}}, source2[415:408], {8{source2[407] & sign}}, source2[407:400]};
  wire [63:0]   extendResult_hi_hi_lo_lo = {extendResult_hi_hi_lo_lo_hi, extendResult_hi_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_hi_lo = {{8{source2[431] & sign}}, source2[431:424], {8{source2[423] & sign}}, source2[423:416]};
  wire [31:0]   extendResult_hi_hi_lo_hi_hi = {{8{source2[447] & sign}}, source2[447:440], {8{source2[439] & sign}}, source2[439:432]};
  wire [63:0]   extendResult_hi_hi_lo_hi = {extendResult_hi_hi_lo_hi_hi, extendResult_hi_hi_lo_hi_lo};
  wire [127:0]  extendResult_hi_hi_lo = {extendResult_hi_hi_lo_hi, extendResult_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_lo_lo = {{8{source2[463] & sign}}, source2[463:456], {8{source2[455] & sign}}, source2[455:448]};
  wire [31:0]   extendResult_hi_hi_hi_lo_hi = {{8{source2[479] & sign}}, source2[479:472], {8{source2[471] & sign}}, source2[471:464]};
  wire [63:0]   extendResult_hi_hi_hi_lo = {extendResult_hi_hi_hi_lo_hi, extendResult_hi_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_hi_lo = {{8{source2[495] & sign}}, source2[495:488], {8{source2[487] & sign}}, source2[487:480]};
  wire [31:0]   extendResult_hi_hi_hi_hi_hi = {{8{source2[511] & sign}}, source2[511:504], {8{source2[503] & sign}}, source2[503:496]};
  wire [63:0]   extendResult_hi_hi_hi_hi = {extendResult_hi_hi_hi_hi_hi, extendResult_hi_hi_hi_hi_lo};
  wire [127:0]  extendResult_hi_hi_hi = {extendResult_hi_hi_hi_hi, extendResult_hi_hi_hi_lo};
  wire [255:0]  extendResult_hi_hi = {extendResult_hi_hi_hi, extendResult_hi_hi_lo};
  wire [511:0]  extendResult_hi = {extendResult_hi_hi, extendResult_hi_lo};
  wire [31:0]   extendResult_lo_lo_lo_lo_lo_lo = {{12{source2[7] & sign}}, source2[7:4], {12{source2[3] & sign}}, source2[3:0]};
  wire [31:0]   extendResult_lo_lo_lo_lo_lo_hi = {{12{source2[15] & sign}}, source2[15:12], {12{source2[11] & sign}}, source2[11:8]};
  wire [63:0]   extendResult_lo_lo_lo_lo_lo_1 = {extendResult_lo_lo_lo_lo_lo_hi, extendResult_lo_lo_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_lo_lo_hi_lo = {{12{source2[23] & sign}}, source2[23:20], {12{source2[19] & sign}}, source2[19:16]};
  wire [31:0]   extendResult_lo_lo_lo_lo_hi_hi = {{12{source2[31] & sign}}, source2[31:28], {12{source2[27] & sign}}, source2[27:24]};
  wire [63:0]   extendResult_lo_lo_lo_lo_hi_1 = {extendResult_lo_lo_lo_lo_hi_hi, extendResult_lo_lo_lo_lo_hi_lo};
  wire [127:0]  extendResult_lo_lo_lo_lo_1 = {extendResult_lo_lo_lo_lo_hi_1, extendResult_lo_lo_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_lo_lo_hi_lo_lo = {{12{source2[39] & sign}}, source2[39:36], {12{source2[35] & sign}}, source2[35:32]};
  wire [31:0]   extendResult_lo_lo_lo_hi_lo_hi = {{12{source2[47] & sign}}, source2[47:44], {12{source2[43] & sign}}, source2[43:40]};
  wire [63:0]   extendResult_lo_lo_lo_hi_lo_1 = {extendResult_lo_lo_lo_hi_lo_hi, extendResult_lo_lo_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_lo_lo_hi_hi_lo = {{12{source2[55] & sign}}, source2[55:52], {12{source2[51] & sign}}, source2[51:48]};
  wire [31:0]   extendResult_lo_lo_lo_hi_hi_hi = {{12{source2[63] & sign}}, source2[63:60], {12{source2[59] & sign}}, source2[59:56]};
  wire [63:0]   extendResult_lo_lo_lo_hi_hi_1 = {extendResult_lo_lo_lo_hi_hi_hi, extendResult_lo_lo_lo_hi_hi_lo};
  wire [127:0]  extendResult_lo_lo_lo_hi_1 = {extendResult_lo_lo_lo_hi_hi_1, extendResult_lo_lo_lo_hi_lo_1};
  wire [255:0]  extendResult_lo_lo_lo_1 = {extendResult_lo_lo_lo_hi_1, extendResult_lo_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_lo_hi_lo_lo_lo = {{12{source2[71] & sign}}, source2[71:68], {12{source2[67] & sign}}, source2[67:64]};
  wire [31:0]   extendResult_lo_lo_hi_lo_lo_hi = {{12{source2[79] & sign}}, source2[79:76], {12{source2[75] & sign}}, source2[75:72]};
  wire [63:0]   extendResult_lo_lo_hi_lo_lo_1 = {extendResult_lo_lo_hi_lo_lo_hi, extendResult_lo_lo_hi_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_lo_hi_lo = {{12{source2[87] & sign}}, source2[87:84], {12{source2[83] & sign}}, source2[83:80]};
  wire [31:0]   extendResult_lo_lo_hi_lo_hi_hi = {{12{source2[95] & sign}}, source2[95:92], {12{source2[91] & sign}}, source2[91:88]};
  wire [63:0]   extendResult_lo_lo_hi_lo_hi_1 = {extendResult_lo_lo_hi_lo_hi_hi, extendResult_lo_lo_hi_lo_hi_lo};
  wire [127:0]  extendResult_lo_lo_hi_lo_1 = {extendResult_lo_lo_hi_lo_hi_1, extendResult_lo_lo_hi_lo_lo_1};
  wire [31:0]   extendResult_lo_lo_hi_hi_lo_lo = {{12{source2[103] & sign}}, source2[103:100], {12{source2[99] & sign}}, source2[99:96]};
  wire [31:0]   extendResult_lo_lo_hi_hi_lo_hi = {{12{source2[111] & sign}}, source2[111:108], {12{source2[107] & sign}}, source2[107:104]};
  wire [63:0]   extendResult_lo_lo_hi_hi_lo_1 = {extendResult_lo_lo_hi_hi_lo_hi, extendResult_lo_lo_hi_hi_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_hi_hi_lo = {{12{source2[119] & sign}}, source2[119:116], {12{source2[115] & sign}}, source2[115:112]};
  wire [31:0]   extendResult_lo_lo_hi_hi_hi_hi = {{12{source2[127] & sign}}, source2[127:124], {12{source2[123] & sign}}, source2[123:120]};
  wire [63:0]   extendResult_lo_lo_hi_hi_hi_1 = {extendResult_lo_lo_hi_hi_hi_hi, extendResult_lo_lo_hi_hi_hi_lo};
  wire [127:0]  extendResult_lo_lo_hi_hi_1 = {extendResult_lo_lo_hi_hi_hi_1, extendResult_lo_lo_hi_hi_lo_1};
  wire [255:0]  extendResult_lo_lo_hi_1 = {extendResult_lo_lo_hi_hi_1, extendResult_lo_lo_hi_lo_1};
  wire [511:0]  extendResult_lo_lo_1 = {extendResult_lo_lo_hi_1, extendResult_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_lo_lo_lo_lo = {{12{source2[135] & sign}}, source2[135:132], {12{source2[131] & sign}}, source2[131:128]};
  wire [31:0]   extendResult_lo_hi_lo_lo_lo_hi = {{12{source2[143] & sign}}, source2[143:140], {12{source2[139] & sign}}, source2[139:136]};
  wire [63:0]   extendResult_lo_hi_lo_lo_lo_1 = {extendResult_lo_hi_lo_lo_lo_hi, extendResult_lo_hi_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_lo_hi_lo = {{12{source2[151] & sign}}, source2[151:148], {12{source2[147] & sign}}, source2[147:144]};
  wire [31:0]   extendResult_lo_hi_lo_lo_hi_hi = {{12{source2[159] & sign}}, source2[159:156], {12{source2[155] & sign}}, source2[155:152]};
  wire [63:0]   extendResult_lo_hi_lo_lo_hi_1 = {extendResult_lo_hi_lo_lo_hi_hi, extendResult_lo_hi_lo_lo_hi_lo};
  wire [127:0]  extendResult_lo_hi_lo_lo_1 = {extendResult_lo_hi_lo_lo_hi_1, extendResult_lo_hi_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_lo_hi_lo_lo = {{12{source2[167] & sign}}, source2[167:164], {12{source2[163] & sign}}, source2[163:160]};
  wire [31:0]   extendResult_lo_hi_lo_hi_lo_hi = {{12{source2[175] & sign}}, source2[175:172], {12{source2[171] & sign}}, source2[171:168]};
  wire [63:0]   extendResult_lo_hi_lo_hi_lo_1 = {extendResult_lo_hi_lo_hi_lo_hi, extendResult_lo_hi_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_hi_hi_lo = {{12{source2[183] & sign}}, source2[183:180], {12{source2[179] & sign}}, source2[179:176]};
  wire [31:0]   extendResult_lo_hi_lo_hi_hi_hi = {{12{source2[191] & sign}}, source2[191:188], {12{source2[187] & sign}}, source2[187:184]};
  wire [63:0]   extendResult_lo_hi_lo_hi_hi_1 = {extendResult_lo_hi_lo_hi_hi_hi, extendResult_lo_hi_lo_hi_hi_lo};
  wire [127:0]  extendResult_lo_hi_lo_hi_1 = {extendResult_lo_hi_lo_hi_hi_1, extendResult_lo_hi_lo_hi_lo_1};
  wire [255:0]  extendResult_lo_hi_lo_1 = {extendResult_lo_hi_lo_hi_1, extendResult_lo_hi_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_hi_lo_lo_lo = {{12{source2[199] & sign}}, source2[199:196], {12{source2[195] & sign}}, source2[195:192]};
  wire [31:0]   extendResult_lo_hi_hi_lo_lo_hi = {{12{source2[207] & sign}}, source2[207:204], {12{source2[203] & sign}}, source2[203:200]};
  wire [63:0]   extendResult_lo_hi_hi_lo_lo_1 = {extendResult_lo_hi_hi_lo_lo_hi, extendResult_lo_hi_hi_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_lo_hi_lo = {{12{source2[215] & sign}}, source2[215:212], {12{source2[211] & sign}}, source2[211:208]};
  wire [31:0]   extendResult_lo_hi_hi_lo_hi_hi = {{12{source2[223] & sign}}, source2[223:220], {12{source2[219] & sign}}, source2[219:216]};
  wire [63:0]   extendResult_lo_hi_hi_lo_hi_1 = {extendResult_lo_hi_hi_lo_hi_hi, extendResult_lo_hi_hi_lo_hi_lo};
  wire [127:0]  extendResult_lo_hi_hi_lo_1 = {extendResult_lo_hi_hi_lo_hi_1, extendResult_lo_hi_hi_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_hi_hi_lo_lo = {{12{source2[231] & sign}}, source2[231:228], {12{source2[227] & sign}}, source2[227:224]};
  wire [31:0]   extendResult_lo_hi_hi_hi_lo_hi = {{12{source2[239] & sign}}, source2[239:236], {12{source2[235] & sign}}, source2[235:232]};
  wire [63:0]   extendResult_lo_hi_hi_hi_lo_1 = {extendResult_lo_hi_hi_hi_lo_hi, extendResult_lo_hi_hi_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_hi_hi_lo = {{12{source2[247] & sign}}, source2[247:244], {12{source2[243] & sign}}, source2[243:240]};
  wire [31:0]   extendResult_lo_hi_hi_hi_hi_hi = {{12{source2[255] & sign}}, source2[255:252], {12{source2[251] & sign}}, source2[251:248]};
  wire [63:0]   extendResult_lo_hi_hi_hi_hi_1 = {extendResult_lo_hi_hi_hi_hi_hi, extendResult_lo_hi_hi_hi_hi_lo};
  wire [127:0]  extendResult_lo_hi_hi_hi_1 = {extendResult_lo_hi_hi_hi_hi_1, extendResult_lo_hi_hi_hi_lo_1};
  wire [255:0]  extendResult_lo_hi_hi_1 = {extendResult_lo_hi_hi_hi_1, extendResult_lo_hi_hi_lo_1};
  wire [511:0]  extendResult_lo_hi_1 = {extendResult_lo_hi_hi_1, extendResult_lo_hi_lo_1};
  wire [1023:0] extendResult_lo_1 = {extendResult_lo_hi_1, extendResult_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_lo_lo_lo_lo = {{12{source2[263] & sign}}, source2[263:260], {12{source2[259] & sign}}, source2[259:256]};
  wire [31:0]   extendResult_hi_lo_lo_lo_lo_hi = {{12{source2[271] & sign}}, source2[271:268], {12{source2[267] & sign}}, source2[267:264]};
  wire [63:0]   extendResult_hi_lo_lo_lo_lo_1 = {extendResult_hi_lo_lo_lo_lo_hi, extendResult_hi_lo_lo_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_lo_hi_lo = {{12{source2[279] & sign}}, source2[279:276], {12{source2[275] & sign}}, source2[275:272]};
  wire [31:0]   extendResult_hi_lo_lo_lo_hi_hi = {{12{source2[287] & sign}}, source2[287:284], {12{source2[283] & sign}}, source2[283:280]};
  wire [63:0]   extendResult_hi_lo_lo_lo_hi_1 = {extendResult_hi_lo_lo_lo_hi_hi, extendResult_hi_lo_lo_lo_hi_lo};
  wire [127:0]  extendResult_hi_lo_lo_lo_1 = {extendResult_hi_lo_lo_lo_hi_1, extendResult_hi_lo_lo_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_lo_hi_lo_lo = {{12{source2[295] & sign}}, source2[295:292], {12{source2[291] & sign}}, source2[291:288]};
  wire [31:0]   extendResult_hi_lo_lo_hi_lo_hi = {{12{source2[303] & sign}}, source2[303:300], {12{source2[299] & sign}}, source2[299:296]};
  wire [63:0]   extendResult_hi_lo_lo_hi_lo_1 = {extendResult_hi_lo_lo_hi_lo_hi, extendResult_hi_lo_lo_hi_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_hi_hi_lo = {{12{source2[311] & sign}}, source2[311:308], {12{source2[307] & sign}}, source2[307:304]};
  wire [31:0]   extendResult_hi_lo_lo_hi_hi_hi = {{12{source2[319] & sign}}, source2[319:316], {12{source2[315] & sign}}, source2[315:312]};
  wire [63:0]   extendResult_hi_lo_lo_hi_hi_1 = {extendResult_hi_lo_lo_hi_hi_hi, extendResult_hi_lo_lo_hi_hi_lo};
  wire [127:0]  extendResult_hi_lo_lo_hi_1 = {extendResult_hi_lo_lo_hi_hi_1, extendResult_hi_lo_lo_hi_lo_1};
  wire [255:0]  extendResult_hi_lo_lo_1 = {extendResult_hi_lo_lo_hi_1, extendResult_hi_lo_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_hi_lo_lo_lo = {{12{source2[327] & sign}}, source2[327:324], {12{source2[323] & sign}}, source2[323:320]};
  wire [31:0]   extendResult_hi_lo_hi_lo_lo_hi = {{12{source2[335] & sign}}, source2[335:332], {12{source2[331] & sign}}, source2[331:328]};
  wire [63:0]   extendResult_hi_lo_hi_lo_lo_1 = {extendResult_hi_lo_hi_lo_lo_hi, extendResult_hi_lo_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_lo_hi_lo = {{12{source2[343] & sign}}, source2[343:340], {12{source2[339] & sign}}, source2[339:336]};
  wire [31:0]   extendResult_hi_lo_hi_lo_hi_hi = {{12{source2[351] & sign}}, source2[351:348], {12{source2[347] & sign}}, source2[347:344]};
  wire [63:0]   extendResult_hi_lo_hi_lo_hi_1 = {extendResult_hi_lo_hi_lo_hi_hi, extendResult_hi_lo_hi_lo_hi_lo};
  wire [127:0]  extendResult_hi_lo_hi_lo_1 = {extendResult_hi_lo_hi_lo_hi_1, extendResult_hi_lo_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_hi_hi_lo_lo = {{12{source2[359] & sign}}, source2[359:356], {12{source2[355] & sign}}, source2[355:352]};
  wire [31:0]   extendResult_hi_lo_hi_hi_lo_hi = {{12{source2[367] & sign}}, source2[367:364], {12{source2[363] & sign}}, source2[363:360]};
  wire [63:0]   extendResult_hi_lo_hi_hi_lo_1 = {extendResult_hi_lo_hi_hi_lo_hi, extendResult_hi_lo_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_hi_hi_lo = {{12{source2[375] & sign}}, source2[375:372], {12{source2[371] & sign}}, source2[371:368]};
  wire [31:0]   extendResult_hi_lo_hi_hi_hi_hi = {{12{source2[383] & sign}}, source2[383:380], {12{source2[379] & sign}}, source2[379:376]};
  wire [63:0]   extendResult_hi_lo_hi_hi_hi_1 = {extendResult_hi_lo_hi_hi_hi_hi, extendResult_hi_lo_hi_hi_hi_lo};
  wire [127:0]  extendResult_hi_lo_hi_hi_1 = {extendResult_hi_lo_hi_hi_hi_1, extendResult_hi_lo_hi_hi_lo_1};
  wire [255:0]  extendResult_hi_lo_hi_1 = {extendResult_hi_lo_hi_hi_1, extendResult_hi_lo_hi_lo_1};
  wire [511:0]  extendResult_hi_lo_1 = {extendResult_hi_lo_hi_1, extendResult_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_lo_lo_lo_lo = {{12{source2[391] & sign}}, source2[391:388], {12{source2[387] & sign}}, source2[387:384]};
  wire [31:0]   extendResult_hi_hi_lo_lo_lo_hi = {{12{source2[399] & sign}}, source2[399:396], {12{source2[395] & sign}}, source2[395:392]};
  wire [63:0]   extendResult_hi_hi_lo_lo_lo_1 = {extendResult_hi_hi_lo_lo_lo_hi, extendResult_hi_hi_lo_lo_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_lo_hi_lo = {{12{source2[407] & sign}}, source2[407:404], {12{source2[403] & sign}}, source2[403:400]};
  wire [31:0]   extendResult_hi_hi_lo_lo_hi_hi = {{12{source2[415] & sign}}, source2[415:412], {12{source2[411] & sign}}, source2[411:408]};
  wire [63:0]   extendResult_hi_hi_lo_lo_hi_1 = {extendResult_hi_hi_lo_lo_hi_hi, extendResult_hi_hi_lo_lo_hi_lo};
  wire [127:0]  extendResult_hi_hi_lo_lo_1 = {extendResult_hi_hi_lo_lo_hi_1, extendResult_hi_hi_lo_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_lo_hi_lo_lo = {{12{source2[423] & sign}}, source2[423:420], {12{source2[419] & sign}}, source2[419:416]};
  wire [31:0]   extendResult_hi_hi_lo_hi_lo_hi = {{12{source2[431] & sign}}, source2[431:428], {12{source2[427] & sign}}, source2[427:424]};
  wire [63:0]   extendResult_hi_hi_lo_hi_lo_1 = {extendResult_hi_hi_lo_hi_lo_hi, extendResult_hi_hi_lo_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_hi_hi_lo = {{12{source2[439] & sign}}, source2[439:436], {12{source2[435] & sign}}, source2[435:432]};
  wire [31:0]   extendResult_hi_hi_lo_hi_hi_hi = {{12{source2[447] & sign}}, source2[447:444], {12{source2[443] & sign}}, source2[443:440]};
  wire [63:0]   extendResult_hi_hi_lo_hi_hi_1 = {extendResult_hi_hi_lo_hi_hi_hi, extendResult_hi_hi_lo_hi_hi_lo};
  wire [127:0]  extendResult_hi_hi_lo_hi_1 = {extendResult_hi_hi_lo_hi_hi_1, extendResult_hi_hi_lo_hi_lo_1};
  wire [255:0]  extendResult_hi_hi_lo_1 = {extendResult_hi_hi_lo_hi_1, extendResult_hi_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_hi_lo_lo_lo = {{12{source2[455] & sign}}, source2[455:452], {12{source2[451] & sign}}, source2[451:448]};
  wire [31:0]   extendResult_hi_hi_hi_lo_lo_hi = {{12{source2[463] & sign}}, source2[463:460], {12{source2[459] & sign}}, source2[459:456]};
  wire [63:0]   extendResult_hi_hi_hi_lo_lo_1 = {extendResult_hi_hi_hi_lo_lo_hi, extendResult_hi_hi_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_lo_hi_lo = {{12{source2[471] & sign}}, source2[471:468], {12{source2[467] & sign}}, source2[467:464]};
  wire [31:0]   extendResult_hi_hi_hi_lo_hi_hi = {{12{source2[479] & sign}}, source2[479:476], {12{source2[475] & sign}}, source2[475:472]};
  wire [63:0]   extendResult_hi_hi_hi_lo_hi_1 = {extendResult_hi_hi_hi_lo_hi_hi, extendResult_hi_hi_hi_lo_hi_lo};
  wire [127:0]  extendResult_hi_hi_hi_lo_1 = {extendResult_hi_hi_hi_lo_hi_1, extendResult_hi_hi_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_hi_hi_lo_lo = {{12{source2[487] & sign}}, source2[487:484], {12{source2[483] & sign}}, source2[483:480]};
  wire [31:0]   extendResult_hi_hi_hi_hi_lo_hi = {{12{source2[495] & sign}}, source2[495:492], {12{source2[491] & sign}}, source2[491:488]};
  wire [63:0]   extendResult_hi_hi_hi_hi_lo_1 = {extendResult_hi_hi_hi_hi_lo_hi, extendResult_hi_hi_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_hi_hi_lo = {{12{source2[503] & sign}}, source2[503:500], {12{source2[499] & sign}}, source2[499:496]};
  wire [31:0]   extendResult_hi_hi_hi_hi_hi_hi = {{12{source2[511] & sign}}, source2[511:508], {12{source2[507] & sign}}, source2[507:504]};
  wire [63:0]   extendResult_hi_hi_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi_hi_hi, extendResult_hi_hi_hi_hi_hi_lo};
  wire [127:0]  extendResult_hi_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi_hi_1, extendResult_hi_hi_hi_hi_lo_1};
  wire [255:0]  extendResult_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi_1, extendResult_hi_hi_hi_lo_1};
  wire [511:0]  extendResult_hi_hi_1 = {extendResult_hi_hi_hi_1, extendResult_hi_hi_lo_1};
  wire [1023:0] extendResult_hi_1 = {extendResult_hi_hi_1, extendResult_hi_lo_1};
  wire [63:0]   extendResult_lo_lo_lo_lo_2 = {{16{source2[31] & sign}}, source2[31:16], {16{source2[15] & sign}}, source2[15:0]};
  wire [63:0]   extendResult_lo_lo_lo_hi_2 = {{16{source2[63] & sign}}, source2[63:48], {16{source2[47] & sign}}, source2[47:32]};
  wire [127:0]  extendResult_lo_lo_lo_2 = {extendResult_lo_lo_lo_hi_2, extendResult_lo_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_lo_hi_lo_2 = {{16{source2[95] & sign}}, source2[95:80], {16{source2[79] & sign}}, source2[79:64]};
  wire [63:0]   extendResult_lo_lo_hi_hi_2 = {{16{source2[127] & sign}}, source2[127:112], {16{source2[111] & sign}}, source2[111:96]};
  wire [127:0]  extendResult_lo_lo_hi_2 = {extendResult_lo_lo_hi_hi_2, extendResult_lo_lo_hi_lo_2};
  wire [255:0]  extendResult_lo_lo_2 = {extendResult_lo_lo_hi_2, extendResult_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_lo_lo_2 = {{16{source2[159] & sign}}, source2[159:144], {16{source2[143] & sign}}, source2[143:128]};
  wire [63:0]   extendResult_lo_hi_lo_hi_2 = {{16{source2[191] & sign}}, source2[191:176], {16{source2[175] & sign}}, source2[175:160]};
  wire [127:0]  extendResult_lo_hi_lo_2 = {extendResult_lo_hi_lo_hi_2, extendResult_lo_hi_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_hi_lo_2 = {{16{source2[223] & sign}}, source2[223:208], {16{source2[207] & sign}}, source2[207:192]};
  wire [63:0]   extendResult_lo_hi_hi_hi_2 = {{16{source2[255] & sign}}, source2[255:240], {16{source2[239] & sign}}, source2[239:224]};
  wire [127:0]  extendResult_lo_hi_hi_2 = {extendResult_lo_hi_hi_hi_2, extendResult_lo_hi_hi_lo_2};
  wire [255:0]  extendResult_lo_hi_2 = {extendResult_lo_hi_hi_2, extendResult_lo_hi_lo_2};
  wire [511:0]  extendResult_lo_2 = {extendResult_lo_hi_2, extendResult_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_lo_lo_2 = {{16{source2[287] & sign}}, source2[287:272], {16{source2[271] & sign}}, source2[271:256]};
  wire [63:0]   extendResult_hi_lo_lo_hi_2 = {{16{source2[319] & sign}}, source2[319:304], {16{source2[303] & sign}}, source2[303:288]};
  wire [127:0]  extendResult_hi_lo_lo_2 = {extendResult_hi_lo_lo_hi_2, extendResult_hi_lo_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_hi_lo_2 = {{16{source2[351] & sign}}, source2[351:336], {16{source2[335] & sign}}, source2[335:320]};
  wire [63:0]   extendResult_hi_lo_hi_hi_2 = {{16{source2[383] & sign}}, source2[383:368], {16{source2[367] & sign}}, source2[367:352]};
  wire [127:0]  extendResult_hi_lo_hi_2 = {extendResult_hi_lo_hi_hi_2, extendResult_hi_lo_hi_lo_2};
  wire [255:0]  extendResult_hi_lo_2 = {extendResult_hi_lo_hi_2, extendResult_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_lo_lo_2 = {{16{source2[415] & sign}}, source2[415:400], {16{source2[399] & sign}}, source2[399:384]};
  wire [63:0]   extendResult_hi_hi_lo_hi_2 = {{16{source2[447] & sign}}, source2[447:432], {16{source2[431] & sign}}, source2[431:416]};
  wire [127:0]  extendResult_hi_hi_lo_2 = {extendResult_hi_hi_lo_hi_2, extendResult_hi_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_hi_lo_2 = {{16{source2[479] & sign}}, source2[479:464], {16{source2[463] & sign}}, source2[463:448]};
  wire [63:0]   extendResult_hi_hi_hi_hi_2 = {{16{source2[511] & sign}}, source2[511:496], {16{source2[495] & sign}}, source2[495:480]};
  wire [127:0]  extendResult_hi_hi_hi_2 = {extendResult_hi_hi_hi_hi_2, extendResult_hi_hi_hi_lo_2};
  wire [255:0]  extendResult_hi_hi_2 = {extendResult_hi_hi_hi_2, extendResult_hi_hi_lo_2};
  wire [511:0]  extendResult_hi_2 = {extendResult_hi_hi_2, extendResult_hi_lo_2};
  wire [63:0]   extendResult_lo_lo_lo_lo_lo_2 = {{24{source2[15] & sign}}, source2[15:8], {24{source2[7] & sign}}, source2[7:0]};
  wire [63:0]   extendResult_lo_lo_lo_lo_hi_2 = {{24{source2[31] & sign}}, source2[31:24], {24{source2[23] & sign}}, source2[23:16]};
  wire [127:0]  extendResult_lo_lo_lo_lo_3 = {extendResult_lo_lo_lo_lo_hi_2, extendResult_lo_lo_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_lo_lo_hi_lo_2 = {{24{source2[47] & sign}}, source2[47:40], {24{source2[39] & sign}}, source2[39:32]};
  wire [63:0]   extendResult_lo_lo_lo_hi_hi_2 = {{24{source2[63] & sign}}, source2[63:56], {24{source2[55] & sign}}, source2[55:48]};
  wire [127:0]  extendResult_lo_lo_lo_hi_3 = {extendResult_lo_lo_lo_hi_hi_2, extendResult_lo_lo_lo_hi_lo_2};
  wire [255:0]  extendResult_lo_lo_lo_3 = {extendResult_lo_lo_lo_hi_3, extendResult_lo_lo_lo_lo_3};
  wire [63:0]   extendResult_lo_lo_hi_lo_lo_2 = {{24{source2[79] & sign}}, source2[79:72], {24{source2[71] & sign}}, source2[71:64]};
  wire [63:0]   extendResult_lo_lo_hi_lo_hi_2 = {{24{source2[95] & sign}}, source2[95:88], {24{source2[87] & sign}}, source2[87:80]};
  wire [127:0]  extendResult_lo_lo_hi_lo_3 = {extendResult_lo_lo_hi_lo_hi_2, extendResult_lo_lo_hi_lo_lo_2};
  wire [63:0]   extendResult_lo_lo_hi_hi_lo_2 = {{24{source2[111] & sign}}, source2[111:104], {24{source2[103] & sign}}, source2[103:96]};
  wire [63:0]   extendResult_lo_lo_hi_hi_hi_2 = {{24{source2[127] & sign}}, source2[127:120], {24{source2[119] & sign}}, source2[119:112]};
  wire [127:0]  extendResult_lo_lo_hi_hi_3 = {extendResult_lo_lo_hi_hi_hi_2, extendResult_lo_lo_hi_hi_lo_2};
  wire [255:0]  extendResult_lo_lo_hi_3 = {extendResult_lo_lo_hi_hi_3, extendResult_lo_lo_hi_lo_3};
  wire [511:0]  extendResult_lo_lo_3 = {extendResult_lo_lo_hi_3, extendResult_lo_lo_lo_3};
  wire [63:0]   extendResult_lo_hi_lo_lo_lo_2 = {{24{source2[143] & sign}}, source2[143:136], {24{source2[135] & sign}}, source2[135:128]};
  wire [63:0]   extendResult_lo_hi_lo_lo_hi_2 = {{24{source2[159] & sign}}, source2[159:152], {24{source2[151] & sign}}, source2[151:144]};
  wire [127:0]  extendResult_lo_hi_lo_lo_3 = {extendResult_lo_hi_lo_lo_hi_2, extendResult_lo_hi_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_lo_hi_lo_2 = {{24{source2[175] & sign}}, source2[175:168], {24{source2[167] & sign}}, source2[167:160]};
  wire [63:0]   extendResult_lo_hi_lo_hi_hi_2 = {{24{source2[191] & sign}}, source2[191:184], {24{source2[183] & sign}}, source2[183:176]};
  wire [127:0]  extendResult_lo_hi_lo_hi_3 = {extendResult_lo_hi_lo_hi_hi_2, extendResult_lo_hi_lo_hi_lo_2};
  wire [255:0]  extendResult_lo_hi_lo_3 = {extendResult_lo_hi_lo_hi_3, extendResult_lo_hi_lo_lo_3};
  wire [63:0]   extendResult_lo_hi_hi_lo_lo_2 = {{24{source2[207] & sign}}, source2[207:200], {24{source2[199] & sign}}, source2[199:192]};
  wire [63:0]   extendResult_lo_hi_hi_lo_hi_2 = {{24{source2[223] & sign}}, source2[223:216], {24{source2[215] & sign}}, source2[215:208]};
  wire [127:0]  extendResult_lo_hi_hi_lo_3 = {extendResult_lo_hi_hi_lo_hi_2, extendResult_lo_hi_hi_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_hi_hi_lo_2 = {{24{source2[239] & sign}}, source2[239:232], {24{source2[231] & sign}}, source2[231:224]};
  wire [63:0]   extendResult_lo_hi_hi_hi_hi_2 = {{24{source2[255] & sign}}, source2[255:248], {24{source2[247] & sign}}, source2[247:240]};
  wire [127:0]  extendResult_lo_hi_hi_hi_3 = {extendResult_lo_hi_hi_hi_hi_2, extendResult_lo_hi_hi_hi_lo_2};
  wire [255:0]  extendResult_lo_hi_hi_3 = {extendResult_lo_hi_hi_hi_3, extendResult_lo_hi_hi_lo_3};
  wire [511:0]  extendResult_lo_hi_3 = {extendResult_lo_hi_hi_3, extendResult_lo_hi_lo_3};
  wire [1023:0] extendResult_lo_3 = {extendResult_lo_hi_3, extendResult_lo_lo_3};
  wire [63:0]   extendResult_hi_lo_lo_lo_lo_2 = {{24{source2[271] & sign}}, source2[271:264], {24{source2[263] & sign}}, source2[263:256]};
  wire [63:0]   extendResult_hi_lo_lo_lo_hi_2 = {{24{source2[287] & sign}}, source2[287:280], {24{source2[279] & sign}}, source2[279:272]};
  wire [127:0]  extendResult_hi_lo_lo_lo_3 = {extendResult_hi_lo_lo_lo_hi_2, extendResult_hi_lo_lo_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_lo_hi_lo_2 = {{24{source2[303] & sign}}, source2[303:296], {24{source2[295] & sign}}, source2[295:288]};
  wire [63:0]   extendResult_hi_lo_lo_hi_hi_2 = {{24{source2[319] & sign}}, source2[319:312], {24{source2[311] & sign}}, source2[311:304]};
  wire [127:0]  extendResult_hi_lo_lo_hi_3 = {extendResult_hi_lo_lo_hi_hi_2, extendResult_hi_lo_lo_hi_lo_2};
  wire [255:0]  extendResult_hi_lo_lo_3 = {extendResult_hi_lo_lo_hi_3, extendResult_hi_lo_lo_lo_3};
  wire [63:0]   extendResult_hi_lo_hi_lo_lo_2 = {{24{source2[335] & sign}}, source2[335:328], {24{source2[327] & sign}}, source2[327:320]};
  wire [63:0]   extendResult_hi_lo_hi_lo_hi_2 = {{24{source2[351] & sign}}, source2[351:344], {24{source2[343] & sign}}, source2[343:336]};
  wire [127:0]  extendResult_hi_lo_hi_lo_3 = {extendResult_hi_lo_hi_lo_hi_2, extendResult_hi_lo_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_hi_hi_lo_2 = {{24{source2[367] & sign}}, source2[367:360], {24{source2[359] & sign}}, source2[359:352]};
  wire [63:0]   extendResult_hi_lo_hi_hi_hi_2 = {{24{source2[383] & sign}}, source2[383:376], {24{source2[375] & sign}}, source2[375:368]};
  wire [127:0]  extendResult_hi_lo_hi_hi_3 = {extendResult_hi_lo_hi_hi_hi_2, extendResult_hi_lo_hi_hi_lo_2};
  wire [255:0]  extendResult_hi_lo_hi_3 = {extendResult_hi_lo_hi_hi_3, extendResult_hi_lo_hi_lo_3};
  wire [511:0]  extendResult_hi_lo_3 = {extendResult_hi_lo_hi_3, extendResult_hi_lo_lo_3};
  wire [63:0]   extendResult_hi_hi_lo_lo_lo_2 = {{24{source2[399] & sign}}, source2[399:392], {24{source2[391] & sign}}, source2[391:384]};
  wire [63:0]   extendResult_hi_hi_lo_lo_hi_2 = {{24{source2[415] & sign}}, source2[415:408], {24{source2[407] & sign}}, source2[407:400]};
  wire [127:0]  extendResult_hi_hi_lo_lo_3 = {extendResult_hi_hi_lo_lo_hi_2, extendResult_hi_hi_lo_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_lo_hi_lo_2 = {{24{source2[431] & sign}}, source2[431:424], {24{source2[423] & sign}}, source2[423:416]};
  wire [63:0]   extendResult_hi_hi_lo_hi_hi_2 = {{24{source2[447] & sign}}, source2[447:440], {24{source2[439] & sign}}, source2[439:432]};
  wire [127:0]  extendResult_hi_hi_lo_hi_3 = {extendResult_hi_hi_lo_hi_hi_2, extendResult_hi_hi_lo_hi_lo_2};
  wire [255:0]  extendResult_hi_hi_lo_3 = {extendResult_hi_hi_lo_hi_3, extendResult_hi_hi_lo_lo_3};
  wire [63:0]   extendResult_hi_hi_hi_lo_lo_2 = {{24{source2[463] & sign}}, source2[463:456], {24{source2[455] & sign}}, source2[455:448]};
  wire [63:0]   extendResult_hi_hi_hi_lo_hi_2 = {{24{source2[479] & sign}}, source2[479:472], {24{source2[471] & sign}}, source2[471:464]};
  wire [127:0]  extendResult_hi_hi_hi_lo_3 = {extendResult_hi_hi_hi_lo_hi_2, extendResult_hi_hi_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_hi_hi_lo_2 = {{24{source2[495] & sign}}, source2[495:488], {24{source2[487] & sign}}, source2[487:480]};
  wire [63:0]   extendResult_hi_hi_hi_hi_hi_2 = {{24{source2[511] & sign}}, source2[511:504], {24{source2[503] & sign}}, source2[503:496]};
  wire [127:0]  extendResult_hi_hi_hi_hi_3 = {extendResult_hi_hi_hi_hi_hi_2, extendResult_hi_hi_hi_hi_lo_2};
  wire [255:0]  extendResult_hi_hi_hi_3 = {extendResult_hi_hi_hi_hi_3, extendResult_hi_hi_hi_lo_3};
  wire [511:0]  extendResult_hi_hi_3 = {extendResult_hi_hi_hi_3, extendResult_hi_hi_lo_3};
  wire [1023:0] extendResult_hi_3 = {extendResult_hi_hi_3, extendResult_hi_lo_3};
  wire [2047:0] extendResult =
    (eew1H[1] ? {1024'h0, _extendResult_T_969[0] ? {extendResult_hi, extendResult_lo} : 1024'h0} | (_extendResult_T_969[1] ? {extendResult_hi_1, extendResult_lo_1} : 2048'h0) : 2048'h0)
    | (eew1H[2] ? {1024'h0, _extendResult_T_969[0] ? {extendResult_hi_2, extendResult_lo_2} : 1024'h0} | (_extendResult_T_969[1] ? {extendResult_hi_3, extendResult_lo_3} : 2048'h0) : 2048'h0);
  assign out = isMaskDestination ? maskDestinationResult : extendResult[1023:0];
endmodule

