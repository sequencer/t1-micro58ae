module MaskExtend(
  input  [1:0]   in_eew,
  input  [2:0]   in_uop,
  input  [511:0] in_source2,
  input  [4:0]   in_groupCounter,
  output [511:0] out
);

  wire [3:0]    _eew1H_T = 4'h1 << in_eew;
  wire [2:0]    eew1H = _eew1H_T[2:0];
  wire          isMaskDestination = in_uop == 3'h0;
  wire [31:0]   sourceDataVec_0 = in_source2[31:0];
  wire [31:0]   sourceDataVec_1 = in_source2[63:32];
  wire [31:0]   sourceDataVec_2 = in_source2[95:64];
  wire [31:0]   sourceDataVec_3 = in_source2[127:96];
  wire [31:0]   sourceDataVec_4 = in_source2[159:128];
  wire [31:0]   sourceDataVec_5 = in_source2[191:160];
  wire [31:0]   sourceDataVec_6 = in_source2[223:192];
  wire [31:0]   sourceDataVec_7 = in_source2[255:224];
  wire [31:0]   sourceDataVec_8 = in_source2[287:256];
  wire [31:0]   sourceDataVec_9 = in_source2[319:288];
  wire [31:0]   sourceDataVec_10 = in_source2[351:320];
  wire [31:0]   sourceDataVec_11 = in_source2[383:352];
  wire [31:0]   sourceDataVec_12 = in_source2[415:384];
  wire [31:0]   sourceDataVec_13 = in_source2[447:416];
  wire [31:0]   sourceDataVec_14 = in_source2[479:448];
  wire [31:0]   sourceDataVec_15 = in_source2[511:480];
  wire [1:0]    maskDestinationResult_lo = sourceDataVec_0[1:0];
  wire [1:0]    maskDestinationResult_hi = sourceDataVec_0[3:2];
  wire [1:0]    maskDestinationResult_lo_1 = sourceDataVec_0[5:4];
  wire [1:0]    maskDestinationResult_hi_1 = sourceDataVec_0[7:6];
  wire [1:0]    maskDestinationResult_lo_2 = sourceDataVec_0[9:8];
  wire [1:0]    maskDestinationResult_hi_2 = sourceDataVec_0[11:10];
  wire [1:0]    maskDestinationResult_lo_3 = sourceDataVec_0[13:12];
  wire [1:0]    maskDestinationResult_hi_3 = sourceDataVec_0[15:14];
  wire [1:0]    maskDestinationResult_lo_4 = sourceDataVec_0[17:16];
  wire [1:0]    maskDestinationResult_hi_4 = sourceDataVec_0[19:18];
  wire [1:0]    maskDestinationResult_lo_5 = sourceDataVec_0[21:20];
  wire [1:0]    maskDestinationResult_hi_5 = sourceDataVec_0[23:22];
  wire [1:0]    maskDestinationResult_lo_6 = sourceDataVec_0[25:24];
  wire [1:0]    maskDestinationResult_hi_6 = sourceDataVec_0[27:26];
  wire [1:0]    maskDestinationResult_lo_7 = sourceDataVec_0[29:28];
  wire [1:0]    maskDestinationResult_hi_7 = sourceDataVec_0[31:30];
  wire [1:0]    maskDestinationResult_lo_8 = sourceDataVec_1[1:0];
  wire [1:0]    maskDestinationResult_hi_8 = sourceDataVec_1[3:2];
  wire [1:0]    maskDestinationResult_lo_9 = sourceDataVec_1[5:4];
  wire [1:0]    maskDestinationResult_hi_9 = sourceDataVec_1[7:6];
  wire [1:0]    maskDestinationResult_lo_10 = sourceDataVec_1[9:8];
  wire [1:0]    maskDestinationResult_hi_10 = sourceDataVec_1[11:10];
  wire [1:0]    maskDestinationResult_lo_11 = sourceDataVec_1[13:12];
  wire [1:0]    maskDestinationResult_hi_11 = sourceDataVec_1[15:14];
  wire [1:0]    maskDestinationResult_lo_12 = sourceDataVec_1[17:16];
  wire [1:0]    maskDestinationResult_hi_12 = sourceDataVec_1[19:18];
  wire [1:0]    maskDestinationResult_lo_13 = sourceDataVec_1[21:20];
  wire [1:0]    maskDestinationResult_hi_13 = sourceDataVec_1[23:22];
  wire [1:0]    maskDestinationResult_lo_14 = sourceDataVec_1[25:24];
  wire [1:0]    maskDestinationResult_hi_14 = sourceDataVec_1[27:26];
  wire [1:0]    maskDestinationResult_lo_15 = sourceDataVec_1[29:28];
  wire [1:0]    maskDestinationResult_hi_15 = sourceDataVec_1[31:30];
  wire [1:0]    maskDestinationResult_lo_16 = sourceDataVec_2[1:0];
  wire [1:0]    maskDestinationResult_hi_16 = sourceDataVec_2[3:2];
  wire [1:0]    maskDestinationResult_lo_17 = sourceDataVec_2[5:4];
  wire [1:0]    maskDestinationResult_hi_17 = sourceDataVec_2[7:6];
  wire [1:0]    maskDestinationResult_lo_18 = sourceDataVec_2[9:8];
  wire [1:0]    maskDestinationResult_hi_18 = sourceDataVec_2[11:10];
  wire [1:0]    maskDestinationResult_lo_19 = sourceDataVec_2[13:12];
  wire [1:0]    maskDestinationResult_hi_19 = sourceDataVec_2[15:14];
  wire [1:0]    maskDestinationResult_lo_20 = sourceDataVec_2[17:16];
  wire [1:0]    maskDestinationResult_hi_20 = sourceDataVec_2[19:18];
  wire [1:0]    maskDestinationResult_lo_21 = sourceDataVec_2[21:20];
  wire [1:0]    maskDestinationResult_hi_21 = sourceDataVec_2[23:22];
  wire [1:0]    maskDestinationResult_lo_22 = sourceDataVec_2[25:24];
  wire [1:0]    maskDestinationResult_hi_22 = sourceDataVec_2[27:26];
  wire [1:0]    maskDestinationResult_lo_23 = sourceDataVec_2[29:28];
  wire [1:0]    maskDestinationResult_hi_23 = sourceDataVec_2[31:30];
  wire [1:0]    maskDestinationResult_lo_24 = sourceDataVec_3[1:0];
  wire [1:0]    maskDestinationResult_hi_24 = sourceDataVec_3[3:2];
  wire [1:0]    maskDestinationResult_lo_25 = sourceDataVec_3[5:4];
  wire [1:0]    maskDestinationResult_hi_25 = sourceDataVec_3[7:6];
  wire [1:0]    maskDestinationResult_lo_26 = sourceDataVec_3[9:8];
  wire [1:0]    maskDestinationResult_hi_26 = sourceDataVec_3[11:10];
  wire [1:0]    maskDestinationResult_lo_27 = sourceDataVec_3[13:12];
  wire [1:0]    maskDestinationResult_hi_27 = sourceDataVec_3[15:14];
  wire [1:0]    maskDestinationResult_lo_28 = sourceDataVec_3[17:16];
  wire [1:0]    maskDestinationResult_hi_28 = sourceDataVec_3[19:18];
  wire [1:0]    maskDestinationResult_lo_29 = sourceDataVec_3[21:20];
  wire [1:0]    maskDestinationResult_hi_29 = sourceDataVec_3[23:22];
  wire [1:0]    maskDestinationResult_lo_30 = sourceDataVec_3[25:24];
  wire [1:0]    maskDestinationResult_hi_30 = sourceDataVec_3[27:26];
  wire [1:0]    maskDestinationResult_lo_31 = sourceDataVec_3[29:28];
  wire [1:0]    maskDestinationResult_hi_31 = sourceDataVec_3[31:30];
  wire [1:0]    maskDestinationResult_lo_32 = sourceDataVec_4[1:0];
  wire [1:0]    maskDestinationResult_hi_32 = sourceDataVec_4[3:2];
  wire [1:0]    maskDestinationResult_lo_33 = sourceDataVec_4[5:4];
  wire [1:0]    maskDestinationResult_hi_33 = sourceDataVec_4[7:6];
  wire [1:0]    maskDestinationResult_lo_34 = sourceDataVec_4[9:8];
  wire [1:0]    maskDestinationResult_hi_34 = sourceDataVec_4[11:10];
  wire [1:0]    maskDestinationResult_lo_35 = sourceDataVec_4[13:12];
  wire [1:0]    maskDestinationResult_hi_35 = sourceDataVec_4[15:14];
  wire [1:0]    maskDestinationResult_lo_36 = sourceDataVec_4[17:16];
  wire [1:0]    maskDestinationResult_hi_36 = sourceDataVec_4[19:18];
  wire [1:0]    maskDestinationResult_lo_37 = sourceDataVec_4[21:20];
  wire [1:0]    maskDestinationResult_hi_37 = sourceDataVec_4[23:22];
  wire [1:0]    maskDestinationResult_lo_38 = sourceDataVec_4[25:24];
  wire [1:0]    maskDestinationResult_hi_38 = sourceDataVec_4[27:26];
  wire [1:0]    maskDestinationResult_lo_39 = sourceDataVec_4[29:28];
  wire [1:0]    maskDestinationResult_hi_39 = sourceDataVec_4[31:30];
  wire [1:0]    maskDestinationResult_lo_40 = sourceDataVec_5[1:0];
  wire [1:0]    maskDestinationResult_hi_40 = sourceDataVec_5[3:2];
  wire [1:0]    maskDestinationResult_lo_41 = sourceDataVec_5[5:4];
  wire [1:0]    maskDestinationResult_hi_41 = sourceDataVec_5[7:6];
  wire [1:0]    maskDestinationResult_lo_42 = sourceDataVec_5[9:8];
  wire [1:0]    maskDestinationResult_hi_42 = sourceDataVec_5[11:10];
  wire [1:0]    maskDestinationResult_lo_43 = sourceDataVec_5[13:12];
  wire [1:0]    maskDestinationResult_hi_43 = sourceDataVec_5[15:14];
  wire [1:0]    maskDestinationResult_lo_44 = sourceDataVec_5[17:16];
  wire [1:0]    maskDestinationResult_hi_44 = sourceDataVec_5[19:18];
  wire [1:0]    maskDestinationResult_lo_45 = sourceDataVec_5[21:20];
  wire [1:0]    maskDestinationResult_hi_45 = sourceDataVec_5[23:22];
  wire [1:0]    maskDestinationResult_lo_46 = sourceDataVec_5[25:24];
  wire [1:0]    maskDestinationResult_hi_46 = sourceDataVec_5[27:26];
  wire [1:0]    maskDestinationResult_lo_47 = sourceDataVec_5[29:28];
  wire [1:0]    maskDestinationResult_hi_47 = sourceDataVec_5[31:30];
  wire [1:0]    maskDestinationResult_lo_48 = sourceDataVec_6[1:0];
  wire [1:0]    maskDestinationResult_hi_48 = sourceDataVec_6[3:2];
  wire [1:0]    maskDestinationResult_lo_49 = sourceDataVec_6[5:4];
  wire [1:0]    maskDestinationResult_hi_49 = sourceDataVec_6[7:6];
  wire [1:0]    maskDestinationResult_lo_50 = sourceDataVec_6[9:8];
  wire [1:0]    maskDestinationResult_hi_50 = sourceDataVec_6[11:10];
  wire [1:0]    maskDestinationResult_lo_51 = sourceDataVec_6[13:12];
  wire [1:0]    maskDestinationResult_hi_51 = sourceDataVec_6[15:14];
  wire [1:0]    maskDestinationResult_lo_52 = sourceDataVec_6[17:16];
  wire [1:0]    maskDestinationResult_hi_52 = sourceDataVec_6[19:18];
  wire [1:0]    maskDestinationResult_lo_53 = sourceDataVec_6[21:20];
  wire [1:0]    maskDestinationResult_hi_53 = sourceDataVec_6[23:22];
  wire [1:0]    maskDestinationResult_lo_54 = sourceDataVec_6[25:24];
  wire [1:0]    maskDestinationResult_hi_54 = sourceDataVec_6[27:26];
  wire [1:0]    maskDestinationResult_lo_55 = sourceDataVec_6[29:28];
  wire [1:0]    maskDestinationResult_hi_55 = sourceDataVec_6[31:30];
  wire [1:0]    maskDestinationResult_lo_56 = sourceDataVec_7[1:0];
  wire [1:0]    maskDestinationResult_hi_56 = sourceDataVec_7[3:2];
  wire [1:0]    maskDestinationResult_lo_57 = sourceDataVec_7[5:4];
  wire [1:0]    maskDestinationResult_hi_57 = sourceDataVec_7[7:6];
  wire [1:0]    maskDestinationResult_lo_58 = sourceDataVec_7[9:8];
  wire [1:0]    maskDestinationResult_hi_58 = sourceDataVec_7[11:10];
  wire [1:0]    maskDestinationResult_lo_59 = sourceDataVec_7[13:12];
  wire [1:0]    maskDestinationResult_hi_59 = sourceDataVec_7[15:14];
  wire [1:0]    maskDestinationResult_lo_60 = sourceDataVec_7[17:16];
  wire [1:0]    maskDestinationResult_hi_60 = sourceDataVec_7[19:18];
  wire [1:0]    maskDestinationResult_lo_61 = sourceDataVec_7[21:20];
  wire [1:0]    maskDestinationResult_hi_61 = sourceDataVec_7[23:22];
  wire [1:0]    maskDestinationResult_lo_62 = sourceDataVec_7[25:24];
  wire [1:0]    maskDestinationResult_hi_62 = sourceDataVec_7[27:26];
  wire [1:0]    maskDestinationResult_lo_63 = sourceDataVec_7[29:28];
  wire [1:0]    maskDestinationResult_hi_63 = sourceDataVec_7[31:30];
  wire [1:0]    maskDestinationResult_lo_64 = sourceDataVec_8[1:0];
  wire [1:0]    maskDestinationResult_hi_64 = sourceDataVec_8[3:2];
  wire [1:0]    maskDestinationResult_lo_65 = sourceDataVec_8[5:4];
  wire [1:0]    maskDestinationResult_hi_65 = sourceDataVec_8[7:6];
  wire [1:0]    maskDestinationResult_lo_66 = sourceDataVec_8[9:8];
  wire [1:0]    maskDestinationResult_hi_66 = sourceDataVec_8[11:10];
  wire [1:0]    maskDestinationResult_lo_67 = sourceDataVec_8[13:12];
  wire [1:0]    maskDestinationResult_hi_67 = sourceDataVec_8[15:14];
  wire [1:0]    maskDestinationResult_lo_68 = sourceDataVec_8[17:16];
  wire [1:0]    maskDestinationResult_hi_68 = sourceDataVec_8[19:18];
  wire [1:0]    maskDestinationResult_lo_69 = sourceDataVec_8[21:20];
  wire [1:0]    maskDestinationResult_hi_69 = sourceDataVec_8[23:22];
  wire [1:0]    maskDestinationResult_lo_70 = sourceDataVec_8[25:24];
  wire [1:0]    maskDestinationResult_hi_70 = sourceDataVec_8[27:26];
  wire [1:0]    maskDestinationResult_lo_71 = sourceDataVec_8[29:28];
  wire [1:0]    maskDestinationResult_hi_71 = sourceDataVec_8[31:30];
  wire [1:0]    maskDestinationResult_lo_72 = sourceDataVec_9[1:0];
  wire [1:0]    maskDestinationResult_hi_72 = sourceDataVec_9[3:2];
  wire [1:0]    maskDestinationResult_lo_73 = sourceDataVec_9[5:4];
  wire [1:0]    maskDestinationResult_hi_73 = sourceDataVec_9[7:6];
  wire [1:0]    maskDestinationResult_lo_74 = sourceDataVec_9[9:8];
  wire [1:0]    maskDestinationResult_hi_74 = sourceDataVec_9[11:10];
  wire [1:0]    maskDestinationResult_lo_75 = sourceDataVec_9[13:12];
  wire [1:0]    maskDestinationResult_hi_75 = sourceDataVec_9[15:14];
  wire [1:0]    maskDestinationResult_lo_76 = sourceDataVec_9[17:16];
  wire [1:0]    maskDestinationResult_hi_76 = sourceDataVec_9[19:18];
  wire [1:0]    maskDestinationResult_lo_77 = sourceDataVec_9[21:20];
  wire [1:0]    maskDestinationResult_hi_77 = sourceDataVec_9[23:22];
  wire [1:0]    maskDestinationResult_lo_78 = sourceDataVec_9[25:24];
  wire [1:0]    maskDestinationResult_hi_78 = sourceDataVec_9[27:26];
  wire [1:0]    maskDestinationResult_lo_79 = sourceDataVec_9[29:28];
  wire [1:0]    maskDestinationResult_hi_79 = sourceDataVec_9[31:30];
  wire [1:0]    maskDestinationResult_lo_80 = sourceDataVec_10[1:0];
  wire [1:0]    maskDestinationResult_hi_80 = sourceDataVec_10[3:2];
  wire [1:0]    maskDestinationResult_lo_81 = sourceDataVec_10[5:4];
  wire [1:0]    maskDestinationResult_hi_81 = sourceDataVec_10[7:6];
  wire [1:0]    maskDestinationResult_lo_82 = sourceDataVec_10[9:8];
  wire [1:0]    maskDestinationResult_hi_82 = sourceDataVec_10[11:10];
  wire [1:0]    maskDestinationResult_lo_83 = sourceDataVec_10[13:12];
  wire [1:0]    maskDestinationResult_hi_83 = sourceDataVec_10[15:14];
  wire [1:0]    maskDestinationResult_lo_84 = sourceDataVec_10[17:16];
  wire [1:0]    maskDestinationResult_hi_84 = sourceDataVec_10[19:18];
  wire [1:0]    maskDestinationResult_lo_85 = sourceDataVec_10[21:20];
  wire [1:0]    maskDestinationResult_hi_85 = sourceDataVec_10[23:22];
  wire [1:0]    maskDestinationResult_lo_86 = sourceDataVec_10[25:24];
  wire [1:0]    maskDestinationResult_hi_86 = sourceDataVec_10[27:26];
  wire [1:0]    maskDestinationResult_lo_87 = sourceDataVec_10[29:28];
  wire [1:0]    maskDestinationResult_hi_87 = sourceDataVec_10[31:30];
  wire [1:0]    maskDestinationResult_lo_88 = sourceDataVec_11[1:0];
  wire [1:0]    maskDestinationResult_hi_88 = sourceDataVec_11[3:2];
  wire [1:0]    maskDestinationResult_lo_89 = sourceDataVec_11[5:4];
  wire [1:0]    maskDestinationResult_hi_89 = sourceDataVec_11[7:6];
  wire [1:0]    maskDestinationResult_lo_90 = sourceDataVec_11[9:8];
  wire [1:0]    maskDestinationResult_hi_90 = sourceDataVec_11[11:10];
  wire [1:0]    maskDestinationResult_lo_91 = sourceDataVec_11[13:12];
  wire [1:0]    maskDestinationResult_hi_91 = sourceDataVec_11[15:14];
  wire [1:0]    maskDestinationResult_lo_92 = sourceDataVec_11[17:16];
  wire [1:0]    maskDestinationResult_hi_92 = sourceDataVec_11[19:18];
  wire [1:0]    maskDestinationResult_lo_93 = sourceDataVec_11[21:20];
  wire [1:0]    maskDestinationResult_hi_93 = sourceDataVec_11[23:22];
  wire [1:0]    maskDestinationResult_lo_94 = sourceDataVec_11[25:24];
  wire [1:0]    maskDestinationResult_hi_94 = sourceDataVec_11[27:26];
  wire [1:0]    maskDestinationResult_lo_95 = sourceDataVec_11[29:28];
  wire [1:0]    maskDestinationResult_hi_95 = sourceDataVec_11[31:30];
  wire [1:0]    maskDestinationResult_lo_96 = sourceDataVec_12[1:0];
  wire [1:0]    maskDestinationResult_hi_96 = sourceDataVec_12[3:2];
  wire [1:0]    maskDestinationResult_lo_97 = sourceDataVec_12[5:4];
  wire [1:0]    maskDestinationResult_hi_97 = sourceDataVec_12[7:6];
  wire [1:0]    maskDestinationResult_lo_98 = sourceDataVec_12[9:8];
  wire [1:0]    maskDestinationResult_hi_98 = sourceDataVec_12[11:10];
  wire [1:0]    maskDestinationResult_lo_99 = sourceDataVec_12[13:12];
  wire [1:0]    maskDestinationResult_hi_99 = sourceDataVec_12[15:14];
  wire [1:0]    maskDestinationResult_lo_100 = sourceDataVec_12[17:16];
  wire [1:0]    maskDestinationResult_hi_100 = sourceDataVec_12[19:18];
  wire [1:0]    maskDestinationResult_lo_101 = sourceDataVec_12[21:20];
  wire [1:0]    maskDestinationResult_hi_101 = sourceDataVec_12[23:22];
  wire [1:0]    maskDestinationResult_lo_102 = sourceDataVec_12[25:24];
  wire [1:0]    maskDestinationResult_hi_102 = sourceDataVec_12[27:26];
  wire [1:0]    maskDestinationResult_lo_103 = sourceDataVec_12[29:28];
  wire [1:0]    maskDestinationResult_hi_103 = sourceDataVec_12[31:30];
  wire [1:0]    maskDestinationResult_lo_104 = sourceDataVec_13[1:0];
  wire [1:0]    maskDestinationResult_hi_104 = sourceDataVec_13[3:2];
  wire [1:0]    maskDestinationResult_lo_105 = sourceDataVec_13[5:4];
  wire [1:0]    maskDestinationResult_hi_105 = sourceDataVec_13[7:6];
  wire [1:0]    maskDestinationResult_lo_106 = sourceDataVec_13[9:8];
  wire [1:0]    maskDestinationResult_hi_106 = sourceDataVec_13[11:10];
  wire [1:0]    maskDestinationResult_lo_107 = sourceDataVec_13[13:12];
  wire [1:0]    maskDestinationResult_hi_107 = sourceDataVec_13[15:14];
  wire [1:0]    maskDestinationResult_lo_108 = sourceDataVec_13[17:16];
  wire [1:0]    maskDestinationResult_hi_108 = sourceDataVec_13[19:18];
  wire [1:0]    maskDestinationResult_lo_109 = sourceDataVec_13[21:20];
  wire [1:0]    maskDestinationResult_hi_109 = sourceDataVec_13[23:22];
  wire [1:0]    maskDestinationResult_lo_110 = sourceDataVec_13[25:24];
  wire [1:0]    maskDestinationResult_hi_110 = sourceDataVec_13[27:26];
  wire [1:0]    maskDestinationResult_lo_111 = sourceDataVec_13[29:28];
  wire [1:0]    maskDestinationResult_hi_111 = sourceDataVec_13[31:30];
  wire [1:0]    maskDestinationResult_lo_112 = sourceDataVec_14[1:0];
  wire [1:0]    maskDestinationResult_hi_112 = sourceDataVec_14[3:2];
  wire [1:0]    maskDestinationResult_lo_113 = sourceDataVec_14[5:4];
  wire [1:0]    maskDestinationResult_hi_113 = sourceDataVec_14[7:6];
  wire [1:0]    maskDestinationResult_lo_114 = sourceDataVec_14[9:8];
  wire [1:0]    maskDestinationResult_hi_114 = sourceDataVec_14[11:10];
  wire [1:0]    maskDestinationResult_lo_115 = sourceDataVec_14[13:12];
  wire [1:0]    maskDestinationResult_hi_115 = sourceDataVec_14[15:14];
  wire [1:0]    maskDestinationResult_lo_116 = sourceDataVec_14[17:16];
  wire [1:0]    maskDestinationResult_hi_116 = sourceDataVec_14[19:18];
  wire [1:0]    maskDestinationResult_lo_117 = sourceDataVec_14[21:20];
  wire [1:0]    maskDestinationResult_hi_117 = sourceDataVec_14[23:22];
  wire [1:0]    maskDestinationResult_lo_118 = sourceDataVec_14[25:24];
  wire [1:0]    maskDestinationResult_hi_118 = sourceDataVec_14[27:26];
  wire [1:0]    maskDestinationResult_lo_119 = sourceDataVec_14[29:28];
  wire [1:0]    maskDestinationResult_hi_119 = sourceDataVec_14[31:30];
  wire [1:0]    maskDestinationResult_lo_120 = sourceDataVec_15[1:0];
  wire [1:0]    maskDestinationResult_hi_120 = sourceDataVec_15[3:2];
  wire [1:0]    maskDestinationResult_lo_121 = sourceDataVec_15[5:4];
  wire [1:0]    maskDestinationResult_hi_121 = sourceDataVec_15[7:6];
  wire [1:0]    maskDestinationResult_lo_122 = sourceDataVec_15[9:8];
  wire [1:0]    maskDestinationResult_hi_122 = sourceDataVec_15[11:10];
  wire [1:0]    maskDestinationResult_lo_123 = sourceDataVec_15[13:12];
  wire [1:0]    maskDestinationResult_hi_123 = sourceDataVec_15[15:14];
  wire [1:0]    maskDestinationResult_lo_124 = sourceDataVec_15[17:16];
  wire [1:0]    maskDestinationResult_hi_124 = sourceDataVec_15[19:18];
  wire [1:0]    maskDestinationResult_lo_125 = sourceDataVec_15[21:20];
  wire [1:0]    maskDestinationResult_hi_125 = sourceDataVec_15[23:22];
  wire [1:0]    maskDestinationResult_lo_126 = sourceDataVec_15[25:24];
  wire [1:0]    maskDestinationResult_hi_126 = sourceDataVec_15[27:26];
  wire [1:0]    maskDestinationResult_lo_127 = sourceDataVec_15[29:28];
  wire [1:0]    maskDestinationResult_hi_127 = sourceDataVec_15[31:30];
  wire [7:0]    maskDestinationResult_lo_lo_lo = {maskDestinationResult_hi_8, maskDestinationResult_lo_8, maskDestinationResult_hi, maskDestinationResult_lo};
  wire [7:0]    maskDestinationResult_lo_lo_hi = {maskDestinationResult_hi_24, maskDestinationResult_lo_24, maskDestinationResult_hi_16, maskDestinationResult_lo_16};
  wire [15:0]   maskDestinationResult_lo_lo = {maskDestinationResult_lo_lo_hi, maskDestinationResult_lo_lo_lo};
  wire [7:0]    maskDestinationResult_lo_hi_lo = {maskDestinationResult_hi_40, maskDestinationResult_lo_40, maskDestinationResult_hi_32, maskDestinationResult_lo_32};
  wire [7:0]    maskDestinationResult_lo_hi_hi = {maskDestinationResult_hi_56, maskDestinationResult_lo_56, maskDestinationResult_hi_48, maskDestinationResult_lo_48};
  wire [15:0]   maskDestinationResult_lo_hi = {maskDestinationResult_lo_hi_hi, maskDestinationResult_lo_hi_lo};
  wire [31:0]   maskDestinationResult_lo_128 = {maskDestinationResult_lo_hi, maskDestinationResult_lo_lo};
  wire [7:0]    maskDestinationResult_hi_lo_lo = {maskDestinationResult_hi_72, maskDestinationResult_lo_72, maskDestinationResult_hi_64, maskDestinationResult_lo_64};
  wire [7:0]    maskDestinationResult_hi_lo_hi = {maskDestinationResult_hi_88, maskDestinationResult_lo_88, maskDestinationResult_hi_80, maskDestinationResult_lo_80};
  wire [15:0]   maskDestinationResult_hi_lo = {maskDestinationResult_hi_lo_hi, maskDestinationResult_hi_lo_lo};
  wire [7:0]    maskDestinationResult_hi_hi_lo = {maskDestinationResult_hi_104, maskDestinationResult_lo_104, maskDestinationResult_hi_96, maskDestinationResult_lo_96};
  wire [7:0]    maskDestinationResult_hi_hi_hi = {maskDestinationResult_hi_120, maskDestinationResult_lo_120, maskDestinationResult_hi_112, maskDestinationResult_lo_112};
  wire [15:0]   maskDestinationResult_hi_hi = {maskDestinationResult_hi_hi_hi, maskDestinationResult_hi_hi_lo};
  wire [31:0]   maskDestinationResult_hi_128 = {maskDestinationResult_hi_hi, maskDestinationResult_hi_lo};
  wire [7:0]    maskDestinationResult_lo_lo_lo_1 = {maskDestinationResult_hi_9, maskDestinationResult_lo_9, maskDestinationResult_hi_1, maskDestinationResult_lo_1};
  wire [7:0]    maskDestinationResult_lo_lo_hi_1 = {maskDestinationResult_hi_25, maskDestinationResult_lo_25, maskDestinationResult_hi_17, maskDestinationResult_lo_17};
  wire [15:0]   maskDestinationResult_lo_lo_1 = {maskDestinationResult_lo_lo_hi_1, maskDestinationResult_lo_lo_lo_1};
  wire [7:0]    maskDestinationResult_lo_hi_lo_1 = {maskDestinationResult_hi_41, maskDestinationResult_lo_41, maskDestinationResult_hi_33, maskDestinationResult_lo_33};
  wire [7:0]    maskDestinationResult_lo_hi_hi_1 = {maskDestinationResult_hi_57, maskDestinationResult_lo_57, maskDestinationResult_hi_49, maskDestinationResult_lo_49};
  wire [15:0]   maskDestinationResult_lo_hi_1 = {maskDestinationResult_lo_hi_hi_1, maskDestinationResult_lo_hi_lo_1};
  wire [31:0]   maskDestinationResult_lo_129 = {maskDestinationResult_lo_hi_1, maskDestinationResult_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_lo_lo_1 = {maskDestinationResult_hi_73, maskDestinationResult_lo_73, maskDestinationResult_hi_65, maskDestinationResult_lo_65};
  wire [7:0]    maskDestinationResult_hi_lo_hi_1 = {maskDestinationResult_hi_89, maskDestinationResult_lo_89, maskDestinationResult_hi_81, maskDestinationResult_lo_81};
  wire [15:0]   maskDestinationResult_hi_lo_1 = {maskDestinationResult_hi_lo_hi_1, maskDestinationResult_hi_lo_lo_1};
  wire [7:0]    maskDestinationResult_hi_hi_lo_1 = {maskDestinationResult_hi_105, maskDestinationResult_lo_105, maskDestinationResult_hi_97, maskDestinationResult_lo_97};
  wire [7:0]    maskDestinationResult_hi_hi_hi_1 = {maskDestinationResult_hi_121, maskDestinationResult_lo_121, maskDestinationResult_hi_113, maskDestinationResult_lo_113};
  wire [15:0]   maskDestinationResult_hi_hi_1 = {maskDestinationResult_hi_hi_hi_1, maskDestinationResult_hi_hi_lo_1};
  wire [31:0]   maskDestinationResult_hi_129 = {maskDestinationResult_hi_hi_1, maskDestinationResult_hi_lo_1};
  wire [7:0]    maskDestinationResult_lo_lo_lo_2 = {maskDestinationResult_hi_10, maskDestinationResult_lo_10, maskDestinationResult_hi_2, maskDestinationResult_lo_2};
  wire [7:0]    maskDestinationResult_lo_lo_hi_2 = {maskDestinationResult_hi_26, maskDestinationResult_lo_26, maskDestinationResult_hi_18, maskDestinationResult_lo_18};
  wire [15:0]   maskDestinationResult_lo_lo_2 = {maskDestinationResult_lo_lo_hi_2, maskDestinationResult_lo_lo_lo_2};
  wire [7:0]    maskDestinationResult_lo_hi_lo_2 = {maskDestinationResult_hi_42, maskDestinationResult_lo_42, maskDestinationResult_hi_34, maskDestinationResult_lo_34};
  wire [7:0]    maskDestinationResult_lo_hi_hi_2 = {maskDestinationResult_hi_58, maskDestinationResult_lo_58, maskDestinationResult_hi_50, maskDestinationResult_lo_50};
  wire [15:0]   maskDestinationResult_lo_hi_2 = {maskDestinationResult_lo_hi_hi_2, maskDestinationResult_lo_hi_lo_2};
  wire [31:0]   maskDestinationResult_lo_130 = {maskDestinationResult_lo_hi_2, maskDestinationResult_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_lo_lo_2 = {maskDestinationResult_hi_74, maskDestinationResult_lo_74, maskDestinationResult_hi_66, maskDestinationResult_lo_66};
  wire [7:0]    maskDestinationResult_hi_lo_hi_2 = {maskDestinationResult_hi_90, maskDestinationResult_lo_90, maskDestinationResult_hi_82, maskDestinationResult_lo_82};
  wire [15:0]   maskDestinationResult_hi_lo_2 = {maskDestinationResult_hi_lo_hi_2, maskDestinationResult_hi_lo_lo_2};
  wire [7:0]    maskDestinationResult_hi_hi_lo_2 = {maskDestinationResult_hi_106, maskDestinationResult_lo_106, maskDestinationResult_hi_98, maskDestinationResult_lo_98};
  wire [7:0]    maskDestinationResult_hi_hi_hi_2 = {maskDestinationResult_hi_122, maskDestinationResult_lo_122, maskDestinationResult_hi_114, maskDestinationResult_lo_114};
  wire [15:0]   maskDestinationResult_hi_hi_2 = {maskDestinationResult_hi_hi_hi_2, maskDestinationResult_hi_hi_lo_2};
  wire [31:0]   maskDestinationResult_hi_130 = {maskDestinationResult_hi_hi_2, maskDestinationResult_hi_lo_2};
  wire [7:0]    maskDestinationResult_lo_lo_lo_3 = {maskDestinationResult_hi_11, maskDestinationResult_lo_11, maskDestinationResult_hi_3, maskDestinationResult_lo_3};
  wire [7:0]    maskDestinationResult_lo_lo_hi_3 = {maskDestinationResult_hi_27, maskDestinationResult_lo_27, maskDestinationResult_hi_19, maskDestinationResult_lo_19};
  wire [15:0]   maskDestinationResult_lo_lo_3 = {maskDestinationResult_lo_lo_hi_3, maskDestinationResult_lo_lo_lo_3};
  wire [7:0]    maskDestinationResult_lo_hi_lo_3 = {maskDestinationResult_hi_43, maskDestinationResult_lo_43, maskDestinationResult_hi_35, maskDestinationResult_lo_35};
  wire [7:0]    maskDestinationResult_lo_hi_hi_3 = {maskDestinationResult_hi_59, maskDestinationResult_lo_59, maskDestinationResult_hi_51, maskDestinationResult_lo_51};
  wire [15:0]   maskDestinationResult_lo_hi_3 = {maskDestinationResult_lo_hi_hi_3, maskDestinationResult_lo_hi_lo_3};
  wire [31:0]   maskDestinationResult_lo_131 = {maskDestinationResult_lo_hi_3, maskDestinationResult_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_lo_lo_3 = {maskDestinationResult_hi_75, maskDestinationResult_lo_75, maskDestinationResult_hi_67, maskDestinationResult_lo_67};
  wire [7:0]    maskDestinationResult_hi_lo_hi_3 = {maskDestinationResult_hi_91, maskDestinationResult_lo_91, maskDestinationResult_hi_83, maskDestinationResult_lo_83};
  wire [15:0]   maskDestinationResult_hi_lo_3 = {maskDestinationResult_hi_lo_hi_3, maskDestinationResult_hi_lo_lo_3};
  wire [7:0]    maskDestinationResult_hi_hi_lo_3 = {maskDestinationResult_hi_107, maskDestinationResult_lo_107, maskDestinationResult_hi_99, maskDestinationResult_lo_99};
  wire [7:0]    maskDestinationResult_hi_hi_hi_3 = {maskDestinationResult_hi_123, maskDestinationResult_lo_123, maskDestinationResult_hi_115, maskDestinationResult_lo_115};
  wire [15:0]   maskDestinationResult_hi_hi_3 = {maskDestinationResult_hi_hi_hi_3, maskDestinationResult_hi_hi_lo_3};
  wire [31:0]   maskDestinationResult_hi_131 = {maskDestinationResult_hi_hi_3, maskDestinationResult_hi_lo_3};
  wire [7:0]    maskDestinationResult_lo_lo_lo_4 = {maskDestinationResult_hi_12, maskDestinationResult_lo_12, maskDestinationResult_hi_4, maskDestinationResult_lo_4};
  wire [7:0]    maskDestinationResult_lo_lo_hi_4 = {maskDestinationResult_hi_28, maskDestinationResult_lo_28, maskDestinationResult_hi_20, maskDestinationResult_lo_20};
  wire [15:0]   maskDestinationResult_lo_lo_4 = {maskDestinationResult_lo_lo_hi_4, maskDestinationResult_lo_lo_lo_4};
  wire [7:0]    maskDestinationResult_lo_hi_lo_4 = {maskDestinationResult_hi_44, maskDestinationResult_lo_44, maskDestinationResult_hi_36, maskDestinationResult_lo_36};
  wire [7:0]    maskDestinationResult_lo_hi_hi_4 = {maskDestinationResult_hi_60, maskDestinationResult_lo_60, maskDestinationResult_hi_52, maskDestinationResult_lo_52};
  wire [15:0]   maskDestinationResult_lo_hi_4 = {maskDestinationResult_lo_hi_hi_4, maskDestinationResult_lo_hi_lo_4};
  wire [31:0]   maskDestinationResult_lo_132 = {maskDestinationResult_lo_hi_4, maskDestinationResult_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_lo_lo_4 = {maskDestinationResult_hi_76, maskDestinationResult_lo_76, maskDestinationResult_hi_68, maskDestinationResult_lo_68};
  wire [7:0]    maskDestinationResult_hi_lo_hi_4 = {maskDestinationResult_hi_92, maskDestinationResult_lo_92, maskDestinationResult_hi_84, maskDestinationResult_lo_84};
  wire [15:0]   maskDestinationResult_hi_lo_4 = {maskDestinationResult_hi_lo_hi_4, maskDestinationResult_hi_lo_lo_4};
  wire [7:0]    maskDestinationResult_hi_hi_lo_4 = {maskDestinationResult_hi_108, maskDestinationResult_lo_108, maskDestinationResult_hi_100, maskDestinationResult_lo_100};
  wire [7:0]    maskDestinationResult_hi_hi_hi_4 = {maskDestinationResult_hi_124, maskDestinationResult_lo_124, maskDestinationResult_hi_116, maskDestinationResult_lo_116};
  wire [15:0]   maskDestinationResult_hi_hi_4 = {maskDestinationResult_hi_hi_hi_4, maskDestinationResult_hi_hi_lo_4};
  wire [31:0]   maskDestinationResult_hi_132 = {maskDestinationResult_hi_hi_4, maskDestinationResult_hi_lo_4};
  wire [7:0]    maskDestinationResult_lo_lo_lo_5 = {maskDestinationResult_hi_13, maskDestinationResult_lo_13, maskDestinationResult_hi_5, maskDestinationResult_lo_5};
  wire [7:0]    maskDestinationResult_lo_lo_hi_5 = {maskDestinationResult_hi_29, maskDestinationResult_lo_29, maskDestinationResult_hi_21, maskDestinationResult_lo_21};
  wire [15:0]   maskDestinationResult_lo_lo_5 = {maskDestinationResult_lo_lo_hi_5, maskDestinationResult_lo_lo_lo_5};
  wire [7:0]    maskDestinationResult_lo_hi_lo_5 = {maskDestinationResult_hi_45, maskDestinationResult_lo_45, maskDestinationResult_hi_37, maskDestinationResult_lo_37};
  wire [7:0]    maskDestinationResult_lo_hi_hi_5 = {maskDestinationResult_hi_61, maskDestinationResult_lo_61, maskDestinationResult_hi_53, maskDestinationResult_lo_53};
  wire [15:0]   maskDestinationResult_lo_hi_5 = {maskDestinationResult_lo_hi_hi_5, maskDestinationResult_lo_hi_lo_5};
  wire [31:0]   maskDestinationResult_lo_133 = {maskDestinationResult_lo_hi_5, maskDestinationResult_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_lo_lo_5 = {maskDestinationResult_hi_77, maskDestinationResult_lo_77, maskDestinationResult_hi_69, maskDestinationResult_lo_69};
  wire [7:0]    maskDestinationResult_hi_lo_hi_5 = {maskDestinationResult_hi_93, maskDestinationResult_lo_93, maskDestinationResult_hi_85, maskDestinationResult_lo_85};
  wire [15:0]   maskDestinationResult_hi_lo_5 = {maskDestinationResult_hi_lo_hi_5, maskDestinationResult_hi_lo_lo_5};
  wire [7:0]    maskDestinationResult_hi_hi_lo_5 = {maskDestinationResult_hi_109, maskDestinationResult_lo_109, maskDestinationResult_hi_101, maskDestinationResult_lo_101};
  wire [7:0]    maskDestinationResult_hi_hi_hi_5 = {maskDestinationResult_hi_125, maskDestinationResult_lo_125, maskDestinationResult_hi_117, maskDestinationResult_lo_117};
  wire [15:0]   maskDestinationResult_hi_hi_5 = {maskDestinationResult_hi_hi_hi_5, maskDestinationResult_hi_hi_lo_5};
  wire [31:0]   maskDestinationResult_hi_133 = {maskDestinationResult_hi_hi_5, maskDestinationResult_hi_lo_5};
  wire [7:0]    maskDestinationResult_lo_lo_lo_6 = {maskDestinationResult_hi_14, maskDestinationResult_lo_14, maskDestinationResult_hi_6, maskDestinationResult_lo_6};
  wire [7:0]    maskDestinationResult_lo_lo_hi_6 = {maskDestinationResult_hi_30, maskDestinationResult_lo_30, maskDestinationResult_hi_22, maskDestinationResult_lo_22};
  wire [15:0]   maskDestinationResult_lo_lo_6 = {maskDestinationResult_lo_lo_hi_6, maskDestinationResult_lo_lo_lo_6};
  wire [7:0]    maskDestinationResult_lo_hi_lo_6 = {maskDestinationResult_hi_46, maskDestinationResult_lo_46, maskDestinationResult_hi_38, maskDestinationResult_lo_38};
  wire [7:0]    maskDestinationResult_lo_hi_hi_6 = {maskDestinationResult_hi_62, maskDestinationResult_lo_62, maskDestinationResult_hi_54, maskDestinationResult_lo_54};
  wire [15:0]   maskDestinationResult_lo_hi_6 = {maskDestinationResult_lo_hi_hi_6, maskDestinationResult_lo_hi_lo_6};
  wire [31:0]   maskDestinationResult_lo_134 = {maskDestinationResult_lo_hi_6, maskDestinationResult_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_lo_lo_6 = {maskDestinationResult_hi_78, maskDestinationResult_lo_78, maskDestinationResult_hi_70, maskDestinationResult_lo_70};
  wire [7:0]    maskDestinationResult_hi_lo_hi_6 = {maskDestinationResult_hi_94, maskDestinationResult_lo_94, maskDestinationResult_hi_86, maskDestinationResult_lo_86};
  wire [15:0]   maskDestinationResult_hi_lo_6 = {maskDestinationResult_hi_lo_hi_6, maskDestinationResult_hi_lo_lo_6};
  wire [7:0]    maskDestinationResult_hi_hi_lo_6 = {maskDestinationResult_hi_110, maskDestinationResult_lo_110, maskDestinationResult_hi_102, maskDestinationResult_lo_102};
  wire [7:0]    maskDestinationResult_hi_hi_hi_6 = {maskDestinationResult_hi_126, maskDestinationResult_lo_126, maskDestinationResult_hi_118, maskDestinationResult_lo_118};
  wire [15:0]   maskDestinationResult_hi_hi_6 = {maskDestinationResult_hi_hi_hi_6, maskDestinationResult_hi_hi_lo_6};
  wire [31:0]   maskDestinationResult_hi_134 = {maskDestinationResult_hi_hi_6, maskDestinationResult_hi_lo_6};
  wire [7:0]    maskDestinationResult_lo_lo_lo_7 = {maskDestinationResult_hi_15, maskDestinationResult_lo_15, maskDestinationResult_hi_7, maskDestinationResult_lo_7};
  wire [7:0]    maskDestinationResult_lo_lo_hi_7 = {maskDestinationResult_hi_31, maskDestinationResult_lo_31, maskDestinationResult_hi_23, maskDestinationResult_lo_23};
  wire [15:0]   maskDestinationResult_lo_lo_7 = {maskDestinationResult_lo_lo_hi_7, maskDestinationResult_lo_lo_lo_7};
  wire [7:0]    maskDestinationResult_lo_hi_lo_7 = {maskDestinationResult_hi_47, maskDestinationResult_lo_47, maskDestinationResult_hi_39, maskDestinationResult_lo_39};
  wire [7:0]    maskDestinationResult_lo_hi_hi_7 = {maskDestinationResult_hi_63, maskDestinationResult_lo_63, maskDestinationResult_hi_55, maskDestinationResult_lo_55};
  wire [15:0]   maskDestinationResult_lo_hi_7 = {maskDestinationResult_lo_hi_hi_7, maskDestinationResult_lo_hi_lo_7};
  wire [31:0]   maskDestinationResult_lo_135 = {maskDestinationResult_lo_hi_7, maskDestinationResult_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_lo_lo_7 = {maskDestinationResult_hi_79, maskDestinationResult_lo_79, maskDestinationResult_hi_71, maskDestinationResult_lo_71};
  wire [7:0]    maskDestinationResult_hi_lo_hi_7 = {maskDestinationResult_hi_95, maskDestinationResult_lo_95, maskDestinationResult_hi_87, maskDestinationResult_lo_87};
  wire [15:0]   maskDestinationResult_hi_lo_7 = {maskDestinationResult_hi_lo_hi_7, maskDestinationResult_hi_lo_lo_7};
  wire [7:0]    maskDestinationResult_hi_hi_lo_7 = {maskDestinationResult_hi_111, maskDestinationResult_lo_111, maskDestinationResult_hi_103, maskDestinationResult_lo_103};
  wire [7:0]    maskDestinationResult_hi_hi_hi_7 = {maskDestinationResult_hi_127, maskDestinationResult_lo_127, maskDestinationResult_hi_119, maskDestinationResult_lo_119};
  wire [15:0]   maskDestinationResult_hi_hi_7 = {maskDestinationResult_hi_hi_hi_7, maskDestinationResult_hi_hi_lo_7};
  wire [31:0]   maskDestinationResult_hi_135 = {maskDestinationResult_hi_hi_7, maskDestinationResult_hi_lo_7};
  wire [127:0]  maskDestinationResult_lo_lo_8 = {maskDestinationResult_hi_129, maskDestinationResult_lo_129, maskDestinationResult_hi_128, maskDestinationResult_lo_128};
  wire [127:0]  maskDestinationResult_lo_hi_8 = {maskDestinationResult_hi_131, maskDestinationResult_lo_131, maskDestinationResult_hi_130, maskDestinationResult_lo_130};
  wire [255:0]  maskDestinationResult_lo_136 = {maskDestinationResult_lo_hi_8, maskDestinationResult_lo_lo_8};
  wire [127:0]  maskDestinationResult_hi_lo_8 = {maskDestinationResult_hi_133, maskDestinationResult_lo_133, maskDestinationResult_hi_132, maskDestinationResult_lo_132};
  wire [127:0]  maskDestinationResult_hi_hi_8 = {maskDestinationResult_hi_135, maskDestinationResult_lo_135, maskDestinationResult_hi_134, maskDestinationResult_lo_134};
  wire [255:0]  maskDestinationResult_hi_136 = {maskDestinationResult_hi_hi_8, maskDestinationResult_hi_lo_8};
  wire [3:0]    maskDestinationResult_lo_lo_lo_8 = {sourceDataVec_1[1:0], sourceDataVec_0[1:0]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_8 = {sourceDataVec_3[1:0], sourceDataVec_2[1:0]};
  wire [7:0]    maskDestinationResult_lo_lo_9 = {maskDestinationResult_lo_lo_hi_8, maskDestinationResult_lo_lo_lo_8};
  wire [3:0]    maskDestinationResult_lo_hi_lo_8 = {sourceDataVec_5[1:0], sourceDataVec_4[1:0]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_8 = {sourceDataVec_7[1:0], sourceDataVec_6[1:0]};
  wire [7:0]    maskDestinationResult_lo_hi_9 = {maskDestinationResult_lo_hi_hi_8, maskDestinationResult_lo_hi_lo_8};
  wire [15:0]   maskDestinationResult_lo_137 = {maskDestinationResult_lo_hi_9, maskDestinationResult_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_lo_lo_8 = {sourceDataVec_9[1:0], sourceDataVec_8[1:0]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_8 = {sourceDataVec_11[1:0], sourceDataVec_10[1:0]};
  wire [7:0]    maskDestinationResult_hi_lo_9 = {maskDestinationResult_hi_lo_hi_8, maskDestinationResult_hi_lo_lo_8};
  wire [3:0]    maskDestinationResult_hi_hi_lo_8 = {sourceDataVec_13[1:0], sourceDataVec_12[1:0]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_8 = {sourceDataVec_15[1:0], sourceDataVec_14[1:0]};
  wire [7:0]    maskDestinationResult_hi_hi_9 = {maskDestinationResult_hi_hi_hi_8, maskDestinationResult_hi_hi_lo_8};
  wire [15:0]   maskDestinationResult_hi_137 = {maskDestinationResult_hi_hi_9, maskDestinationResult_hi_lo_9};
  wire [3:0]    maskDestinationResult_lo_lo_lo_9 = {sourceDataVec_1[3:2], sourceDataVec_0[3:2]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_9 = {sourceDataVec_3[3:2], sourceDataVec_2[3:2]};
  wire [7:0]    maskDestinationResult_lo_lo_10 = {maskDestinationResult_lo_lo_hi_9, maskDestinationResult_lo_lo_lo_9};
  wire [3:0]    maskDestinationResult_lo_hi_lo_9 = {sourceDataVec_5[3:2], sourceDataVec_4[3:2]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_9 = {sourceDataVec_7[3:2], sourceDataVec_6[3:2]};
  wire [7:0]    maskDestinationResult_lo_hi_10 = {maskDestinationResult_lo_hi_hi_9, maskDestinationResult_lo_hi_lo_9};
  wire [15:0]   maskDestinationResult_lo_138 = {maskDestinationResult_lo_hi_10, maskDestinationResult_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_lo_lo_9 = {sourceDataVec_9[3:2], sourceDataVec_8[3:2]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_9 = {sourceDataVec_11[3:2], sourceDataVec_10[3:2]};
  wire [7:0]    maskDestinationResult_hi_lo_10 = {maskDestinationResult_hi_lo_hi_9, maskDestinationResult_hi_lo_lo_9};
  wire [3:0]    maskDestinationResult_hi_hi_lo_9 = {sourceDataVec_13[3:2], sourceDataVec_12[3:2]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_9 = {sourceDataVec_15[3:2], sourceDataVec_14[3:2]};
  wire [7:0]    maskDestinationResult_hi_hi_10 = {maskDestinationResult_hi_hi_hi_9, maskDestinationResult_hi_hi_lo_9};
  wire [15:0]   maskDestinationResult_hi_138 = {maskDestinationResult_hi_hi_10, maskDestinationResult_hi_lo_10};
  wire [3:0]    maskDestinationResult_lo_lo_lo_10 = {sourceDataVec_1[5:4], sourceDataVec_0[5:4]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_10 = {sourceDataVec_3[5:4], sourceDataVec_2[5:4]};
  wire [7:0]    maskDestinationResult_lo_lo_11 = {maskDestinationResult_lo_lo_hi_10, maskDestinationResult_lo_lo_lo_10};
  wire [3:0]    maskDestinationResult_lo_hi_lo_10 = {sourceDataVec_5[5:4], sourceDataVec_4[5:4]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_10 = {sourceDataVec_7[5:4], sourceDataVec_6[5:4]};
  wire [7:0]    maskDestinationResult_lo_hi_11 = {maskDestinationResult_lo_hi_hi_10, maskDestinationResult_lo_hi_lo_10};
  wire [15:0]   maskDestinationResult_lo_139 = {maskDestinationResult_lo_hi_11, maskDestinationResult_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_lo_lo_10 = {sourceDataVec_9[5:4], sourceDataVec_8[5:4]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_10 = {sourceDataVec_11[5:4], sourceDataVec_10[5:4]};
  wire [7:0]    maskDestinationResult_hi_lo_11 = {maskDestinationResult_hi_lo_hi_10, maskDestinationResult_hi_lo_lo_10};
  wire [3:0]    maskDestinationResult_hi_hi_lo_10 = {sourceDataVec_13[5:4], sourceDataVec_12[5:4]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_10 = {sourceDataVec_15[5:4], sourceDataVec_14[5:4]};
  wire [7:0]    maskDestinationResult_hi_hi_11 = {maskDestinationResult_hi_hi_hi_10, maskDestinationResult_hi_hi_lo_10};
  wire [15:0]   maskDestinationResult_hi_139 = {maskDestinationResult_hi_hi_11, maskDestinationResult_hi_lo_11};
  wire [3:0]    maskDestinationResult_lo_lo_lo_11 = {sourceDataVec_1[7:6], sourceDataVec_0[7:6]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_11 = {sourceDataVec_3[7:6], sourceDataVec_2[7:6]};
  wire [7:0]    maskDestinationResult_lo_lo_12 = {maskDestinationResult_lo_lo_hi_11, maskDestinationResult_lo_lo_lo_11};
  wire [3:0]    maskDestinationResult_lo_hi_lo_11 = {sourceDataVec_5[7:6], sourceDataVec_4[7:6]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_11 = {sourceDataVec_7[7:6], sourceDataVec_6[7:6]};
  wire [7:0]    maskDestinationResult_lo_hi_12 = {maskDestinationResult_lo_hi_hi_11, maskDestinationResult_lo_hi_lo_11};
  wire [15:0]   maskDestinationResult_lo_140 = {maskDestinationResult_lo_hi_12, maskDestinationResult_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_lo_lo_11 = {sourceDataVec_9[7:6], sourceDataVec_8[7:6]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_11 = {sourceDataVec_11[7:6], sourceDataVec_10[7:6]};
  wire [7:0]    maskDestinationResult_hi_lo_12 = {maskDestinationResult_hi_lo_hi_11, maskDestinationResult_hi_lo_lo_11};
  wire [3:0]    maskDestinationResult_hi_hi_lo_11 = {sourceDataVec_13[7:6], sourceDataVec_12[7:6]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_11 = {sourceDataVec_15[7:6], sourceDataVec_14[7:6]};
  wire [7:0]    maskDestinationResult_hi_hi_12 = {maskDestinationResult_hi_hi_hi_11, maskDestinationResult_hi_hi_lo_11};
  wire [15:0]   maskDestinationResult_hi_140 = {maskDestinationResult_hi_hi_12, maskDestinationResult_hi_lo_12};
  wire [3:0]    maskDestinationResult_lo_lo_lo_12 = {sourceDataVec_1[9:8], sourceDataVec_0[9:8]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_12 = {sourceDataVec_3[9:8], sourceDataVec_2[9:8]};
  wire [7:0]    maskDestinationResult_lo_lo_13 = {maskDestinationResult_lo_lo_hi_12, maskDestinationResult_lo_lo_lo_12};
  wire [3:0]    maskDestinationResult_lo_hi_lo_12 = {sourceDataVec_5[9:8], sourceDataVec_4[9:8]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_12 = {sourceDataVec_7[9:8], sourceDataVec_6[9:8]};
  wire [7:0]    maskDestinationResult_lo_hi_13 = {maskDestinationResult_lo_hi_hi_12, maskDestinationResult_lo_hi_lo_12};
  wire [15:0]   maskDestinationResult_lo_141 = {maskDestinationResult_lo_hi_13, maskDestinationResult_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_lo_lo_12 = {sourceDataVec_9[9:8], sourceDataVec_8[9:8]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_12 = {sourceDataVec_11[9:8], sourceDataVec_10[9:8]};
  wire [7:0]    maskDestinationResult_hi_lo_13 = {maskDestinationResult_hi_lo_hi_12, maskDestinationResult_hi_lo_lo_12};
  wire [3:0]    maskDestinationResult_hi_hi_lo_12 = {sourceDataVec_13[9:8], sourceDataVec_12[9:8]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_12 = {sourceDataVec_15[9:8], sourceDataVec_14[9:8]};
  wire [7:0]    maskDestinationResult_hi_hi_13 = {maskDestinationResult_hi_hi_hi_12, maskDestinationResult_hi_hi_lo_12};
  wire [15:0]   maskDestinationResult_hi_141 = {maskDestinationResult_hi_hi_13, maskDestinationResult_hi_lo_13};
  wire [3:0]    maskDestinationResult_lo_lo_lo_13 = {sourceDataVec_1[11:10], sourceDataVec_0[11:10]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_13 = {sourceDataVec_3[11:10], sourceDataVec_2[11:10]};
  wire [7:0]    maskDestinationResult_lo_lo_14 = {maskDestinationResult_lo_lo_hi_13, maskDestinationResult_lo_lo_lo_13};
  wire [3:0]    maskDestinationResult_lo_hi_lo_13 = {sourceDataVec_5[11:10], sourceDataVec_4[11:10]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_13 = {sourceDataVec_7[11:10], sourceDataVec_6[11:10]};
  wire [7:0]    maskDestinationResult_lo_hi_14 = {maskDestinationResult_lo_hi_hi_13, maskDestinationResult_lo_hi_lo_13};
  wire [15:0]   maskDestinationResult_lo_142 = {maskDestinationResult_lo_hi_14, maskDestinationResult_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_lo_lo_13 = {sourceDataVec_9[11:10], sourceDataVec_8[11:10]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_13 = {sourceDataVec_11[11:10], sourceDataVec_10[11:10]};
  wire [7:0]    maskDestinationResult_hi_lo_14 = {maskDestinationResult_hi_lo_hi_13, maskDestinationResult_hi_lo_lo_13};
  wire [3:0]    maskDestinationResult_hi_hi_lo_13 = {sourceDataVec_13[11:10], sourceDataVec_12[11:10]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_13 = {sourceDataVec_15[11:10], sourceDataVec_14[11:10]};
  wire [7:0]    maskDestinationResult_hi_hi_14 = {maskDestinationResult_hi_hi_hi_13, maskDestinationResult_hi_hi_lo_13};
  wire [15:0]   maskDestinationResult_hi_142 = {maskDestinationResult_hi_hi_14, maskDestinationResult_hi_lo_14};
  wire [3:0]    maskDestinationResult_lo_lo_lo_14 = {sourceDataVec_1[13:12], sourceDataVec_0[13:12]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_14 = {sourceDataVec_3[13:12], sourceDataVec_2[13:12]};
  wire [7:0]    maskDestinationResult_lo_lo_15 = {maskDestinationResult_lo_lo_hi_14, maskDestinationResult_lo_lo_lo_14};
  wire [3:0]    maskDestinationResult_lo_hi_lo_14 = {sourceDataVec_5[13:12], sourceDataVec_4[13:12]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_14 = {sourceDataVec_7[13:12], sourceDataVec_6[13:12]};
  wire [7:0]    maskDestinationResult_lo_hi_15 = {maskDestinationResult_lo_hi_hi_14, maskDestinationResult_lo_hi_lo_14};
  wire [15:0]   maskDestinationResult_lo_143 = {maskDestinationResult_lo_hi_15, maskDestinationResult_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_lo_lo_14 = {sourceDataVec_9[13:12], sourceDataVec_8[13:12]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_14 = {sourceDataVec_11[13:12], sourceDataVec_10[13:12]};
  wire [7:0]    maskDestinationResult_hi_lo_15 = {maskDestinationResult_hi_lo_hi_14, maskDestinationResult_hi_lo_lo_14};
  wire [3:0]    maskDestinationResult_hi_hi_lo_14 = {sourceDataVec_13[13:12], sourceDataVec_12[13:12]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_14 = {sourceDataVec_15[13:12], sourceDataVec_14[13:12]};
  wire [7:0]    maskDestinationResult_hi_hi_15 = {maskDestinationResult_hi_hi_hi_14, maskDestinationResult_hi_hi_lo_14};
  wire [15:0]   maskDestinationResult_hi_143 = {maskDestinationResult_hi_hi_15, maskDestinationResult_hi_lo_15};
  wire [3:0]    maskDestinationResult_lo_lo_lo_15 = {sourceDataVec_1[15:14], sourceDataVec_0[15:14]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_15 = {sourceDataVec_3[15:14], sourceDataVec_2[15:14]};
  wire [7:0]    maskDestinationResult_lo_lo_16 = {maskDestinationResult_lo_lo_hi_15, maskDestinationResult_lo_lo_lo_15};
  wire [3:0]    maskDestinationResult_lo_hi_lo_15 = {sourceDataVec_5[15:14], sourceDataVec_4[15:14]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_15 = {sourceDataVec_7[15:14], sourceDataVec_6[15:14]};
  wire [7:0]    maskDestinationResult_lo_hi_16 = {maskDestinationResult_lo_hi_hi_15, maskDestinationResult_lo_hi_lo_15};
  wire [15:0]   maskDestinationResult_lo_144 = {maskDestinationResult_lo_hi_16, maskDestinationResult_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_lo_lo_15 = {sourceDataVec_9[15:14], sourceDataVec_8[15:14]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_15 = {sourceDataVec_11[15:14], sourceDataVec_10[15:14]};
  wire [7:0]    maskDestinationResult_hi_lo_16 = {maskDestinationResult_hi_lo_hi_15, maskDestinationResult_hi_lo_lo_15};
  wire [3:0]    maskDestinationResult_hi_hi_lo_15 = {sourceDataVec_13[15:14], sourceDataVec_12[15:14]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_15 = {sourceDataVec_15[15:14], sourceDataVec_14[15:14]};
  wire [7:0]    maskDestinationResult_hi_hi_16 = {maskDestinationResult_hi_hi_hi_15, maskDestinationResult_hi_hi_lo_15};
  wire [15:0]   maskDestinationResult_hi_144 = {maskDestinationResult_hi_hi_16, maskDestinationResult_hi_lo_16};
  wire [3:0]    maskDestinationResult_lo_lo_lo_16 = {sourceDataVec_1[17:16], sourceDataVec_0[17:16]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_16 = {sourceDataVec_3[17:16], sourceDataVec_2[17:16]};
  wire [7:0]    maskDestinationResult_lo_lo_17 = {maskDestinationResult_lo_lo_hi_16, maskDestinationResult_lo_lo_lo_16};
  wire [3:0]    maskDestinationResult_lo_hi_lo_16 = {sourceDataVec_5[17:16], sourceDataVec_4[17:16]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_16 = {sourceDataVec_7[17:16], sourceDataVec_6[17:16]};
  wire [7:0]    maskDestinationResult_lo_hi_17 = {maskDestinationResult_lo_hi_hi_16, maskDestinationResult_lo_hi_lo_16};
  wire [15:0]   maskDestinationResult_lo_145 = {maskDestinationResult_lo_hi_17, maskDestinationResult_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_lo_lo_16 = {sourceDataVec_9[17:16], sourceDataVec_8[17:16]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_16 = {sourceDataVec_11[17:16], sourceDataVec_10[17:16]};
  wire [7:0]    maskDestinationResult_hi_lo_17 = {maskDestinationResult_hi_lo_hi_16, maskDestinationResult_hi_lo_lo_16};
  wire [3:0]    maskDestinationResult_hi_hi_lo_16 = {sourceDataVec_13[17:16], sourceDataVec_12[17:16]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_16 = {sourceDataVec_15[17:16], sourceDataVec_14[17:16]};
  wire [7:0]    maskDestinationResult_hi_hi_17 = {maskDestinationResult_hi_hi_hi_16, maskDestinationResult_hi_hi_lo_16};
  wire [15:0]   maskDestinationResult_hi_145 = {maskDestinationResult_hi_hi_17, maskDestinationResult_hi_lo_17};
  wire [3:0]    maskDestinationResult_lo_lo_lo_17 = {sourceDataVec_1[19:18], sourceDataVec_0[19:18]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_17 = {sourceDataVec_3[19:18], sourceDataVec_2[19:18]};
  wire [7:0]    maskDestinationResult_lo_lo_18 = {maskDestinationResult_lo_lo_hi_17, maskDestinationResult_lo_lo_lo_17};
  wire [3:0]    maskDestinationResult_lo_hi_lo_17 = {sourceDataVec_5[19:18], sourceDataVec_4[19:18]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_17 = {sourceDataVec_7[19:18], sourceDataVec_6[19:18]};
  wire [7:0]    maskDestinationResult_lo_hi_18 = {maskDestinationResult_lo_hi_hi_17, maskDestinationResult_lo_hi_lo_17};
  wire [15:0]   maskDestinationResult_lo_146 = {maskDestinationResult_lo_hi_18, maskDestinationResult_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_lo_lo_17 = {sourceDataVec_9[19:18], sourceDataVec_8[19:18]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_17 = {sourceDataVec_11[19:18], sourceDataVec_10[19:18]};
  wire [7:0]    maskDestinationResult_hi_lo_18 = {maskDestinationResult_hi_lo_hi_17, maskDestinationResult_hi_lo_lo_17};
  wire [3:0]    maskDestinationResult_hi_hi_lo_17 = {sourceDataVec_13[19:18], sourceDataVec_12[19:18]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_17 = {sourceDataVec_15[19:18], sourceDataVec_14[19:18]};
  wire [7:0]    maskDestinationResult_hi_hi_18 = {maskDestinationResult_hi_hi_hi_17, maskDestinationResult_hi_hi_lo_17};
  wire [15:0]   maskDestinationResult_hi_146 = {maskDestinationResult_hi_hi_18, maskDestinationResult_hi_lo_18};
  wire [3:0]    maskDestinationResult_lo_lo_lo_18 = {sourceDataVec_1[21:20], sourceDataVec_0[21:20]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_18 = {sourceDataVec_3[21:20], sourceDataVec_2[21:20]};
  wire [7:0]    maskDestinationResult_lo_lo_19 = {maskDestinationResult_lo_lo_hi_18, maskDestinationResult_lo_lo_lo_18};
  wire [3:0]    maskDestinationResult_lo_hi_lo_18 = {sourceDataVec_5[21:20], sourceDataVec_4[21:20]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_18 = {sourceDataVec_7[21:20], sourceDataVec_6[21:20]};
  wire [7:0]    maskDestinationResult_lo_hi_19 = {maskDestinationResult_lo_hi_hi_18, maskDestinationResult_lo_hi_lo_18};
  wire [15:0]   maskDestinationResult_lo_147 = {maskDestinationResult_lo_hi_19, maskDestinationResult_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_lo_lo_18 = {sourceDataVec_9[21:20], sourceDataVec_8[21:20]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_18 = {sourceDataVec_11[21:20], sourceDataVec_10[21:20]};
  wire [7:0]    maskDestinationResult_hi_lo_19 = {maskDestinationResult_hi_lo_hi_18, maskDestinationResult_hi_lo_lo_18};
  wire [3:0]    maskDestinationResult_hi_hi_lo_18 = {sourceDataVec_13[21:20], sourceDataVec_12[21:20]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_18 = {sourceDataVec_15[21:20], sourceDataVec_14[21:20]};
  wire [7:0]    maskDestinationResult_hi_hi_19 = {maskDestinationResult_hi_hi_hi_18, maskDestinationResult_hi_hi_lo_18};
  wire [15:0]   maskDestinationResult_hi_147 = {maskDestinationResult_hi_hi_19, maskDestinationResult_hi_lo_19};
  wire [3:0]    maskDestinationResult_lo_lo_lo_19 = {sourceDataVec_1[23:22], sourceDataVec_0[23:22]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_19 = {sourceDataVec_3[23:22], sourceDataVec_2[23:22]};
  wire [7:0]    maskDestinationResult_lo_lo_20 = {maskDestinationResult_lo_lo_hi_19, maskDestinationResult_lo_lo_lo_19};
  wire [3:0]    maskDestinationResult_lo_hi_lo_19 = {sourceDataVec_5[23:22], sourceDataVec_4[23:22]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_19 = {sourceDataVec_7[23:22], sourceDataVec_6[23:22]};
  wire [7:0]    maskDestinationResult_lo_hi_20 = {maskDestinationResult_lo_hi_hi_19, maskDestinationResult_lo_hi_lo_19};
  wire [15:0]   maskDestinationResult_lo_148 = {maskDestinationResult_lo_hi_20, maskDestinationResult_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_lo_lo_19 = {sourceDataVec_9[23:22], sourceDataVec_8[23:22]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_19 = {sourceDataVec_11[23:22], sourceDataVec_10[23:22]};
  wire [7:0]    maskDestinationResult_hi_lo_20 = {maskDestinationResult_hi_lo_hi_19, maskDestinationResult_hi_lo_lo_19};
  wire [3:0]    maskDestinationResult_hi_hi_lo_19 = {sourceDataVec_13[23:22], sourceDataVec_12[23:22]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_19 = {sourceDataVec_15[23:22], sourceDataVec_14[23:22]};
  wire [7:0]    maskDestinationResult_hi_hi_20 = {maskDestinationResult_hi_hi_hi_19, maskDestinationResult_hi_hi_lo_19};
  wire [15:0]   maskDestinationResult_hi_148 = {maskDestinationResult_hi_hi_20, maskDestinationResult_hi_lo_20};
  wire [3:0]    maskDestinationResult_lo_lo_lo_20 = {sourceDataVec_1[25:24], sourceDataVec_0[25:24]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_20 = {sourceDataVec_3[25:24], sourceDataVec_2[25:24]};
  wire [7:0]    maskDestinationResult_lo_lo_21 = {maskDestinationResult_lo_lo_hi_20, maskDestinationResult_lo_lo_lo_20};
  wire [3:0]    maskDestinationResult_lo_hi_lo_20 = {sourceDataVec_5[25:24], sourceDataVec_4[25:24]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_20 = {sourceDataVec_7[25:24], sourceDataVec_6[25:24]};
  wire [7:0]    maskDestinationResult_lo_hi_21 = {maskDestinationResult_lo_hi_hi_20, maskDestinationResult_lo_hi_lo_20};
  wire [15:0]   maskDestinationResult_lo_149 = {maskDestinationResult_lo_hi_21, maskDestinationResult_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_lo_lo_20 = {sourceDataVec_9[25:24], sourceDataVec_8[25:24]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_20 = {sourceDataVec_11[25:24], sourceDataVec_10[25:24]};
  wire [7:0]    maskDestinationResult_hi_lo_21 = {maskDestinationResult_hi_lo_hi_20, maskDestinationResult_hi_lo_lo_20};
  wire [3:0]    maskDestinationResult_hi_hi_lo_20 = {sourceDataVec_13[25:24], sourceDataVec_12[25:24]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_20 = {sourceDataVec_15[25:24], sourceDataVec_14[25:24]};
  wire [7:0]    maskDestinationResult_hi_hi_21 = {maskDestinationResult_hi_hi_hi_20, maskDestinationResult_hi_hi_lo_20};
  wire [15:0]   maskDestinationResult_hi_149 = {maskDestinationResult_hi_hi_21, maskDestinationResult_hi_lo_21};
  wire [3:0]    maskDestinationResult_lo_lo_lo_21 = {sourceDataVec_1[27:26], sourceDataVec_0[27:26]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_21 = {sourceDataVec_3[27:26], sourceDataVec_2[27:26]};
  wire [7:0]    maskDestinationResult_lo_lo_22 = {maskDestinationResult_lo_lo_hi_21, maskDestinationResult_lo_lo_lo_21};
  wire [3:0]    maskDestinationResult_lo_hi_lo_21 = {sourceDataVec_5[27:26], sourceDataVec_4[27:26]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_21 = {sourceDataVec_7[27:26], sourceDataVec_6[27:26]};
  wire [7:0]    maskDestinationResult_lo_hi_22 = {maskDestinationResult_lo_hi_hi_21, maskDestinationResult_lo_hi_lo_21};
  wire [15:0]   maskDestinationResult_lo_150 = {maskDestinationResult_lo_hi_22, maskDestinationResult_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_lo_lo_21 = {sourceDataVec_9[27:26], sourceDataVec_8[27:26]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_21 = {sourceDataVec_11[27:26], sourceDataVec_10[27:26]};
  wire [7:0]    maskDestinationResult_hi_lo_22 = {maskDestinationResult_hi_lo_hi_21, maskDestinationResult_hi_lo_lo_21};
  wire [3:0]    maskDestinationResult_hi_hi_lo_21 = {sourceDataVec_13[27:26], sourceDataVec_12[27:26]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_21 = {sourceDataVec_15[27:26], sourceDataVec_14[27:26]};
  wire [7:0]    maskDestinationResult_hi_hi_22 = {maskDestinationResult_hi_hi_hi_21, maskDestinationResult_hi_hi_lo_21};
  wire [15:0]   maskDestinationResult_hi_150 = {maskDestinationResult_hi_hi_22, maskDestinationResult_hi_lo_22};
  wire [3:0]    maskDestinationResult_lo_lo_lo_22 = {sourceDataVec_1[29:28], sourceDataVec_0[29:28]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_22 = {sourceDataVec_3[29:28], sourceDataVec_2[29:28]};
  wire [7:0]    maskDestinationResult_lo_lo_23 = {maskDestinationResult_lo_lo_hi_22, maskDestinationResult_lo_lo_lo_22};
  wire [3:0]    maskDestinationResult_lo_hi_lo_22 = {sourceDataVec_5[29:28], sourceDataVec_4[29:28]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_22 = {sourceDataVec_7[29:28], sourceDataVec_6[29:28]};
  wire [7:0]    maskDestinationResult_lo_hi_23 = {maskDestinationResult_lo_hi_hi_22, maskDestinationResult_lo_hi_lo_22};
  wire [15:0]   maskDestinationResult_lo_151 = {maskDestinationResult_lo_hi_23, maskDestinationResult_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_lo_lo_22 = {sourceDataVec_9[29:28], sourceDataVec_8[29:28]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_22 = {sourceDataVec_11[29:28], sourceDataVec_10[29:28]};
  wire [7:0]    maskDestinationResult_hi_lo_23 = {maskDestinationResult_hi_lo_hi_22, maskDestinationResult_hi_lo_lo_22};
  wire [3:0]    maskDestinationResult_hi_hi_lo_22 = {sourceDataVec_13[29:28], sourceDataVec_12[29:28]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_22 = {sourceDataVec_15[29:28], sourceDataVec_14[29:28]};
  wire [7:0]    maskDestinationResult_hi_hi_23 = {maskDestinationResult_hi_hi_hi_22, maskDestinationResult_hi_hi_lo_22};
  wire [15:0]   maskDestinationResult_hi_151 = {maskDestinationResult_hi_hi_23, maskDestinationResult_hi_lo_23};
  wire [3:0]    maskDestinationResult_lo_lo_lo_23 = {sourceDataVec_1[31:30], sourceDataVec_0[31:30]};
  wire [3:0]    maskDestinationResult_lo_lo_hi_23 = {sourceDataVec_3[31:30], sourceDataVec_2[31:30]};
  wire [7:0]    maskDestinationResult_lo_lo_24 = {maskDestinationResult_lo_lo_hi_23, maskDestinationResult_lo_lo_lo_23};
  wire [3:0]    maskDestinationResult_lo_hi_lo_23 = {sourceDataVec_5[31:30], sourceDataVec_4[31:30]};
  wire [3:0]    maskDestinationResult_lo_hi_hi_23 = {sourceDataVec_7[31:30], sourceDataVec_6[31:30]};
  wire [7:0]    maskDestinationResult_lo_hi_24 = {maskDestinationResult_lo_hi_hi_23, maskDestinationResult_lo_hi_lo_23};
  wire [15:0]   maskDestinationResult_lo_152 = {maskDestinationResult_lo_hi_24, maskDestinationResult_lo_lo_24};
  wire [3:0]    maskDestinationResult_hi_lo_lo_23 = {sourceDataVec_9[31:30], sourceDataVec_8[31:30]};
  wire [3:0]    maskDestinationResult_hi_lo_hi_23 = {sourceDataVec_11[31:30], sourceDataVec_10[31:30]};
  wire [7:0]    maskDestinationResult_hi_lo_24 = {maskDestinationResult_hi_lo_hi_23, maskDestinationResult_hi_lo_lo_23};
  wire [3:0]    maskDestinationResult_hi_hi_lo_23 = {sourceDataVec_13[31:30], sourceDataVec_12[31:30]};
  wire [3:0]    maskDestinationResult_hi_hi_hi_23 = {sourceDataVec_15[31:30], sourceDataVec_14[31:30]};
  wire [7:0]    maskDestinationResult_hi_hi_24 = {maskDestinationResult_hi_hi_hi_23, maskDestinationResult_hi_hi_lo_23};
  wire [15:0]   maskDestinationResult_hi_152 = {maskDestinationResult_hi_hi_24, maskDestinationResult_hi_lo_24};
  wire [63:0]   maskDestinationResult_lo_lo_lo_24 = {maskDestinationResult_hi_138, maskDestinationResult_lo_138, maskDestinationResult_hi_137, maskDestinationResult_lo_137};
  wire [63:0]   maskDestinationResult_lo_lo_hi_24 = {maskDestinationResult_hi_140, maskDestinationResult_lo_140, maskDestinationResult_hi_139, maskDestinationResult_lo_139};
  wire [127:0]  maskDestinationResult_lo_lo_25 = {maskDestinationResult_lo_lo_hi_24, maskDestinationResult_lo_lo_lo_24};
  wire [63:0]   maskDestinationResult_lo_hi_lo_24 = {maskDestinationResult_hi_142, maskDestinationResult_lo_142, maskDestinationResult_hi_141, maskDestinationResult_lo_141};
  wire [63:0]   maskDestinationResult_lo_hi_hi_24 = {maskDestinationResult_hi_144, maskDestinationResult_lo_144, maskDestinationResult_hi_143, maskDestinationResult_lo_143};
  wire [127:0]  maskDestinationResult_lo_hi_25 = {maskDestinationResult_lo_hi_hi_24, maskDestinationResult_lo_hi_lo_24};
  wire [255:0]  maskDestinationResult_lo_153 = {maskDestinationResult_lo_hi_25, maskDestinationResult_lo_lo_25};
  wire [63:0]   maskDestinationResult_hi_lo_lo_24 = {maskDestinationResult_hi_146, maskDestinationResult_lo_146, maskDestinationResult_hi_145, maskDestinationResult_lo_145};
  wire [63:0]   maskDestinationResult_hi_lo_hi_24 = {maskDestinationResult_hi_148, maskDestinationResult_lo_148, maskDestinationResult_hi_147, maskDestinationResult_lo_147};
  wire [127:0]  maskDestinationResult_hi_lo_25 = {maskDestinationResult_hi_lo_hi_24, maskDestinationResult_hi_lo_lo_24};
  wire [63:0]   maskDestinationResult_hi_hi_lo_24 = {maskDestinationResult_hi_150, maskDestinationResult_lo_150, maskDestinationResult_hi_149, maskDestinationResult_lo_149};
  wire [63:0]   maskDestinationResult_hi_hi_hi_24 = {maskDestinationResult_hi_152, maskDestinationResult_lo_152, maskDestinationResult_hi_151, maskDestinationResult_lo_151};
  wire [127:0]  maskDestinationResult_hi_hi_25 = {maskDestinationResult_hi_hi_hi_24, maskDestinationResult_hi_hi_lo_24};
  wire [255:0]  maskDestinationResult_hi_153 = {maskDestinationResult_hi_hi_25, maskDestinationResult_hi_lo_25};
  wire [1:0]    maskDestinationResult_lo_lo_lo_25 = {sourceDataVec_1[0], sourceDataVec_0[0]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_25 = {sourceDataVec_3[0], sourceDataVec_2[0]};
  wire [3:0]    maskDestinationResult_lo_lo_26 = {maskDestinationResult_lo_lo_hi_25, maskDestinationResult_lo_lo_lo_25};
  wire [1:0]    maskDestinationResult_lo_hi_lo_25 = {sourceDataVec_5[0], sourceDataVec_4[0]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_25 = {sourceDataVec_7[0], sourceDataVec_6[0]};
  wire [3:0]    maskDestinationResult_lo_hi_26 = {maskDestinationResult_lo_hi_hi_25, maskDestinationResult_lo_hi_lo_25};
  wire [7:0]    maskDestinationResult_lo_154 = {maskDestinationResult_lo_hi_26, maskDestinationResult_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_lo_lo_25 = {sourceDataVec_9[0], sourceDataVec_8[0]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_25 = {sourceDataVec_11[0], sourceDataVec_10[0]};
  wire [3:0]    maskDestinationResult_hi_lo_26 = {maskDestinationResult_hi_lo_hi_25, maskDestinationResult_hi_lo_lo_25};
  wire [1:0]    maskDestinationResult_hi_hi_lo_25 = {sourceDataVec_13[0], sourceDataVec_12[0]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_25 = {sourceDataVec_15[0], sourceDataVec_14[0]};
  wire [3:0]    maskDestinationResult_hi_hi_26 = {maskDestinationResult_hi_hi_hi_25, maskDestinationResult_hi_hi_lo_25};
  wire [7:0]    maskDestinationResult_hi_154 = {maskDestinationResult_hi_hi_26, maskDestinationResult_hi_lo_26};
  wire [1:0]    maskDestinationResult_lo_lo_lo_26 = {sourceDataVec_1[1], sourceDataVec_0[1]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_26 = {sourceDataVec_3[1], sourceDataVec_2[1]};
  wire [3:0]    maskDestinationResult_lo_lo_27 = {maskDestinationResult_lo_lo_hi_26, maskDestinationResult_lo_lo_lo_26};
  wire [1:0]    maskDestinationResult_lo_hi_lo_26 = {sourceDataVec_5[1], sourceDataVec_4[1]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_26 = {sourceDataVec_7[1], sourceDataVec_6[1]};
  wire [3:0]    maskDestinationResult_lo_hi_27 = {maskDestinationResult_lo_hi_hi_26, maskDestinationResult_lo_hi_lo_26};
  wire [7:0]    maskDestinationResult_lo_155 = {maskDestinationResult_lo_hi_27, maskDestinationResult_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_lo_lo_26 = {sourceDataVec_9[1], sourceDataVec_8[1]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_26 = {sourceDataVec_11[1], sourceDataVec_10[1]};
  wire [3:0]    maskDestinationResult_hi_lo_27 = {maskDestinationResult_hi_lo_hi_26, maskDestinationResult_hi_lo_lo_26};
  wire [1:0]    maskDestinationResult_hi_hi_lo_26 = {sourceDataVec_13[1], sourceDataVec_12[1]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_26 = {sourceDataVec_15[1], sourceDataVec_14[1]};
  wire [3:0]    maskDestinationResult_hi_hi_27 = {maskDestinationResult_hi_hi_hi_26, maskDestinationResult_hi_hi_lo_26};
  wire [7:0]    maskDestinationResult_hi_155 = {maskDestinationResult_hi_hi_27, maskDestinationResult_hi_lo_27};
  wire [1:0]    maskDestinationResult_lo_lo_lo_27 = {sourceDataVec_1[2], sourceDataVec_0[2]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_27 = {sourceDataVec_3[2], sourceDataVec_2[2]};
  wire [3:0]    maskDestinationResult_lo_lo_28 = {maskDestinationResult_lo_lo_hi_27, maskDestinationResult_lo_lo_lo_27};
  wire [1:0]    maskDestinationResult_lo_hi_lo_27 = {sourceDataVec_5[2], sourceDataVec_4[2]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_27 = {sourceDataVec_7[2], sourceDataVec_6[2]};
  wire [3:0]    maskDestinationResult_lo_hi_28 = {maskDestinationResult_lo_hi_hi_27, maskDestinationResult_lo_hi_lo_27};
  wire [7:0]    maskDestinationResult_lo_156 = {maskDestinationResult_lo_hi_28, maskDestinationResult_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_lo_lo_27 = {sourceDataVec_9[2], sourceDataVec_8[2]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_27 = {sourceDataVec_11[2], sourceDataVec_10[2]};
  wire [3:0]    maskDestinationResult_hi_lo_28 = {maskDestinationResult_hi_lo_hi_27, maskDestinationResult_hi_lo_lo_27};
  wire [1:0]    maskDestinationResult_hi_hi_lo_27 = {sourceDataVec_13[2], sourceDataVec_12[2]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_27 = {sourceDataVec_15[2], sourceDataVec_14[2]};
  wire [3:0]    maskDestinationResult_hi_hi_28 = {maskDestinationResult_hi_hi_hi_27, maskDestinationResult_hi_hi_lo_27};
  wire [7:0]    maskDestinationResult_hi_156 = {maskDestinationResult_hi_hi_28, maskDestinationResult_hi_lo_28};
  wire [1:0]    maskDestinationResult_lo_lo_lo_28 = {sourceDataVec_1[3], sourceDataVec_0[3]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_28 = {sourceDataVec_3[3], sourceDataVec_2[3]};
  wire [3:0]    maskDestinationResult_lo_lo_29 = {maskDestinationResult_lo_lo_hi_28, maskDestinationResult_lo_lo_lo_28};
  wire [1:0]    maskDestinationResult_lo_hi_lo_28 = {sourceDataVec_5[3], sourceDataVec_4[3]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_28 = {sourceDataVec_7[3], sourceDataVec_6[3]};
  wire [3:0]    maskDestinationResult_lo_hi_29 = {maskDestinationResult_lo_hi_hi_28, maskDestinationResult_lo_hi_lo_28};
  wire [7:0]    maskDestinationResult_lo_157 = {maskDestinationResult_lo_hi_29, maskDestinationResult_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_lo_lo_28 = {sourceDataVec_9[3], sourceDataVec_8[3]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_28 = {sourceDataVec_11[3], sourceDataVec_10[3]};
  wire [3:0]    maskDestinationResult_hi_lo_29 = {maskDestinationResult_hi_lo_hi_28, maskDestinationResult_hi_lo_lo_28};
  wire [1:0]    maskDestinationResult_hi_hi_lo_28 = {sourceDataVec_13[3], sourceDataVec_12[3]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_28 = {sourceDataVec_15[3], sourceDataVec_14[3]};
  wire [3:0]    maskDestinationResult_hi_hi_29 = {maskDestinationResult_hi_hi_hi_28, maskDestinationResult_hi_hi_lo_28};
  wire [7:0]    maskDestinationResult_hi_157 = {maskDestinationResult_hi_hi_29, maskDestinationResult_hi_lo_29};
  wire [1:0]    maskDestinationResult_lo_lo_lo_29 = {sourceDataVec_1[4], sourceDataVec_0[4]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_29 = {sourceDataVec_3[4], sourceDataVec_2[4]};
  wire [3:0]    maskDestinationResult_lo_lo_30 = {maskDestinationResult_lo_lo_hi_29, maskDestinationResult_lo_lo_lo_29};
  wire [1:0]    maskDestinationResult_lo_hi_lo_29 = {sourceDataVec_5[4], sourceDataVec_4[4]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_29 = {sourceDataVec_7[4], sourceDataVec_6[4]};
  wire [3:0]    maskDestinationResult_lo_hi_30 = {maskDestinationResult_lo_hi_hi_29, maskDestinationResult_lo_hi_lo_29};
  wire [7:0]    maskDestinationResult_lo_158 = {maskDestinationResult_lo_hi_30, maskDestinationResult_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_lo_lo_29 = {sourceDataVec_9[4], sourceDataVec_8[4]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_29 = {sourceDataVec_11[4], sourceDataVec_10[4]};
  wire [3:0]    maskDestinationResult_hi_lo_30 = {maskDestinationResult_hi_lo_hi_29, maskDestinationResult_hi_lo_lo_29};
  wire [1:0]    maskDestinationResult_hi_hi_lo_29 = {sourceDataVec_13[4], sourceDataVec_12[4]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_29 = {sourceDataVec_15[4], sourceDataVec_14[4]};
  wire [3:0]    maskDestinationResult_hi_hi_30 = {maskDestinationResult_hi_hi_hi_29, maskDestinationResult_hi_hi_lo_29};
  wire [7:0]    maskDestinationResult_hi_158 = {maskDestinationResult_hi_hi_30, maskDestinationResult_hi_lo_30};
  wire [1:0]    maskDestinationResult_lo_lo_lo_30 = {sourceDataVec_1[5], sourceDataVec_0[5]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_30 = {sourceDataVec_3[5], sourceDataVec_2[5]};
  wire [3:0]    maskDestinationResult_lo_lo_31 = {maskDestinationResult_lo_lo_hi_30, maskDestinationResult_lo_lo_lo_30};
  wire [1:0]    maskDestinationResult_lo_hi_lo_30 = {sourceDataVec_5[5], sourceDataVec_4[5]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_30 = {sourceDataVec_7[5], sourceDataVec_6[5]};
  wire [3:0]    maskDestinationResult_lo_hi_31 = {maskDestinationResult_lo_hi_hi_30, maskDestinationResult_lo_hi_lo_30};
  wire [7:0]    maskDestinationResult_lo_159 = {maskDestinationResult_lo_hi_31, maskDestinationResult_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_lo_lo_30 = {sourceDataVec_9[5], sourceDataVec_8[5]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_30 = {sourceDataVec_11[5], sourceDataVec_10[5]};
  wire [3:0]    maskDestinationResult_hi_lo_31 = {maskDestinationResult_hi_lo_hi_30, maskDestinationResult_hi_lo_lo_30};
  wire [1:0]    maskDestinationResult_hi_hi_lo_30 = {sourceDataVec_13[5], sourceDataVec_12[5]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_30 = {sourceDataVec_15[5], sourceDataVec_14[5]};
  wire [3:0]    maskDestinationResult_hi_hi_31 = {maskDestinationResult_hi_hi_hi_30, maskDestinationResult_hi_hi_lo_30};
  wire [7:0]    maskDestinationResult_hi_159 = {maskDestinationResult_hi_hi_31, maskDestinationResult_hi_lo_31};
  wire [1:0]    maskDestinationResult_lo_lo_lo_31 = {sourceDataVec_1[6], sourceDataVec_0[6]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_31 = {sourceDataVec_3[6], sourceDataVec_2[6]};
  wire [3:0]    maskDestinationResult_lo_lo_32 = {maskDestinationResult_lo_lo_hi_31, maskDestinationResult_lo_lo_lo_31};
  wire [1:0]    maskDestinationResult_lo_hi_lo_31 = {sourceDataVec_5[6], sourceDataVec_4[6]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_31 = {sourceDataVec_7[6], sourceDataVec_6[6]};
  wire [3:0]    maskDestinationResult_lo_hi_32 = {maskDestinationResult_lo_hi_hi_31, maskDestinationResult_lo_hi_lo_31};
  wire [7:0]    maskDestinationResult_lo_160 = {maskDestinationResult_lo_hi_32, maskDestinationResult_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_lo_lo_31 = {sourceDataVec_9[6], sourceDataVec_8[6]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_31 = {sourceDataVec_11[6], sourceDataVec_10[6]};
  wire [3:0]    maskDestinationResult_hi_lo_32 = {maskDestinationResult_hi_lo_hi_31, maskDestinationResult_hi_lo_lo_31};
  wire [1:0]    maskDestinationResult_hi_hi_lo_31 = {sourceDataVec_13[6], sourceDataVec_12[6]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_31 = {sourceDataVec_15[6], sourceDataVec_14[6]};
  wire [3:0]    maskDestinationResult_hi_hi_32 = {maskDestinationResult_hi_hi_hi_31, maskDestinationResult_hi_hi_lo_31};
  wire [7:0]    maskDestinationResult_hi_160 = {maskDestinationResult_hi_hi_32, maskDestinationResult_hi_lo_32};
  wire [1:0]    maskDestinationResult_lo_lo_lo_32 = {sourceDataVec_1[7], sourceDataVec_0[7]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_32 = {sourceDataVec_3[7], sourceDataVec_2[7]};
  wire [3:0]    maskDestinationResult_lo_lo_33 = {maskDestinationResult_lo_lo_hi_32, maskDestinationResult_lo_lo_lo_32};
  wire [1:0]    maskDestinationResult_lo_hi_lo_32 = {sourceDataVec_5[7], sourceDataVec_4[7]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_32 = {sourceDataVec_7[7], sourceDataVec_6[7]};
  wire [3:0]    maskDestinationResult_lo_hi_33 = {maskDestinationResult_lo_hi_hi_32, maskDestinationResult_lo_hi_lo_32};
  wire [7:0]    maskDestinationResult_lo_161 = {maskDestinationResult_lo_hi_33, maskDestinationResult_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_lo_lo_32 = {sourceDataVec_9[7], sourceDataVec_8[7]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_32 = {sourceDataVec_11[7], sourceDataVec_10[7]};
  wire [3:0]    maskDestinationResult_hi_lo_33 = {maskDestinationResult_hi_lo_hi_32, maskDestinationResult_hi_lo_lo_32};
  wire [1:0]    maskDestinationResult_hi_hi_lo_32 = {sourceDataVec_13[7], sourceDataVec_12[7]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_32 = {sourceDataVec_15[7], sourceDataVec_14[7]};
  wire [3:0]    maskDestinationResult_hi_hi_33 = {maskDestinationResult_hi_hi_hi_32, maskDestinationResult_hi_hi_lo_32};
  wire [7:0]    maskDestinationResult_hi_161 = {maskDestinationResult_hi_hi_33, maskDestinationResult_hi_lo_33};
  wire [1:0]    maskDestinationResult_lo_lo_lo_33 = {sourceDataVec_1[8], sourceDataVec_0[8]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_33 = {sourceDataVec_3[8], sourceDataVec_2[8]};
  wire [3:0]    maskDestinationResult_lo_lo_34 = {maskDestinationResult_lo_lo_hi_33, maskDestinationResult_lo_lo_lo_33};
  wire [1:0]    maskDestinationResult_lo_hi_lo_33 = {sourceDataVec_5[8], sourceDataVec_4[8]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_33 = {sourceDataVec_7[8], sourceDataVec_6[8]};
  wire [3:0]    maskDestinationResult_lo_hi_34 = {maskDestinationResult_lo_hi_hi_33, maskDestinationResult_lo_hi_lo_33};
  wire [7:0]    maskDestinationResult_lo_162 = {maskDestinationResult_lo_hi_34, maskDestinationResult_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_lo_lo_33 = {sourceDataVec_9[8], sourceDataVec_8[8]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_33 = {sourceDataVec_11[8], sourceDataVec_10[8]};
  wire [3:0]    maskDestinationResult_hi_lo_34 = {maskDestinationResult_hi_lo_hi_33, maskDestinationResult_hi_lo_lo_33};
  wire [1:0]    maskDestinationResult_hi_hi_lo_33 = {sourceDataVec_13[8], sourceDataVec_12[8]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_33 = {sourceDataVec_15[8], sourceDataVec_14[8]};
  wire [3:0]    maskDestinationResult_hi_hi_34 = {maskDestinationResult_hi_hi_hi_33, maskDestinationResult_hi_hi_lo_33};
  wire [7:0]    maskDestinationResult_hi_162 = {maskDestinationResult_hi_hi_34, maskDestinationResult_hi_lo_34};
  wire [1:0]    maskDestinationResult_lo_lo_lo_34 = {sourceDataVec_1[9], sourceDataVec_0[9]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_34 = {sourceDataVec_3[9], sourceDataVec_2[9]};
  wire [3:0]    maskDestinationResult_lo_lo_35 = {maskDestinationResult_lo_lo_hi_34, maskDestinationResult_lo_lo_lo_34};
  wire [1:0]    maskDestinationResult_lo_hi_lo_34 = {sourceDataVec_5[9], sourceDataVec_4[9]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_34 = {sourceDataVec_7[9], sourceDataVec_6[9]};
  wire [3:0]    maskDestinationResult_lo_hi_35 = {maskDestinationResult_lo_hi_hi_34, maskDestinationResult_lo_hi_lo_34};
  wire [7:0]    maskDestinationResult_lo_163 = {maskDestinationResult_lo_hi_35, maskDestinationResult_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_lo_lo_34 = {sourceDataVec_9[9], sourceDataVec_8[9]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_34 = {sourceDataVec_11[9], sourceDataVec_10[9]};
  wire [3:0]    maskDestinationResult_hi_lo_35 = {maskDestinationResult_hi_lo_hi_34, maskDestinationResult_hi_lo_lo_34};
  wire [1:0]    maskDestinationResult_hi_hi_lo_34 = {sourceDataVec_13[9], sourceDataVec_12[9]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_34 = {sourceDataVec_15[9], sourceDataVec_14[9]};
  wire [3:0]    maskDestinationResult_hi_hi_35 = {maskDestinationResult_hi_hi_hi_34, maskDestinationResult_hi_hi_lo_34};
  wire [7:0]    maskDestinationResult_hi_163 = {maskDestinationResult_hi_hi_35, maskDestinationResult_hi_lo_35};
  wire [1:0]    maskDestinationResult_lo_lo_lo_35 = {sourceDataVec_1[10], sourceDataVec_0[10]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_35 = {sourceDataVec_3[10], sourceDataVec_2[10]};
  wire [3:0]    maskDestinationResult_lo_lo_36 = {maskDestinationResult_lo_lo_hi_35, maskDestinationResult_lo_lo_lo_35};
  wire [1:0]    maskDestinationResult_lo_hi_lo_35 = {sourceDataVec_5[10], sourceDataVec_4[10]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_35 = {sourceDataVec_7[10], sourceDataVec_6[10]};
  wire [3:0]    maskDestinationResult_lo_hi_36 = {maskDestinationResult_lo_hi_hi_35, maskDestinationResult_lo_hi_lo_35};
  wire [7:0]    maskDestinationResult_lo_164 = {maskDestinationResult_lo_hi_36, maskDestinationResult_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_lo_lo_35 = {sourceDataVec_9[10], sourceDataVec_8[10]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_35 = {sourceDataVec_11[10], sourceDataVec_10[10]};
  wire [3:0]    maskDestinationResult_hi_lo_36 = {maskDestinationResult_hi_lo_hi_35, maskDestinationResult_hi_lo_lo_35};
  wire [1:0]    maskDestinationResult_hi_hi_lo_35 = {sourceDataVec_13[10], sourceDataVec_12[10]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_35 = {sourceDataVec_15[10], sourceDataVec_14[10]};
  wire [3:0]    maskDestinationResult_hi_hi_36 = {maskDestinationResult_hi_hi_hi_35, maskDestinationResult_hi_hi_lo_35};
  wire [7:0]    maskDestinationResult_hi_164 = {maskDestinationResult_hi_hi_36, maskDestinationResult_hi_lo_36};
  wire [1:0]    maskDestinationResult_lo_lo_lo_36 = {sourceDataVec_1[11], sourceDataVec_0[11]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_36 = {sourceDataVec_3[11], sourceDataVec_2[11]};
  wire [3:0]    maskDestinationResult_lo_lo_37 = {maskDestinationResult_lo_lo_hi_36, maskDestinationResult_lo_lo_lo_36};
  wire [1:0]    maskDestinationResult_lo_hi_lo_36 = {sourceDataVec_5[11], sourceDataVec_4[11]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_36 = {sourceDataVec_7[11], sourceDataVec_6[11]};
  wire [3:0]    maskDestinationResult_lo_hi_37 = {maskDestinationResult_lo_hi_hi_36, maskDestinationResult_lo_hi_lo_36};
  wire [7:0]    maskDestinationResult_lo_165 = {maskDestinationResult_lo_hi_37, maskDestinationResult_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_lo_lo_36 = {sourceDataVec_9[11], sourceDataVec_8[11]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_36 = {sourceDataVec_11[11], sourceDataVec_10[11]};
  wire [3:0]    maskDestinationResult_hi_lo_37 = {maskDestinationResult_hi_lo_hi_36, maskDestinationResult_hi_lo_lo_36};
  wire [1:0]    maskDestinationResult_hi_hi_lo_36 = {sourceDataVec_13[11], sourceDataVec_12[11]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_36 = {sourceDataVec_15[11], sourceDataVec_14[11]};
  wire [3:0]    maskDestinationResult_hi_hi_37 = {maskDestinationResult_hi_hi_hi_36, maskDestinationResult_hi_hi_lo_36};
  wire [7:0]    maskDestinationResult_hi_165 = {maskDestinationResult_hi_hi_37, maskDestinationResult_hi_lo_37};
  wire [1:0]    maskDestinationResult_lo_lo_lo_37 = {sourceDataVec_1[12], sourceDataVec_0[12]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_37 = {sourceDataVec_3[12], sourceDataVec_2[12]};
  wire [3:0]    maskDestinationResult_lo_lo_38 = {maskDestinationResult_lo_lo_hi_37, maskDestinationResult_lo_lo_lo_37};
  wire [1:0]    maskDestinationResult_lo_hi_lo_37 = {sourceDataVec_5[12], sourceDataVec_4[12]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_37 = {sourceDataVec_7[12], sourceDataVec_6[12]};
  wire [3:0]    maskDestinationResult_lo_hi_38 = {maskDestinationResult_lo_hi_hi_37, maskDestinationResult_lo_hi_lo_37};
  wire [7:0]    maskDestinationResult_lo_166 = {maskDestinationResult_lo_hi_38, maskDestinationResult_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_lo_lo_37 = {sourceDataVec_9[12], sourceDataVec_8[12]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_37 = {sourceDataVec_11[12], sourceDataVec_10[12]};
  wire [3:0]    maskDestinationResult_hi_lo_38 = {maskDestinationResult_hi_lo_hi_37, maskDestinationResult_hi_lo_lo_37};
  wire [1:0]    maskDestinationResult_hi_hi_lo_37 = {sourceDataVec_13[12], sourceDataVec_12[12]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_37 = {sourceDataVec_15[12], sourceDataVec_14[12]};
  wire [3:0]    maskDestinationResult_hi_hi_38 = {maskDestinationResult_hi_hi_hi_37, maskDestinationResult_hi_hi_lo_37};
  wire [7:0]    maskDestinationResult_hi_166 = {maskDestinationResult_hi_hi_38, maskDestinationResult_hi_lo_38};
  wire [1:0]    maskDestinationResult_lo_lo_lo_38 = {sourceDataVec_1[13], sourceDataVec_0[13]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_38 = {sourceDataVec_3[13], sourceDataVec_2[13]};
  wire [3:0]    maskDestinationResult_lo_lo_39 = {maskDestinationResult_lo_lo_hi_38, maskDestinationResult_lo_lo_lo_38};
  wire [1:0]    maskDestinationResult_lo_hi_lo_38 = {sourceDataVec_5[13], sourceDataVec_4[13]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_38 = {sourceDataVec_7[13], sourceDataVec_6[13]};
  wire [3:0]    maskDestinationResult_lo_hi_39 = {maskDestinationResult_lo_hi_hi_38, maskDestinationResult_lo_hi_lo_38};
  wire [7:0]    maskDestinationResult_lo_167 = {maskDestinationResult_lo_hi_39, maskDestinationResult_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_lo_lo_38 = {sourceDataVec_9[13], sourceDataVec_8[13]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_38 = {sourceDataVec_11[13], sourceDataVec_10[13]};
  wire [3:0]    maskDestinationResult_hi_lo_39 = {maskDestinationResult_hi_lo_hi_38, maskDestinationResult_hi_lo_lo_38};
  wire [1:0]    maskDestinationResult_hi_hi_lo_38 = {sourceDataVec_13[13], sourceDataVec_12[13]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_38 = {sourceDataVec_15[13], sourceDataVec_14[13]};
  wire [3:0]    maskDestinationResult_hi_hi_39 = {maskDestinationResult_hi_hi_hi_38, maskDestinationResult_hi_hi_lo_38};
  wire [7:0]    maskDestinationResult_hi_167 = {maskDestinationResult_hi_hi_39, maskDestinationResult_hi_lo_39};
  wire [1:0]    maskDestinationResult_lo_lo_lo_39 = {sourceDataVec_1[14], sourceDataVec_0[14]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_39 = {sourceDataVec_3[14], sourceDataVec_2[14]};
  wire [3:0]    maskDestinationResult_lo_lo_40 = {maskDestinationResult_lo_lo_hi_39, maskDestinationResult_lo_lo_lo_39};
  wire [1:0]    maskDestinationResult_lo_hi_lo_39 = {sourceDataVec_5[14], sourceDataVec_4[14]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_39 = {sourceDataVec_7[14], sourceDataVec_6[14]};
  wire [3:0]    maskDestinationResult_lo_hi_40 = {maskDestinationResult_lo_hi_hi_39, maskDestinationResult_lo_hi_lo_39};
  wire [7:0]    maskDestinationResult_lo_168 = {maskDestinationResult_lo_hi_40, maskDestinationResult_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_lo_lo_39 = {sourceDataVec_9[14], sourceDataVec_8[14]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_39 = {sourceDataVec_11[14], sourceDataVec_10[14]};
  wire [3:0]    maskDestinationResult_hi_lo_40 = {maskDestinationResult_hi_lo_hi_39, maskDestinationResult_hi_lo_lo_39};
  wire [1:0]    maskDestinationResult_hi_hi_lo_39 = {sourceDataVec_13[14], sourceDataVec_12[14]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_39 = {sourceDataVec_15[14], sourceDataVec_14[14]};
  wire [3:0]    maskDestinationResult_hi_hi_40 = {maskDestinationResult_hi_hi_hi_39, maskDestinationResult_hi_hi_lo_39};
  wire [7:0]    maskDestinationResult_hi_168 = {maskDestinationResult_hi_hi_40, maskDestinationResult_hi_lo_40};
  wire [1:0]    maskDestinationResult_lo_lo_lo_40 = {sourceDataVec_1[15], sourceDataVec_0[15]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_40 = {sourceDataVec_3[15], sourceDataVec_2[15]};
  wire [3:0]    maskDestinationResult_lo_lo_41 = {maskDestinationResult_lo_lo_hi_40, maskDestinationResult_lo_lo_lo_40};
  wire [1:0]    maskDestinationResult_lo_hi_lo_40 = {sourceDataVec_5[15], sourceDataVec_4[15]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_40 = {sourceDataVec_7[15], sourceDataVec_6[15]};
  wire [3:0]    maskDestinationResult_lo_hi_41 = {maskDestinationResult_lo_hi_hi_40, maskDestinationResult_lo_hi_lo_40};
  wire [7:0]    maskDestinationResult_lo_169 = {maskDestinationResult_lo_hi_41, maskDestinationResult_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_lo_lo_40 = {sourceDataVec_9[15], sourceDataVec_8[15]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_40 = {sourceDataVec_11[15], sourceDataVec_10[15]};
  wire [3:0]    maskDestinationResult_hi_lo_41 = {maskDestinationResult_hi_lo_hi_40, maskDestinationResult_hi_lo_lo_40};
  wire [1:0]    maskDestinationResult_hi_hi_lo_40 = {sourceDataVec_13[15], sourceDataVec_12[15]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_40 = {sourceDataVec_15[15], sourceDataVec_14[15]};
  wire [3:0]    maskDestinationResult_hi_hi_41 = {maskDestinationResult_hi_hi_hi_40, maskDestinationResult_hi_hi_lo_40};
  wire [7:0]    maskDestinationResult_hi_169 = {maskDestinationResult_hi_hi_41, maskDestinationResult_hi_lo_41};
  wire [1:0]    maskDestinationResult_lo_lo_lo_41 = {sourceDataVec_1[16], sourceDataVec_0[16]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_41 = {sourceDataVec_3[16], sourceDataVec_2[16]};
  wire [3:0]    maskDestinationResult_lo_lo_42 = {maskDestinationResult_lo_lo_hi_41, maskDestinationResult_lo_lo_lo_41};
  wire [1:0]    maskDestinationResult_lo_hi_lo_41 = {sourceDataVec_5[16], sourceDataVec_4[16]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_41 = {sourceDataVec_7[16], sourceDataVec_6[16]};
  wire [3:0]    maskDestinationResult_lo_hi_42 = {maskDestinationResult_lo_hi_hi_41, maskDestinationResult_lo_hi_lo_41};
  wire [7:0]    maskDestinationResult_lo_170 = {maskDestinationResult_lo_hi_42, maskDestinationResult_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_lo_lo_41 = {sourceDataVec_9[16], sourceDataVec_8[16]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_41 = {sourceDataVec_11[16], sourceDataVec_10[16]};
  wire [3:0]    maskDestinationResult_hi_lo_42 = {maskDestinationResult_hi_lo_hi_41, maskDestinationResult_hi_lo_lo_41};
  wire [1:0]    maskDestinationResult_hi_hi_lo_41 = {sourceDataVec_13[16], sourceDataVec_12[16]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_41 = {sourceDataVec_15[16], sourceDataVec_14[16]};
  wire [3:0]    maskDestinationResult_hi_hi_42 = {maskDestinationResult_hi_hi_hi_41, maskDestinationResult_hi_hi_lo_41};
  wire [7:0]    maskDestinationResult_hi_170 = {maskDestinationResult_hi_hi_42, maskDestinationResult_hi_lo_42};
  wire [1:0]    maskDestinationResult_lo_lo_lo_42 = {sourceDataVec_1[17], sourceDataVec_0[17]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_42 = {sourceDataVec_3[17], sourceDataVec_2[17]};
  wire [3:0]    maskDestinationResult_lo_lo_43 = {maskDestinationResult_lo_lo_hi_42, maskDestinationResult_lo_lo_lo_42};
  wire [1:0]    maskDestinationResult_lo_hi_lo_42 = {sourceDataVec_5[17], sourceDataVec_4[17]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_42 = {sourceDataVec_7[17], sourceDataVec_6[17]};
  wire [3:0]    maskDestinationResult_lo_hi_43 = {maskDestinationResult_lo_hi_hi_42, maskDestinationResult_lo_hi_lo_42};
  wire [7:0]    maskDestinationResult_lo_171 = {maskDestinationResult_lo_hi_43, maskDestinationResult_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_lo_lo_42 = {sourceDataVec_9[17], sourceDataVec_8[17]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_42 = {sourceDataVec_11[17], sourceDataVec_10[17]};
  wire [3:0]    maskDestinationResult_hi_lo_43 = {maskDestinationResult_hi_lo_hi_42, maskDestinationResult_hi_lo_lo_42};
  wire [1:0]    maskDestinationResult_hi_hi_lo_42 = {sourceDataVec_13[17], sourceDataVec_12[17]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_42 = {sourceDataVec_15[17], sourceDataVec_14[17]};
  wire [3:0]    maskDestinationResult_hi_hi_43 = {maskDestinationResult_hi_hi_hi_42, maskDestinationResult_hi_hi_lo_42};
  wire [7:0]    maskDestinationResult_hi_171 = {maskDestinationResult_hi_hi_43, maskDestinationResult_hi_lo_43};
  wire [1:0]    maskDestinationResult_lo_lo_lo_43 = {sourceDataVec_1[18], sourceDataVec_0[18]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_43 = {sourceDataVec_3[18], sourceDataVec_2[18]};
  wire [3:0]    maskDestinationResult_lo_lo_44 = {maskDestinationResult_lo_lo_hi_43, maskDestinationResult_lo_lo_lo_43};
  wire [1:0]    maskDestinationResult_lo_hi_lo_43 = {sourceDataVec_5[18], sourceDataVec_4[18]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_43 = {sourceDataVec_7[18], sourceDataVec_6[18]};
  wire [3:0]    maskDestinationResult_lo_hi_44 = {maskDestinationResult_lo_hi_hi_43, maskDestinationResult_lo_hi_lo_43};
  wire [7:0]    maskDestinationResult_lo_172 = {maskDestinationResult_lo_hi_44, maskDestinationResult_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_lo_lo_43 = {sourceDataVec_9[18], sourceDataVec_8[18]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_43 = {sourceDataVec_11[18], sourceDataVec_10[18]};
  wire [3:0]    maskDestinationResult_hi_lo_44 = {maskDestinationResult_hi_lo_hi_43, maskDestinationResult_hi_lo_lo_43};
  wire [1:0]    maskDestinationResult_hi_hi_lo_43 = {sourceDataVec_13[18], sourceDataVec_12[18]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_43 = {sourceDataVec_15[18], sourceDataVec_14[18]};
  wire [3:0]    maskDestinationResult_hi_hi_44 = {maskDestinationResult_hi_hi_hi_43, maskDestinationResult_hi_hi_lo_43};
  wire [7:0]    maskDestinationResult_hi_172 = {maskDestinationResult_hi_hi_44, maskDestinationResult_hi_lo_44};
  wire [1:0]    maskDestinationResult_lo_lo_lo_44 = {sourceDataVec_1[19], sourceDataVec_0[19]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_44 = {sourceDataVec_3[19], sourceDataVec_2[19]};
  wire [3:0]    maskDestinationResult_lo_lo_45 = {maskDestinationResult_lo_lo_hi_44, maskDestinationResult_lo_lo_lo_44};
  wire [1:0]    maskDestinationResult_lo_hi_lo_44 = {sourceDataVec_5[19], sourceDataVec_4[19]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_44 = {sourceDataVec_7[19], sourceDataVec_6[19]};
  wire [3:0]    maskDestinationResult_lo_hi_45 = {maskDestinationResult_lo_hi_hi_44, maskDestinationResult_lo_hi_lo_44};
  wire [7:0]    maskDestinationResult_lo_173 = {maskDestinationResult_lo_hi_45, maskDestinationResult_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_lo_lo_44 = {sourceDataVec_9[19], sourceDataVec_8[19]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_44 = {sourceDataVec_11[19], sourceDataVec_10[19]};
  wire [3:0]    maskDestinationResult_hi_lo_45 = {maskDestinationResult_hi_lo_hi_44, maskDestinationResult_hi_lo_lo_44};
  wire [1:0]    maskDestinationResult_hi_hi_lo_44 = {sourceDataVec_13[19], sourceDataVec_12[19]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_44 = {sourceDataVec_15[19], sourceDataVec_14[19]};
  wire [3:0]    maskDestinationResult_hi_hi_45 = {maskDestinationResult_hi_hi_hi_44, maskDestinationResult_hi_hi_lo_44};
  wire [7:0]    maskDestinationResult_hi_173 = {maskDestinationResult_hi_hi_45, maskDestinationResult_hi_lo_45};
  wire [1:0]    maskDestinationResult_lo_lo_lo_45 = {sourceDataVec_1[20], sourceDataVec_0[20]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_45 = {sourceDataVec_3[20], sourceDataVec_2[20]};
  wire [3:0]    maskDestinationResult_lo_lo_46 = {maskDestinationResult_lo_lo_hi_45, maskDestinationResult_lo_lo_lo_45};
  wire [1:0]    maskDestinationResult_lo_hi_lo_45 = {sourceDataVec_5[20], sourceDataVec_4[20]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_45 = {sourceDataVec_7[20], sourceDataVec_6[20]};
  wire [3:0]    maskDestinationResult_lo_hi_46 = {maskDestinationResult_lo_hi_hi_45, maskDestinationResult_lo_hi_lo_45};
  wire [7:0]    maskDestinationResult_lo_174 = {maskDestinationResult_lo_hi_46, maskDestinationResult_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_lo_lo_45 = {sourceDataVec_9[20], sourceDataVec_8[20]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_45 = {sourceDataVec_11[20], sourceDataVec_10[20]};
  wire [3:0]    maskDestinationResult_hi_lo_46 = {maskDestinationResult_hi_lo_hi_45, maskDestinationResult_hi_lo_lo_45};
  wire [1:0]    maskDestinationResult_hi_hi_lo_45 = {sourceDataVec_13[20], sourceDataVec_12[20]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_45 = {sourceDataVec_15[20], sourceDataVec_14[20]};
  wire [3:0]    maskDestinationResult_hi_hi_46 = {maskDestinationResult_hi_hi_hi_45, maskDestinationResult_hi_hi_lo_45};
  wire [7:0]    maskDestinationResult_hi_174 = {maskDestinationResult_hi_hi_46, maskDestinationResult_hi_lo_46};
  wire [1:0]    maskDestinationResult_lo_lo_lo_46 = {sourceDataVec_1[21], sourceDataVec_0[21]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_46 = {sourceDataVec_3[21], sourceDataVec_2[21]};
  wire [3:0]    maskDestinationResult_lo_lo_47 = {maskDestinationResult_lo_lo_hi_46, maskDestinationResult_lo_lo_lo_46};
  wire [1:0]    maskDestinationResult_lo_hi_lo_46 = {sourceDataVec_5[21], sourceDataVec_4[21]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_46 = {sourceDataVec_7[21], sourceDataVec_6[21]};
  wire [3:0]    maskDestinationResult_lo_hi_47 = {maskDestinationResult_lo_hi_hi_46, maskDestinationResult_lo_hi_lo_46};
  wire [7:0]    maskDestinationResult_lo_175 = {maskDestinationResult_lo_hi_47, maskDestinationResult_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_lo_lo_46 = {sourceDataVec_9[21], sourceDataVec_8[21]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_46 = {sourceDataVec_11[21], sourceDataVec_10[21]};
  wire [3:0]    maskDestinationResult_hi_lo_47 = {maskDestinationResult_hi_lo_hi_46, maskDestinationResult_hi_lo_lo_46};
  wire [1:0]    maskDestinationResult_hi_hi_lo_46 = {sourceDataVec_13[21], sourceDataVec_12[21]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_46 = {sourceDataVec_15[21], sourceDataVec_14[21]};
  wire [3:0]    maskDestinationResult_hi_hi_47 = {maskDestinationResult_hi_hi_hi_46, maskDestinationResult_hi_hi_lo_46};
  wire [7:0]    maskDestinationResult_hi_175 = {maskDestinationResult_hi_hi_47, maskDestinationResult_hi_lo_47};
  wire [1:0]    maskDestinationResult_lo_lo_lo_47 = {sourceDataVec_1[22], sourceDataVec_0[22]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_47 = {sourceDataVec_3[22], sourceDataVec_2[22]};
  wire [3:0]    maskDestinationResult_lo_lo_48 = {maskDestinationResult_lo_lo_hi_47, maskDestinationResult_lo_lo_lo_47};
  wire [1:0]    maskDestinationResult_lo_hi_lo_47 = {sourceDataVec_5[22], sourceDataVec_4[22]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_47 = {sourceDataVec_7[22], sourceDataVec_6[22]};
  wire [3:0]    maskDestinationResult_lo_hi_48 = {maskDestinationResult_lo_hi_hi_47, maskDestinationResult_lo_hi_lo_47};
  wire [7:0]    maskDestinationResult_lo_176 = {maskDestinationResult_lo_hi_48, maskDestinationResult_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_lo_lo_47 = {sourceDataVec_9[22], sourceDataVec_8[22]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_47 = {sourceDataVec_11[22], sourceDataVec_10[22]};
  wire [3:0]    maskDestinationResult_hi_lo_48 = {maskDestinationResult_hi_lo_hi_47, maskDestinationResult_hi_lo_lo_47};
  wire [1:0]    maskDestinationResult_hi_hi_lo_47 = {sourceDataVec_13[22], sourceDataVec_12[22]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_47 = {sourceDataVec_15[22], sourceDataVec_14[22]};
  wire [3:0]    maskDestinationResult_hi_hi_48 = {maskDestinationResult_hi_hi_hi_47, maskDestinationResult_hi_hi_lo_47};
  wire [7:0]    maskDestinationResult_hi_176 = {maskDestinationResult_hi_hi_48, maskDestinationResult_hi_lo_48};
  wire [1:0]    maskDestinationResult_lo_lo_lo_48 = {sourceDataVec_1[23], sourceDataVec_0[23]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_48 = {sourceDataVec_3[23], sourceDataVec_2[23]};
  wire [3:0]    maskDestinationResult_lo_lo_49 = {maskDestinationResult_lo_lo_hi_48, maskDestinationResult_lo_lo_lo_48};
  wire [1:0]    maskDestinationResult_lo_hi_lo_48 = {sourceDataVec_5[23], sourceDataVec_4[23]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_48 = {sourceDataVec_7[23], sourceDataVec_6[23]};
  wire [3:0]    maskDestinationResult_lo_hi_49 = {maskDestinationResult_lo_hi_hi_48, maskDestinationResult_lo_hi_lo_48};
  wire [7:0]    maskDestinationResult_lo_177 = {maskDestinationResult_lo_hi_49, maskDestinationResult_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_lo_lo_48 = {sourceDataVec_9[23], sourceDataVec_8[23]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_48 = {sourceDataVec_11[23], sourceDataVec_10[23]};
  wire [3:0]    maskDestinationResult_hi_lo_49 = {maskDestinationResult_hi_lo_hi_48, maskDestinationResult_hi_lo_lo_48};
  wire [1:0]    maskDestinationResult_hi_hi_lo_48 = {sourceDataVec_13[23], sourceDataVec_12[23]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_48 = {sourceDataVec_15[23], sourceDataVec_14[23]};
  wire [3:0]    maskDestinationResult_hi_hi_49 = {maskDestinationResult_hi_hi_hi_48, maskDestinationResult_hi_hi_lo_48};
  wire [7:0]    maskDestinationResult_hi_177 = {maskDestinationResult_hi_hi_49, maskDestinationResult_hi_lo_49};
  wire [1:0]    maskDestinationResult_lo_lo_lo_49 = {sourceDataVec_1[24], sourceDataVec_0[24]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_49 = {sourceDataVec_3[24], sourceDataVec_2[24]};
  wire [3:0]    maskDestinationResult_lo_lo_50 = {maskDestinationResult_lo_lo_hi_49, maskDestinationResult_lo_lo_lo_49};
  wire [1:0]    maskDestinationResult_lo_hi_lo_49 = {sourceDataVec_5[24], sourceDataVec_4[24]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_49 = {sourceDataVec_7[24], sourceDataVec_6[24]};
  wire [3:0]    maskDestinationResult_lo_hi_50 = {maskDestinationResult_lo_hi_hi_49, maskDestinationResult_lo_hi_lo_49};
  wire [7:0]    maskDestinationResult_lo_178 = {maskDestinationResult_lo_hi_50, maskDestinationResult_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_lo_lo_49 = {sourceDataVec_9[24], sourceDataVec_8[24]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_49 = {sourceDataVec_11[24], sourceDataVec_10[24]};
  wire [3:0]    maskDestinationResult_hi_lo_50 = {maskDestinationResult_hi_lo_hi_49, maskDestinationResult_hi_lo_lo_49};
  wire [1:0]    maskDestinationResult_hi_hi_lo_49 = {sourceDataVec_13[24], sourceDataVec_12[24]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_49 = {sourceDataVec_15[24], sourceDataVec_14[24]};
  wire [3:0]    maskDestinationResult_hi_hi_50 = {maskDestinationResult_hi_hi_hi_49, maskDestinationResult_hi_hi_lo_49};
  wire [7:0]    maskDestinationResult_hi_178 = {maskDestinationResult_hi_hi_50, maskDestinationResult_hi_lo_50};
  wire [1:0]    maskDestinationResult_lo_lo_lo_50 = {sourceDataVec_1[25], sourceDataVec_0[25]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_50 = {sourceDataVec_3[25], sourceDataVec_2[25]};
  wire [3:0]    maskDestinationResult_lo_lo_51 = {maskDestinationResult_lo_lo_hi_50, maskDestinationResult_lo_lo_lo_50};
  wire [1:0]    maskDestinationResult_lo_hi_lo_50 = {sourceDataVec_5[25], sourceDataVec_4[25]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_50 = {sourceDataVec_7[25], sourceDataVec_6[25]};
  wire [3:0]    maskDestinationResult_lo_hi_51 = {maskDestinationResult_lo_hi_hi_50, maskDestinationResult_lo_hi_lo_50};
  wire [7:0]    maskDestinationResult_lo_179 = {maskDestinationResult_lo_hi_51, maskDestinationResult_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_lo_lo_50 = {sourceDataVec_9[25], sourceDataVec_8[25]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_50 = {sourceDataVec_11[25], sourceDataVec_10[25]};
  wire [3:0]    maskDestinationResult_hi_lo_51 = {maskDestinationResult_hi_lo_hi_50, maskDestinationResult_hi_lo_lo_50};
  wire [1:0]    maskDestinationResult_hi_hi_lo_50 = {sourceDataVec_13[25], sourceDataVec_12[25]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_50 = {sourceDataVec_15[25], sourceDataVec_14[25]};
  wire [3:0]    maskDestinationResult_hi_hi_51 = {maskDestinationResult_hi_hi_hi_50, maskDestinationResult_hi_hi_lo_50};
  wire [7:0]    maskDestinationResult_hi_179 = {maskDestinationResult_hi_hi_51, maskDestinationResult_hi_lo_51};
  wire [1:0]    maskDestinationResult_lo_lo_lo_51 = {sourceDataVec_1[26], sourceDataVec_0[26]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_51 = {sourceDataVec_3[26], sourceDataVec_2[26]};
  wire [3:0]    maskDestinationResult_lo_lo_52 = {maskDestinationResult_lo_lo_hi_51, maskDestinationResult_lo_lo_lo_51};
  wire [1:0]    maskDestinationResult_lo_hi_lo_51 = {sourceDataVec_5[26], sourceDataVec_4[26]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_51 = {sourceDataVec_7[26], sourceDataVec_6[26]};
  wire [3:0]    maskDestinationResult_lo_hi_52 = {maskDestinationResult_lo_hi_hi_51, maskDestinationResult_lo_hi_lo_51};
  wire [7:0]    maskDestinationResult_lo_180 = {maskDestinationResult_lo_hi_52, maskDestinationResult_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_lo_lo_51 = {sourceDataVec_9[26], sourceDataVec_8[26]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_51 = {sourceDataVec_11[26], sourceDataVec_10[26]};
  wire [3:0]    maskDestinationResult_hi_lo_52 = {maskDestinationResult_hi_lo_hi_51, maskDestinationResult_hi_lo_lo_51};
  wire [1:0]    maskDestinationResult_hi_hi_lo_51 = {sourceDataVec_13[26], sourceDataVec_12[26]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_51 = {sourceDataVec_15[26], sourceDataVec_14[26]};
  wire [3:0]    maskDestinationResult_hi_hi_52 = {maskDestinationResult_hi_hi_hi_51, maskDestinationResult_hi_hi_lo_51};
  wire [7:0]    maskDestinationResult_hi_180 = {maskDestinationResult_hi_hi_52, maskDestinationResult_hi_lo_52};
  wire [1:0]    maskDestinationResult_lo_lo_lo_52 = {sourceDataVec_1[27], sourceDataVec_0[27]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_52 = {sourceDataVec_3[27], sourceDataVec_2[27]};
  wire [3:0]    maskDestinationResult_lo_lo_53 = {maskDestinationResult_lo_lo_hi_52, maskDestinationResult_lo_lo_lo_52};
  wire [1:0]    maskDestinationResult_lo_hi_lo_52 = {sourceDataVec_5[27], sourceDataVec_4[27]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_52 = {sourceDataVec_7[27], sourceDataVec_6[27]};
  wire [3:0]    maskDestinationResult_lo_hi_53 = {maskDestinationResult_lo_hi_hi_52, maskDestinationResult_lo_hi_lo_52};
  wire [7:0]    maskDestinationResult_lo_181 = {maskDestinationResult_lo_hi_53, maskDestinationResult_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_lo_lo_52 = {sourceDataVec_9[27], sourceDataVec_8[27]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_52 = {sourceDataVec_11[27], sourceDataVec_10[27]};
  wire [3:0]    maskDestinationResult_hi_lo_53 = {maskDestinationResult_hi_lo_hi_52, maskDestinationResult_hi_lo_lo_52};
  wire [1:0]    maskDestinationResult_hi_hi_lo_52 = {sourceDataVec_13[27], sourceDataVec_12[27]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_52 = {sourceDataVec_15[27], sourceDataVec_14[27]};
  wire [3:0]    maskDestinationResult_hi_hi_53 = {maskDestinationResult_hi_hi_hi_52, maskDestinationResult_hi_hi_lo_52};
  wire [7:0]    maskDestinationResult_hi_181 = {maskDestinationResult_hi_hi_53, maskDestinationResult_hi_lo_53};
  wire [1:0]    maskDestinationResult_lo_lo_lo_53 = {sourceDataVec_1[28], sourceDataVec_0[28]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_53 = {sourceDataVec_3[28], sourceDataVec_2[28]};
  wire [3:0]    maskDestinationResult_lo_lo_54 = {maskDestinationResult_lo_lo_hi_53, maskDestinationResult_lo_lo_lo_53};
  wire [1:0]    maskDestinationResult_lo_hi_lo_53 = {sourceDataVec_5[28], sourceDataVec_4[28]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_53 = {sourceDataVec_7[28], sourceDataVec_6[28]};
  wire [3:0]    maskDestinationResult_lo_hi_54 = {maskDestinationResult_lo_hi_hi_53, maskDestinationResult_lo_hi_lo_53};
  wire [7:0]    maskDestinationResult_lo_182 = {maskDestinationResult_lo_hi_54, maskDestinationResult_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_lo_lo_53 = {sourceDataVec_9[28], sourceDataVec_8[28]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_53 = {sourceDataVec_11[28], sourceDataVec_10[28]};
  wire [3:0]    maskDestinationResult_hi_lo_54 = {maskDestinationResult_hi_lo_hi_53, maskDestinationResult_hi_lo_lo_53};
  wire [1:0]    maskDestinationResult_hi_hi_lo_53 = {sourceDataVec_13[28], sourceDataVec_12[28]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_53 = {sourceDataVec_15[28], sourceDataVec_14[28]};
  wire [3:0]    maskDestinationResult_hi_hi_54 = {maskDestinationResult_hi_hi_hi_53, maskDestinationResult_hi_hi_lo_53};
  wire [7:0]    maskDestinationResult_hi_182 = {maskDestinationResult_hi_hi_54, maskDestinationResult_hi_lo_54};
  wire [1:0]    maskDestinationResult_lo_lo_lo_54 = {sourceDataVec_1[29], sourceDataVec_0[29]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_54 = {sourceDataVec_3[29], sourceDataVec_2[29]};
  wire [3:0]    maskDestinationResult_lo_lo_55 = {maskDestinationResult_lo_lo_hi_54, maskDestinationResult_lo_lo_lo_54};
  wire [1:0]    maskDestinationResult_lo_hi_lo_54 = {sourceDataVec_5[29], sourceDataVec_4[29]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_54 = {sourceDataVec_7[29], sourceDataVec_6[29]};
  wire [3:0]    maskDestinationResult_lo_hi_55 = {maskDestinationResult_lo_hi_hi_54, maskDestinationResult_lo_hi_lo_54};
  wire [7:0]    maskDestinationResult_lo_183 = {maskDestinationResult_lo_hi_55, maskDestinationResult_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_lo_lo_54 = {sourceDataVec_9[29], sourceDataVec_8[29]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_54 = {sourceDataVec_11[29], sourceDataVec_10[29]};
  wire [3:0]    maskDestinationResult_hi_lo_55 = {maskDestinationResult_hi_lo_hi_54, maskDestinationResult_hi_lo_lo_54};
  wire [1:0]    maskDestinationResult_hi_hi_lo_54 = {sourceDataVec_13[29], sourceDataVec_12[29]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_54 = {sourceDataVec_15[29], sourceDataVec_14[29]};
  wire [3:0]    maskDestinationResult_hi_hi_55 = {maskDestinationResult_hi_hi_hi_54, maskDestinationResult_hi_hi_lo_54};
  wire [7:0]    maskDestinationResult_hi_183 = {maskDestinationResult_hi_hi_55, maskDestinationResult_hi_lo_55};
  wire [1:0]    maskDestinationResult_lo_lo_lo_55 = {sourceDataVec_1[30], sourceDataVec_0[30]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_55 = {sourceDataVec_3[30], sourceDataVec_2[30]};
  wire [3:0]    maskDestinationResult_lo_lo_56 = {maskDestinationResult_lo_lo_hi_55, maskDestinationResult_lo_lo_lo_55};
  wire [1:0]    maskDestinationResult_lo_hi_lo_55 = {sourceDataVec_5[30], sourceDataVec_4[30]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_55 = {sourceDataVec_7[30], sourceDataVec_6[30]};
  wire [3:0]    maskDestinationResult_lo_hi_56 = {maskDestinationResult_lo_hi_hi_55, maskDestinationResult_lo_hi_lo_55};
  wire [7:0]    maskDestinationResult_lo_184 = {maskDestinationResult_lo_hi_56, maskDestinationResult_lo_lo_56};
  wire [1:0]    maskDestinationResult_hi_lo_lo_55 = {sourceDataVec_9[30], sourceDataVec_8[30]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_55 = {sourceDataVec_11[30], sourceDataVec_10[30]};
  wire [3:0]    maskDestinationResult_hi_lo_56 = {maskDestinationResult_hi_lo_hi_55, maskDestinationResult_hi_lo_lo_55};
  wire [1:0]    maskDestinationResult_hi_hi_lo_55 = {sourceDataVec_13[30], sourceDataVec_12[30]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_55 = {sourceDataVec_15[30], sourceDataVec_14[30]};
  wire [3:0]    maskDestinationResult_hi_hi_56 = {maskDestinationResult_hi_hi_hi_55, maskDestinationResult_hi_hi_lo_55};
  wire [7:0]    maskDestinationResult_hi_184 = {maskDestinationResult_hi_hi_56, maskDestinationResult_hi_lo_56};
  wire [1:0]    maskDestinationResult_lo_lo_lo_56 = {sourceDataVec_1[31], sourceDataVec_0[31]};
  wire [1:0]    maskDestinationResult_lo_lo_hi_56 = {sourceDataVec_3[31], sourceDataVec_2[31]};
  wire [3:0]    maskDestinationResult_lo_lo_57 = {maskDestinationResult_lo_lo_hi_56, maskDestinationResult_lo_lo_lo_56};
  wire [1:0]    maskDestinationResult_lo_hi_lo_56 = {sourceDataVec_5[31], sourceDataVec_4[31]};
  wire [1:0]    maskDestinationResult_lo_hi_hi_56 = {sourceDataVec_7[31], sourceDataVec_6[31]};
  wire [3:0]    maskDestinationResult_lo_hi_57 = {maskDestinationResult_lo_hi_hi_56, maskDestinationResult_lo_hi_lo_56};
  wire [7:0]    maskDestinationResult_lo_185 = {maskDestinationResult_lo_hi_57, maskDestinationResult_lo_lo_57};
  wire [1:0]    maskDestinationResult_hi_lo_lo_56 = {sourceDataVec_9[31], sourceDataVec_8[31]};
  wire [1:0]    maskDestinationResult_hi_lo_hi_56 = {sourceDataVec_11[31], sourceDataVec_10[31]};
  wire [3:0]    maskDestinationResult_hi_lo_57 = {maskDestinationResult_hi_lo_hi_56, maskDestinationResult_hi_lo_lo_56};
  wire [1:0]    maskDestinationResult_hi_hi_lo_56 = {sourceDataVec_13[31], sourceDataVec_12[31]};
  wire [1:0]    maskDestinationResult_hi_hi_hi_56 = {sourceDataVec_15[31], sourceDataVec_14[31]};
  wire [3:0]    maskDestinationResult_hi_hi_57 = {maskDestinationResult_hi_hi_hi_56, maskDestinationResult_hi_hi_lo_56};
  wire [7:0]    maskDestinationResult_hi_185 = {maskDestinationResult_hi_hi_57, maskDestinationResult_hi_lo_57};
  wire [31:0]   maskDestinationResult_lo_lo_lo_lo = {maskDestinationResult_hi_155, maskDestinationResult_lo_155, maskDestinationResult_hi_154, maskDestinationResult_lo_154};
  wire [31:0]   maskDestinationResult_lo_lo_lo_hi = {maskDestinationResult_hi_157, maskDestinationResult_lo_157, maskDestinationResult_hi_156, maskDestinationResult_lo_156};
  wire [63:0]   maskDestinationResult_lo_lo_lo_57 = {maskDestinationResult_lo_lo_lo_hi, maskDestinationResult_lo_lo_lo_lo};
  wire [31:0]   maskDestinationResult_lo_lo_hi_lo = {maskDestinationResult_hi_159, maskDestinationResult_lo_159, maskDestinationResult_hi_158, maskDestinationResult_lo_158};
  wire [31:0]   maskDestinationResult_lo_lo_hi_hi = {maskDestinationResult_hi_161, maskDestinationResult_lo_161, maskDestinationResult_hi_160, maskDestinationResult_lo_160};
  wire [63:0]   maskDestinationResult_lo_lo_hi_57 = {maskDestinationResult_lo_lo_hi_hi, maskDestinationResult_lo_lo_hi_lo};
  wire [127:0]  maskDestinationResult_lo_lo_58 = {maskDestinationResult_lo_lo_hi_57, maskDestinationResult_lo_lo_lo_57};
  wire [31:0]   maskDestinationResult_lo_hi_lo_lo = {maskDestinationResult_hi_163, maskDestinationResult_lo_163, maskDestinationResult_hi_162, maskDestinationResult_lo_162};
  wire [31:0]   maskDestinationResult_lo_hi_lo_hi = {maskDestinationResult_hi_165, maskDestinationResult_lo_165, maskDestinationResult_hi_164, maskDestinationResult_lo_164};
  wire [63:0]   maskDestinationResult_lo_hi_lo_57 = {maskDestinationResult_lo_hi_lo_hi, maskDestinationResult_lo_hi_lo_lo};
  wire [31:0]   maskDestinationResult_lo_hi_hi_lo = {maskDestinationResult_hi_167, maskDestinationResult_lo_167, maskDestinationResult_hi_166, maskDestinationResult_lo_166};
  wire [31:0]   maskDestinationResult_lo_hi_hi_hi = {maskDestinationResult_hi_169, maskDestinationResult_lo_169, maskDestinationResult_hi_168, maskDestinationResult_lo_168};
  wire [63:0]   maskDestinationResult_lo_hi_hi_57 = {maskDestinationResult_lo_hi_hi_hi, maskDestinationResult_lo_hi_hi_lo};
  wire [127:0]  maskDestinationResult_lo_hi_58 = {maskDestinationResult_lo_hi_hi_57, maskDestinationResult_lo_hi_lo_57};
  wire [255:0]  maskDestinationResult_lo_186 = {maskDestinationResult_lo_hi_58, maskDestinationResult_lo_lo_58};
  wire [31:0]   maskDestinationResult_hi_lo_lo_lo = {maskDestinationResult_hi_171, maskDestinationResult_lo_171, maskDestinationResult_hi_170, maskDestinationResult_lo_170};
  wire [31:0]   maskDestinationResult_hi_lo_lo_hi = {maskDestinationResult_hi_173, maskDestinationResult_lo_173, maskDestinationResult_hi_172, maskDestinationResult_lo_172};
  wire [63:0]   maskDestinationResult_hi_lo_lo_57 = {maskDestinationResult_hi_lo_lo_hi, maskDestinationResult_hi_lo_lo_lo};
  wire [31:0]   maskDestinationResult_hi_lo_hi_lo = {maskDestinationResult_hi_175, maskDestinationResult_lo_175, maskDestinationResult_hi_174, maskDestinationResult_lo_174};
  wire [31:0]   maskDestinationResult_hi_lo_hi_hi = {maskDestinationResult_hi_177, maskDestinationResult_lo_177, maskDestinationResult_hi_176, maskDestinationResult_lo_176};
  wire [63:0]   maskDestinationResult_hi_lo_hi_57 = {maskDestinationResult_hi_lo_hi_hi, maskDestinationResult_hi_lo_hi_lo};
  wire [127:0]  maskDestinationResult_hi_lo_58 = {maskDestinationResult_hi_lo_hi_57, maskDestinationResult_hi_lo_lo_57};
  wire [31:0]   maskDestinationResult_hi_hi_lo_lo = {maskDestinationResult_hi_179, maskDestinationResult_lo_179, maskDestinationResult_hi_178, maskDestinationResult_lo_178};
  wire [31:0]   maskDestinationResult_hi_hi_lo_hi = {maskDestinationResult_hi_181, maskDestinationResult_lo_181, maskDestinationResult_hi_180, maskDestinationResult_lo_180};
  wire [63:0]   maskDestinationResult_hi_hi_lo_57 = {maskDestinationResult_hi_hi_lo_hi, maskDestinationResult_hi_hi_lo_lo};
  wire [31:0]   maskDestinationResult_hi_hi_hi_lo = {maskDestinationResult_hi_183, maskDestinationResult_lo_183, maskDestinationResult_hi_182, maskDestinationResult_lo_182};
  wire [31:0]   maskDestinationResult_hi_hi_hi_hi = {maskDestinationResult_hi_185, maskDestinationResult_lo_185, maskDestinationResult_hi_184, maskDestinationResult_lo_184};
  wire [63:0]   maskDestinationResult_hi_hi_hi_57 = {maskDestinationResult_hi_hi_hi_hi, maskDestinationResult_hi_hi_hi_lo};
  wire [127:0]  maskDestinationResult_hi_hi_58 = {maskDestinationResult_hi_hi_hi_57, maskDestinationResult_hi_hi_lo_57};
  wire [255:0]  maskDestinationResult_hi_186 = {maskDestinationResult_hi_hi_58, maskDestinationResult_hi_lo_58};
  wire [511:0]  maskDestinationResult =
    (eew1H[0] ? {maskDestinationResult_hi_136, maskDestinationResult_lo_136} : 512'h0) | (eew1H[1] ? {maskDestinationResult_hi_153, maskDestinationResult_lo_153} : 512'h0)
    | (eew1H[2] ? {maskDestinationResult_hi_186, maskDestinationResult_lo_186} : 512'h0);
  wire          sign = in_uop[0];
  wire          extendRatio = in_uop[2];
  wire [3:0]    _source2_T_1 = 4'h1 << in_groupCounter[1:0];
  wire [1:0]    _source2_T_18 = 2'h1 << in_groupCounter[0];
  wire [255:0]  source2 =
    extendRatio
      ? {128'h0, (_source2_T_1[0] ? in_source2[127:0] : 128'h0) | (_source2_T_1[1] ? in_source2[255:128] : 128'h0) | (_source2_T_1[2] ? in_source2[383:256] : 128'h0) | (_source2_T_1[3] ? in_source2[511:384] : 128'h0)}
      : (_source2_T_18[0] ? in_source2[255:0] : 256'h0) | (_source2_T_18[1] ? in_source2[511:256] : 256'h0);
  wire [1:0]    _extendResult_T_489 = 2'h1 << extendRatio;
  wire [31:0]   extendResult_lo_lo_lo_lo = {{8{source2[15] & sign}}, source2[15:8], {8{source2[7] & sign}}, source2[7:0]};
  wire [31:0]   extendResult_lo_lo_lo_hi = {{8{source2[31] & sign}}, source2[31:24], {8{source2[23] & sign}}, source2[23:16]};
  wire [63:0]   extendResult_lo_lo_lo = {extendResult_lo_lo_lo_hi, extendResult_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_lo = {{8{source2[47] & sign}}, source2[47:40], {8{source2[39] & sign}}, source2[39:32]};
  wire [31:0]   extendResult_lo_lo_hi_hi = {{8{source2[63] & sign}}, source2[63:56], {8{source2[55] & sign}}, source2[55:48]};
  wire [63:0]   extendResult_lo_lo_hi = {extendResult_lo_lo_hi_hi, extendResult_lo_lo_hi_lo};
  wire [127:0]  extendResult_lo_lo = {extendResult_lo_lo_hi, extendResult_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_lo = {{8{source2[79] & sign}}, source2[79:72], {8{source2[71] & sign}}, source2[71:64]};
  wire [31:0]   extendResult_lo_hi_lo_hi = {{8{source2[95] & sign}}, source2[95:88], {8{source2[87] & sign}}, source2[87:80]};
  wire [63:0]   extendResult_lo_hi_lo = {extendResult_lo_hi_lo_hi, extendResult_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_lo = {{8{source2[111] & sign}}, source2[111:104], {8{source2[103] & sign}}, source2[103:96]};
  wire [31:0]   extendResult_lo_hi_hi_hi = {{8{source2[127] & sign}}, source2[127:120], {8{source2[119] & sign}}, source2[119:112]};
  wire [63:0]   extendResult_lo_hi_hi = {extendResult_lo_hi_hi_hi, extendResult_lo_hi_hi_lo};
  wire [127:0]  extendResult_lo_hi = {extendResult_lo_hi_hi, extendResult_lo_hi_lo};
  wire [255:0]  extendResult_lo = {extendResult_lo_hi, extendResult_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_lo = {{8{source2[143] & sign}}, source2[143:136], {8{source2[135] & sign}}, source2[135:128]};
  wire [31:0]   extendResult_hi_lo_lo_hi = {{8{source2[159] & sign}}, source2[159:152], {8{source2[151] & sign}}, source2[151:144]};
  wire [63:0]   extendResult_hi_lo_lo = {extendResult_hi_lo_lo_hi, extendResult_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_lo = {{8{source2[175] & sign}}, source2[175:168], {8{source2[167] & sign}}, source2[167:160]};
  wire [31:0]   extendResult_hi_lo_hi_hi = {{8{source2[191] & sign}}, source2[191:184], {8{source2[183] & sign}}, source2[183:176]};
  wire [63:0]   extendResult_hi_lo_hi = {extendResult_hi_lo_hi_hi, extendResult_hi_lo_hi_lo};
  wire [127:0]  extendResult_hi_lo = {extendResult_hi_lo_hi, extendResult_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_lo = {{8{source2[207] & sign}}, source2[207:200], {8{source2[199] & sign}}, source2[199:192]};
  wire [31:0]   extendResult_hi_hi_lo_hi = {{8{source2[223] & sign}}, source2[223:216], {8{source2[215] & sign}}, source2[215:208]};
  wire [63:0]   extendResult_hi_hi_lo = {extendResult_hi_hi_lo_hi, extendResult_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_lo = {{8{source2[239] & sign}}, source2[239:232], {8{source2[231] & sign}}, source2[231:224]};
  wire [31:0]   extendResult_hi_hi_hi_hi = {{8{source2[255] & sign}}, source2[255:248], {8{source2[247] & sign}}, source2[247:240]};
  wire [63:0]   extendResult_hi_hi_hi = {extendResult_hi_hi_hi_hi, extendResult_hi_hi_hi_lo};
  wire [127:0]  extendResult_hi_hi = {extendResult_hi_hi_hi, extendResult_hi_hi_lo};
  wire [255:0]  extendResult_hi = {extendResult_hi_hi, extendResult_hi_lo};
  wire [31:0]   extendResult_lo_lo_lo_lo_lo = {{12{source2[7] & sign}}, source2[7:4], {12{source2[3] & sign}}, source2[3:0]};
  wire [31:0]   extendResult_lo_lo_lo_lo_hi = {{12{source2[15] & sign}}, source2[15:12], {12{source2[11] & sign}}, source2[11:8]};
  wire [63:0]   extendResult_lo_lo_lo_lo_1 = {extendResult_lo_lo_lo_lo_hi, extendResult_lo_lo_lo_lo_lo};
  wire [31:0]   extendResult_lo_lo_lo_hi_lo = {{12{source2[23] & sign}}, source2[23:20], {12{source2[19] & sign}}, source2[19:16]};
  wire [31:0]   extendResult_lo_lo_lo_hi_hi = {{12{source2[31] & sign}}, source2[31:28], {12{source2[27] & sign}}, source2[27:24]};
  wire [63:0]   extendResult_lo_lo_lo_hi_1 = {extendResult_lo_lo_lo_hi_hi, extendResult_lo_lo_lo_hi_lo};
  wire [127:0]  extendResult_lo_lo_lo_1 = {extendResult_lo_lo_lo_hi_1, extendResult_lo_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_lo_hi_lo_lo = {{12{source2[39] & sign}}, source2[39:36], {12{source2[35] & sign}}, source2[35:32]};
  wire [31:0]   extendResult_lo_lo_hi_lo_hi = {{12{source2[47] & sign}}, source2[47:44], {12{source2[43] & sign}}, source2[43:40]};
  wire [63:0]   extendResult_lo_lo_hi_lo_1 = {extendResult_lo_lo_hi_lo_hi, extendResult_lo_lo_hi_lo_lo};
  wire [31:0]   extendResult_lo_lo_hi_hi_lo = {{12{source2[55] & sign}}, source2[55:52], {12{source2[51] & sign}}, source2[51:48]};
  wire [31:0]   extendResult_lo_lo_hi_hi_hi = {{12{source2[63] & sign}}, source2[63:60], {12{source2[59] & sign}}, source2[59:56]};
  wire [63:0]   extendResult_lo_lo_hi_hi_1 = {extendResult_lo_lo_hi_hi_hi, extendResult_lo_lo_hi_hi_lo};
  wire [127:0]  extendResult_lo_lo_hi_1 = {extendResult_lo_lo_hi_hi_1, extendResult_lo_lo_hi_lo_1};
  wire [255:0]  extendResult_lo_lo_1 = {extendResult_lo_lo_hi_1, extendResult_lo_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_lo_lo_lo = {{12{source2[71] & sign}}, source2[71:68], {12{source2[67] & sign}}, source2[67:64]};
  wire [31:0]   extendResult_lo_hi_lo_lo_hi = {{12{source2[79] & sign}}, source2[79:76], {12{source2[75] & sign}}, source2[75:72]};
  wire [63:0]   extendResult_lo_hi_lo_lo_1 = {extendResult_lo_hi_lo_lo_hi, extendResult_lo_hi_lo_lo_lo};
  wire [31:0]   extendResult_lo_hi_lo_hi_lo = {{12{source2[87] & sign}}, source2[87:84], {12{source2[83] & sign}}, source2[83:80]};
  wire [31:0]   extendResult_lo_hi_lo_hi_hi = {{12{source2[95] & sign}}, source2[95:92], {12{source2[91] & sign}}, source2[91:88]};
  wire [63:0]   extendResult_lo_hi_lo_hi_1 = {extendResult_lo_hi_lo_hi_hi, extendResult_lo_hi_lo_hi_lo};
  wire [127:0]  extendResult_lo_hi_lo_1 = {extendResult_lo_hi_lo_hi_1, extendResult_lo_hi_lo_lo_1};
  wire [31:0]   extendResult_lo_hi_hi_lo_lo = {{12{source2[103] & sign}}, source2[103:100], {12{source2[99] & sign}}, source2[99:96]};
  wire [31:0]   extendResult_lo_hi_hi_lo_hi = {{12{source2[111] & sign}}, source2[111:108], {12{source2[107] & sign}}, source2[107:104]};
  wire [63:0]   extendResult_lo_hi_hi_lo_1 = {extendResult_lo_hi_hi_lo_hi, extendResult_lo_hi_hi_lo_lo};
  wire [31:0]   extendResult_lo_hi_hi_hi_lo = {{12{source2[119] & sign}}, source2[119:116], {12{source2[115] & sign}}, source2[115:112]};
  wire [31:0]   extendResult_lo_hi_hi_hi_hi = {{12{source2[127] & sign}}, source2[127:124], {12{source2[123] & sign}}, source2[123:120]};
  wire [63:0]   extendResult_lo_hi_hi_hi_1 = {extendResult_lo_hi_hi_hi_hi, extendResult_lo_hi_hi_hi_lo};
  wire [127:0]  extendResult_lo_hi_hi_1 = {extendResult_lo_hi_hi_hi_1, extendResult_lo_hi_hi_lo_1};
  wire [255:0]  extendResult_lo_hi_1 = {extendResult_lo_hi_hi_1, extendResult_lo_hi_lo_1};
  wire [511:0]  extendResult_lo_1 = {extendResult_lo_hi_1, extendResult_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_lo_lo_lo = {{12{source2[135] & sign}}, source2[135:132], {12{source2[131] & sign}}, source2[131:128]};
  wire [31:0]   extendResult_hi_lo_lo_lo_hi = {{12{source2[143] & sign}}, source2[143:140], {12{source2[139] & sign}}, source2[139:136]};
  wire [63:0]   extendResult_hi_lo_lo_lo_1 = {extendResult_hi_lo_lo_lo_hi, extendResult_hi_lo_lo_lo_lo};
  wire [31:0]   extendResult_hi_lo_lo_hi_lo = {{12{source2[151] & sign}}, source2[151:148], {12{source2[147] & sign}}, source2[147:144]};
  wire [31:0]   extendResult_hi_lo_lo_hi_hi = {{12{source2[159] & sign}}, source2[159:156], {12{source2[155] & sign}}, source2[155:152]};
  wire [63:0]   extendResult_hi_lo_lo_hi_1 = {extendResult_hi_lo_lo_hi_hi, extendResult_hi_lo_lo_hi_lo};
  wire [127:0]  extendResult_hi_lo_lo_1 = {extendResult_hi_lo_lo_hi_1, extendResult_hi_lo_lo_lo_1};
  wire [31:0]   extendResult_hi_lo_hi_lo_lo = {{12{source2[167] & sign}}, source2[167:164], {12{source2[163] & sign}}, source2[163:160]};
  wire [31:0]   extendResult_hi_lo_hi_lo_hi = {{12{source2[175] & sign}}, source2[175:172], {12{source2[171] & sign}}, source2[171:168]};
  wire [63:0]   extendResult_hi_lo_hi_lo_1 = {extendResult_hi_lo_hi_lo_hi, extendResult_hi_lo_hi_lo_lo};
  wire [31:0]   extendResult_hi_lo_hi_hi_lo = {{12{source2[183] & sign}}, source2[183:180], {12{source2[179] & sign}}, source2[179:176]};
  wire [31:0]   extendResult_hi_lo_hi_hi_hi = {{12{source2[191] & sign}}, source2[191:188], {12{source2[187] & sign}}, source2[187:184]};
  wire [63:0]   extendResult_hi_lo_hi_hi_1 = {extendResult_hi_lo_hi_hi_hi, extendResult_hi_lo_hi_hi_lo};
  wire [127:0]  extendResult_hi_lo_hi_1 = {extendResult_hi_lo_hi_hi_1, extendResult_hi_lo_hi_lo_1};
  wire [255:0]  extendResult_hi_lo_1 = {extendResult_hi_lo_hi_1, extendResult_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_lo_lo_lo = {{12{source2[199] & sign}}, source2[199:196], {12{source2[195] & sign}}, source2[195:192]};
  wire [31:0]   extendResult_hi_hi_lo_lo_hi = {{12{source2[207] & sign}}, source2[207:204], {12{source2[203] & sign}}, source2[203:200]};
  wire [63:0]   extendResult_hi_hi_lo_lo_1 = {extendResult_hi_hi_lo_lo_hi, extendResult_hi_hi_lo_lo_lo};
  wire [31:0]   extendResult_hi_hi_lo_hi_lo = {{12{source2[215] & sign}}, source2[215:212], {12{source2[211] & sign}}, source2[211:208]};
  wire [31:0]   extendResult_hi_hi_lo_hi_hi = {{12{source2[223] & sign}}, source2[223:220], {12{source2[219] & sign}}, source2[219:216]};
  wire [63:0]   extendResult_hi_hi_lo_hi_1 = {extendResult_hi_hi_lo_hi_hi, extendResult_hi_hi_lo_hi_lo};
  wire [127:0]  extendResult_hi_hi_lo_1 = {extendResult_hi_hi_lo_hi_1, extendResult_hi_hi_lo_lo_1};
  wire [31:0]   extendResult_hi_hi_hi_lo_lo = {{12{source2[231] & sign}}, source2[231:228], {12{source2[227] & sign}}, source2[227:224]};
  wire [31:0]   extendResult_hi_hi_hi_lo_hi = {{12{source2[239] & sign}}, source2[239:236], {12{source2[235] & sign}}, source2[235:232]};
  wire [63:0]   extendResult_hi_hi_hi_lo_1 = {extendResult_hi_hi_hi_lo_hi, extendResult_hi_hi_hi_lo_lo};
  wire [31:0]   extendResult_hi_hi_hi_hi_lo = {{12{source2[247] & sign}}, source2[247:244], {12{source2[243] & sign}}, source2[243:240]};
  wire [31:0]   extendResult_hi_hi_hi_hi_hi = {{12{source2[255] & sign}}, source2[255:252], {12{source2[251] & sign}}, source2[251:248]};
  wire [63:0]   extendResult_hi_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi_hi, extendResult_hi_hi_hi_hi_lo};
  wire [127:0]  extendResult_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi_1, extendResult_hi_hi_hi_lo_1};
  wire [255:0]  extendResult_hi_hi_1 = {extendResult_hi_hi_hi_1, extendResult_hi_hi_lo_1};
  wire [511:0]  extendResult_hi_1 = {extendResult_hi_hi_1, extendResult_hi_lo_1};
  wire [63:0]   extendResult_lo_lo_lo_2 = {{16{source2[31] & sign}}, source2[31:16], {16{source2[15] & sign}}, source2[15:0]};
  wire [63:0]   extendResult_lo_lo_hi_2 = {{16{source2[63] & sign}}, source2[63:48], {16{source2[47] & sign}}, source2[47:32]};
  wire [127:0]  extendResult_lo_lo_2 = {extendResult_lo_lo_hi_2, extendResult_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_lo_2 = {{16{source2[95] & sign}}, source2[95:80], {16{source2[79] & sign}}, source2[79:64]};
  wire [63:0]   extendResult_lo_hi_hi_2 = {{16{source2[127] & sign}}, source2[127:112], {16{source2[111] & sign}}, source2[111:96]};
  wire [127:0]  extendResult_lo_hi_2 = {extendResult_lo_hi_hi_2, extendResult_lo_hi_lo_2};
  wire [255:0]  extendResult_lo_2 = {extendResult_lo_hi_2, extendResult_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_lo_2 = {{16{source2[159] & sign}}, source2[159:144], {16{source2[143] & sign}}, source2[143:128]};
  wire [63:0]   extendResult_hi_lo_hi_2 = {{16{source2[191] & sign}}, source2[191:176], {16{source2[175] & sign}}, source2[175:160]};
  wire [127:0]  extendResult_hi_lo_2 = {extendResult_hi_lo_hi_2, extendResult_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_lo_2 = {{16{source2[223] & sign}}, source2[223:208], {16{source2[207] & sign}}, source2[207:192]};
  wire [63:0]   extendResult_hi_hi_hi_2 = {{16{source2[255] & sign}}, source2[255:240], {16{source2[239] & sign}}, source2[239:224]};
  wire [127:0]  extendResult_hi_hi_2 = {extendResult_hi_hi_hi_2, extendResult_hi_hi_lo_2};
  wire [255:0]  extendResult_hi_2 = {extendResult_hi_hi_2, extendResult_hi_lo_2};
  wire [63:0]   extendResult_lo_lo_lo_lo_2 = {{24{source2[15] & sign}}, source2[15:8], {24{source2[7] & sign}}, source2[7:0]};
  wire [63:0]   extendResult_lo_lo_lo_hi_2 = {{24{source2[31] & sign}}, source2[31:24], {24{source2[23] & sign}}, source2[23:16]};
  wire [127:0]  extendResult_lo_lo_lo_3 = {extendResult_lo_lo_lo_hi_2, extendResult_lo_lo_lo_lo_2};
  wire [63:0]   extendResult_lo_lo_hi_lo_2 = {{24{source2[47] & sign}}, source2[47:40], {24{source2[39] & sign}}, source2[39:32]};
  wire [63:0]   extendResult_lo_lo_hi_hi_2 = {{24{source2[63] & sign}}, source2[63:56], {24{source2[55] & sign}}, source2[55:48]};
  wire [127:0]  extendResult_lo_lo_hi_3 = {extendResult_lo_lo_hi_hi_2, extendResult_lo_lo_hi_lo_2};
  wire [255:0]  extendResult_lo_lo_3 = {extendResult_lo_lo_hi_3, extendResult_lo_lo_lo_3};
  wire [63:0]   extendResult_lo_hi_lo_lo_2 = {{24{source2[79] & sign}}, source2[79:72], {24{source2[71] & sign}}, source2[71:64]};
  wire [63:0]   extendResult_lo_hi_lo_hi_2 = {{24{source2[95] & sign}}, source2[95:88], {24{source2[87] & sign}}, source2[87:80]};
  wire [127:0]  extendResult_lo_hi_lo_3 = {extendResult_lo_hi_lo_hi_2, extendResult_lo_hi_lo_lo_2};
  wire [63:0]   extendResult_lo_hi_hi_lo_2 = {{24{source2[111] & sign}}, source2[111:104], {24{source2[103] & sign}}, source2[103:96]};
  wire [63:0]   extendResult_lo_hi_hi_hi_2 = {{24{source2[127] & sign}}, source2[127:120], {24{source2[119] & sign}}, source2[119:112]};
  wire [127:0]  extendResult_lo_hi_hi_3 = {extendResult_lo_hi_hi_hi_2, extendResult_lo_hi_hi_lo_2};
  wire [255:0]  extendResult_lo_hi_3 = {extendResult_lo_hi_hi_3, extendResult_lo_hi_lo_3};
  wire [511:0]  extendResult_lo_3 = {extendResult_lo_hi_3, extendResult_lo_lo_3};
  wire [63:0]   extendResult_hi_lo_lo_lo_2 = {{24{source2[143] & sign}}, source2[143:136], {24{source2[135] & sign}}, source2[135:128]};
  wire [63:0]   extendResult_hi_lo_lo_hi_2 = {{24{source2[159] & sign}}, source2[159:152], {24{source2[151] & sign}}, source2[151:144]};
  wire [127:0]  extendResult_hi_lo_lo_3 = {extendResult_hi_lo_lo_hi_2, extendResult_hi_lo_lo_lo_2};
  wire [63:0]   extendResult_hi_lo_hi_lo_2 = {{24{source2[175] & sign}}, source2[175:168], {24{source2[167] & sign}}, source2[167:160]};
  wire [63:0]   extendResult_hi_lo_hi_hi_2 = {{24{source2[191] & sign}}, source2[191:184], {24{source2[183] & sign}}, source2[183:176]};
  wire [127:0]  extendResult_hi_lo_hi_3 = {extendResult_hi_lo_hi_hi_2, extendResult_hi_lo_hi_lo_2};
  wire [255:0]  extendResult_hi_lo_3 = {extendResult_hi_lo_hi_3, extendResult_hi_lo_lo_3};
  wire [63:0]   extendResult_hi_hi_lo_lo_2 = {{24{source2[207] & sign}}, source2[207:200], {24{source2[199] & sign}}, source2[199:192]};
  wire [63:0]   extendResult_hi_hi_lo_hi_2 = {{24{source2[223] & sign}}, source2[223:216], {24{source2[215] & sign}}, source2[215:208]};
  wire [127:0]  extendResult_hi_hi_lo_3 = {extendResult_hi_hi_lo_hi_2, extendResult_hi_hi_lo_lo_2};
  wire [63:0]   extendResult_hi_hi_hi_lo_2 = {{24{source2[239] & sign}}, source2[239:232], {24{source2[231] & sign}}, source2[231:224]};
  wire [63:0]   extendResult_hi_hi_hi_hi_2 = {{24{source2[255] & sign}}, source2[255:248], {24{source2[247] & sign}}, source2[247:240]};
  wire [127:0]  extendResult_hi_hi_hi_3 = {extendResult_hi_hi_hi_hi_2, extendResult_hi_hi_hi_lo_2};
  wire [255:0]  extendResult_hi_hi_3 = {extendResult_hi_hi_hi_3, extendResult_hi_hi_lo_3};
  wire [511:0]  extendResult_hi_3 = {extendResult_hi_hi_3, extendResult_hi_lo_3};
  wire [1023:0] extendResult =
    (eew1H[1] ? {512'h0, _extendResult_T_489[0] ? {extendResult_hi, extendResult_lo} : 512'h0} | (_extendResult_T_489[1] ? {extendResult_hi_1, extendResult_lo_1} : 1024'h0) : 1024'h0)
    | (eew1H[2] ? {512'h0, _extendResult_T_489[0] ? {extendResult_hi_2, extendResult_lo_2} : 512'h0} | (_extendResult_T_489[1] ? {extendResult_hi_3, extendResult_lo_3} : 1024'h0) : 1024'h0);
  assign out = isMaskDestination ? maskDestinationResult : extendResult[511:0];
endmodule

