
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_orderReduce,
                instReq_bits_decodeResult_floatMul,
  input  [1:0]  instReq_bits_decodeResult_fpExecutionType,
  input         instReq_bits_decodeResult_float,
                instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [10:0] instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_0_bits_fpReduceValid,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_1_bits_fpReduceValid,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_2_bits_fpReduceValid,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeReq_3_bits_fpReduceValid,
                exeReq_4_valid,
  input  [31:0] exeReq_4_bits_source1,
                exeReq_4_bits_source2,
  input  [2:0]  exeReq_4_bits_index,
  input         exeReq_4_bits_ffo,
                exeReq_4_bits_fpReduceValid,
                exeReq_5_valid,
  input  [31:0] exeReq_5_bits_source1,
                exeReq_5_bits_source2,
  input  [2:0]  exeReq_5_bits_index,
  input         exeReq_5_bits_ffo,
                exeReq_5_bits_fpReduceValid,
                exeReq_6_valid,
  input  [31:0] exeReq_6_bits_source1,
                exeReq_6_bits_source2,
  input  [2:0]  exeReq_6_bits_index,
  input         exeReq_6_bits_ffo,
                exeReq_6_bits_fpReduceValid,
                exeReq_7_valid,
  input  [31:0] exeReq_7_bits_source1,
                exeReq_7_bits_source2,
  input  [2:0]  exeReq_7_bits_index,
  input         exeReq_7_bits_ffo,
                exeReq_7_bits_fpReduceValid,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output [1:0]  exeResp_0_bits_offset,
  output [3:0]  exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output [1:0]  exeResp_1_bits_offset,
  output [3:0]  exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output [1:0]  exeResp_2_bits_offset,
  output [3:0]  exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output [1:0]  exeResp_3_bits_offset,
  output [3:0]  exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         exeResp_4_ready,
  output        exeResp_4_valid,
  output [4:0]  exeResp_4_bits_vd,
  output [1:0]  exeResp_4_bits_offset,
  output [3:0]  exeResp_4_bits_mask,
  output [31:0] exeResp_4_bits_data,
  output [2:0]  exeResp_4_bits_instructionIndex,
  input         exeResp_5_ready,
  output        exeResp_5_valid,
  output [4:0]  exeResp_5_bits_vd,
  output [1:0]  exeResp_5_bits_offset,
  output [3:0]  exeResp_5_bits_mask,
  output [31:0] exeResp_5_bits_data,
  output [2:0]  exeResp_5_bits_instructionIndex,
  input         exeResp_6_ready,
  output        exeResp_6_valid,
  output [4:0]  exeResp_6_bits_vd,
  output [1:0]  exeResp_6_bits_offset,
  output [3:0]  exeResp_6_bits_mask,
  output [31:0] exeResp_6_bits_data,
  output [2:0]  exeResp_6_bits_instructionIndex,
  input         exeResp_7_ready,
  output        exeResp_7_valid,
  output [4:0]  exeResp_7_bits_vd,
  output [1:0]  exeResp_7_bits_offset,
  output [3:0]  exeResp_7_bits_mask,
  output [31:0] exeResp_7_bits_data,
  output [2:0]  exeResp_7_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
                writeRelease_4,
                writeRelease_5,
                writeRelease_6,
                writeRelease_7,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
                tokenIO_4_maskRequestRelease,
                tokenIO_5_maskRequestRelease,
                tokenIO_6_maskRequestRelease,
                tokenIO_7_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output [1:0]  readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output [1:0]  readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output [1:0]  readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output [1:0]  readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readChannel_4_ready,
  output        readChannel_4_valid,
  output [4:0]  readChannel_4_bits_vs,
  output [1:0]  readChannel_4_bits_offset,
  output [2:0]  readChannel_4_bits_instructionIndex,
  input         readChannel_5_ready,
  output        readChannel_5_valid,
  output [4:0]  readChannel_5_bits_vs,
  output [1:0]  readChannel_5_bits_offset,
  output [2:0]  readChannel_5_bits_instructionIndex,
  input         readChannel_6_ready,
  output        readChannel_6_valid,
  output [4:0]  readChannel_6_bits_vs,
  output [1:0]  readChannel_6_bits_offset,
  output [2:0]  readChannel_6_bits_instructionIndex,
  input         readChannel_7_ready,
  output        readChannel_7_valid,
  output [4:0]  readChannel_7_bits_vs,
  output [1:0]  readChannel_7_bits_offset,
  output [2:0]  readChannel_7_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  input         readResult_4_valid,
  input  [31:0] readResult_4_bits,
  input         readResult_5_valid,
  input  [31:0] readResult_5_bits,
  input         readResult_6_valid,
  input  [31:0] readResult_6_bits,
  input         readResult_7_valid,
  input  [31:0] readResult_7_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
                laneMaskInput_4,
                laneMaskInput_5,
                laneMaskInput_6,
                laneMaskInput_7,
  input  [4:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
                laneMaskSelect_4,
                laneMaskSelect_5,
                laneMaskSelect_6,
                laneMaskSelect_7,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
                laneMaskSewSelect_4,
                laneMaskSewSelect_5,
                laneMaskSewSelect_6,
                laneMaskSewSelect_7,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input  [1:0]  v0UpdateVec_0_bits_offset,
  input  [3:0]  v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input  [1:0]  v0UpdateVec_1_bits_offset,
  input  [3:0]  v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input  [1:0]  v0UpdateVec_2_bits_offset,
  input  [3:0]  v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input  [1:0]  v0UpdateVec_3_bits_offset,
  input  [3:0]  v0UpdateVec_3_bits_mask,
  input         v0UpdateVec_4_valid,
  input  [31:0] v0UpdateVec_4_bits_data,
  input  [1:0]  v0UpdateVec_4_bits_offset,
  input  [3:0]  v0UpdateVec_4_bits_mask,
  input         v0UpdateVec_5_valid,
  input  [31:0] v0UpdateVec_5_bits_data,
  input  [1:0]  v0UpdateVec_5_bits_offset,
  input  [3:0]  v0UpdateVec_5_bits_mask,
  input         v0UpdateVec_6_valid,
  input  [31:0] v0UpdateVec_6_bits_data,
  input  [1:0]  v0UpdateVec_6_bits_offset,
  input  [3:0]  v0UpdateVec_6_bits_mask,
  input         v0UpdateVec_7_valid,
  input  [31:0] v0UpdateVec_7_bits_data,
  input  [1:0]  v0UpdateVec_7_bits_offset,
  input  [3:0]  v0UpdateVec_7_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire              readCrossBar_input_7_valid;
  wire              readCrossBar_input_6_valid;
  wire              readCrossBar_input_5_valid;
  wire              readCrossBar_input_4_valid;
  wire              readCrossBar_input_3_valid;
  wire              readCrossBar_input_2_valid;
  wire              readCrossBar_input_1_valid;
  wire              readCrossBar_input_0_valid;
  wire              _writeQueue_fifo_7_empty;
  wire              _writeQueue_fifo_7_full;
  wire              _writeQueue_fifo_7_error;
  wire [50:0]       _writeQueue_fifo_7_data_out;
  wire              _writeQueue_fifo_6_empty;
  wire              _writeQueue_fifo_6_full;
  wire              _writeQueue_fifo_6_error;
  wire [50:0]       _writeQueue_fifo_6_data_out;
  wire              _writeQueue_fifo_5_empty;
  wire              _writeQueue_fifo_5_full;
  wire              _writeQueue_fifo_5_error;
  wire [50:0]       _writeQueue_fifo_5_data_out;
  wire              _writeQueue_fifo_4_empty;
  wire              _writeQueue_fifo_4_full;
  wire              _writeQueue_fifo_4_error;
  wire [50:0]       _writeQueue_fifo_4_data_out;
  wire              _writeQueue_fifo_3_empty;
  wire              _writeQueue_fifo_3_full;
  wire              _writeQueue_fifo_3_error;
  wire [50:0]       _writeQueue_fifo_3_data_out;
  wire              _writeQueue_fifo_2_empty;
  wire              _writeQueue_fifo_2_full;
  wire              _writeQueue_fifo_2_error;
  wire [50:0]       _writeQueue_fifo_2_data_out;
  wire              _writeQueue_fifo_1_empty;
  wire              _writeQueue_fifo_1_full;
  wire              _writeQueue_fifo_1_error;
  wire [50:0]       _writeQueue_fifo_1_data_out;
  wire              _writeQueue_fifo_empty;
  wire              _writeQueue_fifo_full;
  wire              _writeQueue_fifo_error;
  wire [50:0]       _writeQueue_fifo_data_out;
  wire [255:0]      _extendUnit_out;
  wire              _reduceUnit_in_ready;
  wire              _reduceUnit_out_valid;
  wire [31:0]       _reduceUnit_out_bits_data;
  wire [3:0]        _reduceUnit_out_bits_mask;
  wire              _compressUnit_out_compressValid;
  wire [31:0]       _compressUnit_writeData;
  wire              _compressUnit_stageValid;
  wire              _readData_readDataQueue_fifo_7_empty;
  wire              _readData_readDataQueue_fifo_7_full;
  wire              _readData_readDataQueue_fifo_7_error;
  wire [31:0]       _readData_readDataQueue_fifo_7_data_out;
  wire              _readData_readDataQueue_fifo_6_empty;
  wire              _readData_readDataQueue_fifo_6_full;
  wire              _readData_readDataQueue_fifo_6_error;
  wire [31:0]       _readData_readDataQueue_fifo_6_data_out;
  wire              _readData_readDataQueue_fifo_5_empty;
  wire              _readData_readDataQueue_fifo_5_full;
  wire              _readData_readDataQueue_fifo_5_error;
  wire [31:0]       _readData_readDataQueue_fifo_5_data_out;
  wire              _readData_readDataQueue_fifo_4_empty;
  wire              _readData_readDataQueue_fifo_4_full;
  wire              _readData_readDataQueue_fifo_4_error;
  wire [31:0]       _readData_readDataQueue_fifo_4_data_out;
  wire              _readData_readDataQueue_fifo_3_empty;
  wire              _readData_readDataQueue_fifo_3_full;
  wire              _readData_readDataQueue_fifo_3_error;
  wire [31:0]       _readData_readDataQueue_fifo_3_data_out;
  wire              _readData_readDataQueue_fifo_2_empty;
  wire              _readData_readDataQueue_fifo_2_full;
  wire              _readData_readDataQueue_fifo_2_error;
  wire [31:0]       _readData_readDataQueue_fifo_2_data_out;
  wire              _readData_readDataQueue_fifo_1_empty;
  wire              _readData_readDataQueue_fifo_1_full;
  wire              _readData_readDataQueue_fifo_1_error;
  wire [31:0]       _readData_readDataQueue_fifo_1_data_out;
  wire              _readData_readDataQueue_fifo_empty;
  wire              _readData_readDataQueue_fifo_full;
  wire              _readData_readDataQueue_fifo_error;
  wire [31:0]       _readData_readDataQueue_fifo_data_out;
  wire              _readMessageQueue_fifo_7_empty;
  wire              _readMessageQueue_fifo_7_full;
  wire              _readMessageQueue_fifo_7_error;
  wire [9:0]        _readMessageQueue_fifo_7_data_out;
  wire              _readMessageQueue_fifo_6_empty;
  wire              _readMessageQueue_fifo_6_full;
  wire              _readMessageQueue_fifo_6_error;
  wire [9:0]        _readMessageQueue_fifo_6_data_out;
  wire              _readMessageQueue_fifo_5_empty;
  wire              _readMessageQueue_fifo_5_full;
  wire              _readMessageQueue_fifo_5_error;
  wire [9:0]        _readMessageQueue_fifo_5_data_out;
  wire              _readMessageQueue_fifo_4_empty;
  wire              _readMessageQueue_fifo_4_full;
  wire              _readMessageQueue_fifo_4_error;
  wire [9:0]        _readMessageQueue_fifo_4_data_out;
  wire              _readMessageQueue_fifo_3_empty;
  wire              _readMessageQueue_fifo_3_full;
  wire              _readMessageQueue_fifo_3_error;
  wire [9:0]        _readMessageQueue_fifo_3_data_out;
  wire              _readMessageQueue_fifo_2_empty;
  wire              _readMessageQueue_fifo_2_full;
  wire              _readMessageQueue_fifo_2_error;
  wire [9:0]        _readMessageQueue_fifo_2_data_out;
  wire              _readMessageQueue_fifo_1_empty;
  wire              _readMessageQueue_fifo_1_full;
  wire              _readMessageQueue_fifo_1_error;
  wire [9:0]        _readMessageQueue_fifo_1_data_out;
  wire              _readMessageQueue_fifo_empty;
  wire              _readMessageQueue_fifo_full;
  wire              _readMessageQueue_fifo_error;
  wire [9:0]        _readMessageQueue_fifo_data_out;
  wire              _reorderQueueVec_fifo_7_empty;
  wire              _reorderQueueVec_fifo_7_full;
  wire              _reorderQueueVec_fifo_7_error;
  wire [39:0]       _reorderQueueVec_fifo_7_data_out;
  wire              _reorderQueueVec_fifo_6_empty;
  wire              _reorderQueueVec_fifo_6_full;
  wire              _reorderQueueVec_fifo_6_error;
  wire [39:0]       _reorderQueueVec_fifo_6_data_out;
  wire              _reorderQueueVec_fifo_5_empty;
  wire              _reorderQueueVec_fifo_5_full;
  wire              _reorderQueueVec_fifo_5_error;
  wire [39:0]       _reorderQueueVec_fifo_5_data_out;
  wire              _reorderQueueVec_fifo_4_empty;
  wire              _reorderQueueVec_fifo_4_full;
  wire              _reorderQueueVec_fifo_4_error;
  wire [39:0]       _reorderQueueVec_fifo_4_data_out;
  wire              _reorderQueueVec_fifo_3_empty;
  wire              _reorderQueueVec_fifo_3_full;
  wire              _reorderQueueVec_fifo_3_error;
  wire [39:0]       _reorderQueueVec_fifo_3_data_out;
  wire              _reorderQueueVec_fifo_2_empty;
  wire              _reorderQueueVec_fifo_2_full;
  wire              _reorderQueueVec_fifo_2_error;
  wire [39:0]       _reorderQueueVec_fifo_2_data_out;
  wire              _reorderQueueVec_fifo_1_empty;
  wire              _reorderQueueVec_fifo_1_full;
  wire              _reorderQueueVec_fifo_1_error;
  wire [39:0]       _reorderQueueVec_fifo_1_data_out;
  wire              _reorderQueueVec_fifo_empty;
  wire              _reorderQueueVec_fifo_full;
  wire              _reorderQueueVec_fifo_error;
  wire [39:0]       _reorderQueueVec_fifo_data_out;
  wire              _compressUnitResultQueue_fifo_empty;
  wire              _compressUnitResultQueue_fifo_full;
  wire              _compressUnitResultQueue_fifo_error;
  wire [302:0]      _compressUnitResultQueue_fifo_data_out;
  wire              _readWaitQueue_fifo_empty;
  wire              _readWaitQueue_fifo_full;
  wire              _readWaitQueue_fifo_error;
  wire [32:0]       _readWaitQueue_fifo_data_out;
  wire              _readCrossBar_input_0_ready;
  wire              _readCrossBar_input_1_ready;
  wire              _readCrossBar_input_2_ready;
  wire              _readCrossBar_input_3_ready;
  wire              _readCrossBar_input_4_ready;
  wire              _readCrossBar_input_5_ready;
  wire              _readCrossBar_input_6_ready;
  wire              _readCrossBar_input_7_ready;
  wire              _readCrossBar_output_0_valid;
  wire [4:0]        _readCrossBar_output_0_bits_vs;
  wire [1:0]        _readCrossBar_output_0_bits_offset;
  wire [2:0]        _readCrossBar_output_0_bits_writeIndex;
  wire              _readCrossBar_output_1_valid;
  wire [4:0]        _readCrossBar_output_1_bits_vs;
  wire [1:0]        _readCrossBar_output_1_bits_offset;
  wire [2:0]        _readCrossBar_output_1_bits_writeIndex;
  wire              _readCrossBar_output_2_valid;
  wire [4:0]        _readCrossBar_output_2_bits_vs;
  wire [1:0]        _readCrossBar_output_2_bits_offset;
  wire [2:0]        _readCrossBar_output_2_bits_writeIndex;
  wire              _readCrossBar_output_3_valid;
  wire [4:0]        _readCrossBar_output_3_bits_vs;
  wire [1:0]        _readCrossBar_output_3_bits_offset;
  wire [2:0]        _readCrossBar_output_3_bits_writeIndex;
  wire              _readCrossBar_output_4_valid;
  wire [4:0]        _readCrossBar_output_4_bits_vs;
  wire [1:0]        _readCrossBar_output_4_bits_offset;
  wire [2:0]        _readCrossBar_output_4_bits_writeIndex;
  wire              _readCrossBar_output_5_valid;
  wire [4:0]        _readCrossBar_output_5_bits_vs;
  wire [1:0]        _readCrossBar_output_5_bits_offset;
  wire [2:0]        _readCrossBar_output_5_bits_writeIndex;
  wire              _readCrossBar_output_6_valid;
  wire [4:0]        _readCrossBar_output_6_bits_vs;
  wire [1:0]        _readCrossBar_output_6_bits_offset;
  wire [2:0]        _readCrossBar_output_6_bits_writeIndex;
  wire              _readCrossBar_output_7_valid;
  wire [4:0]        _readCrossBar_output_7_bits_vs;
  wire [1:0]        _readCrossBar_output_7_bits_offset;
  wire [2:0]        _readCrossBar_output_7_bits_writeIndex;
  wire              _accessCountQueue_fifo_empty;
  wire              _accessCountQueue_fifo_full;
  wire              _accessCountQueue_fifo_error;
  wire [31:0]       _accessCountQueue_fifo_data_out;
  wire              _slideAddressGen_indexDeq_valid;
  wire [7:0]        _slideAddressGen_indexDeq_bits_needRead;
  wire [7:0]        _slideAddressGen_indexDeq_bits_elementValid;
  wire [7:0]        _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [15:0]       _slideAddressGen_indexDeq_bits_readOffset;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_4;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_5;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_6;
  wire [2:0]        _slideAddressGen_indexDeq_bits_accessLane_7;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_4;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_5;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_6;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_7;
  wire [7:0]        _slideAddressGen_indexDeq_bits_executeGroup;
  wire [15:0]       _slideAddressGen_indexDeq_bits_readDataOffset;
  wire              _slideAddressGen_indexDeq_bits_last;
  wire [7:0]        _slideAddressGen_slideGroupOut;
  wire              _exeRequestQueue_queue_fifo_7_empty;
  wire              _exeRequestQueue_queue_fifo_7_full;
  wire              _exeRequestQueue_queue_fifo_7_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_7_data_out;
  wire              _exeRequestQueue_queue_fifo_6_empty;
  wire              _exeRequestQueue_queue_fifo_6_full;
  wire              _exeRequestQueue_queue_fifo_6_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_6_data_out;
  wire              _exeRequestQueue_queue_fifo_5_empty;
  wire              _exeRequestQueue_queue_fifo_5_full;
  wire              _exeRequestQueue_queue_fifo_5_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_5_data_out;
  wire              _exeRequestQueue_queue_fifo_4_empty;
  wire              _exeRequestQueue_queue_fifo_4_full;
  wire              _exeRequestQueue_queue_fifo_4_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_4_data_out;
  wire              _exeRequestQueue_queue_fifo_3_empty;
  wire              _exeRequestQueue_queue_fifo_3_full;
  wire              _exeRequestQueue_queue_fifo_3_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_3_data_out;
  wire              _exeRequestQueue_queue_fifo_2_empty;
  wire              _exeRequestQueue_queue_fifo_2_full;
  wire              _exeRequestQueue_queue_fifo_2_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_2_data_out;
  wire              _exeRequestQueue_queue_fifo_1_empty;
  wire              _exeRequestQueue_queue_fifo_1_full;
  wire              _exeRequestQueue_queue_fifo_1_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_1_data_out;
  wire              _exeRequestQueue_queue_fifo_empty;
  wire              _exeRequestQueue_queue_fifo_full;
  wire              _exeRequestQueue_queue_fifo_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_data_out;
  wire              _maskedWrite_in_0_ready;
  wire              _maskedWrite_in_1_ready;
  wire              _maskedWrite_in_2_ready;
  wire              _maskedWrite_in_3_ready;
  wire              _maskedWrite_in_4_ready;
  wire              _maskedWrite_in_5_ready;
  wire              _maskedWrite_in_6_ready;
  wire              _maskedWrite_in_7_ready;
  wire              _maskedWrite_out_0_valid;
  wire              _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_0_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_0_bits_writeData_groupCounter;
  wire              _maskedWrite_out_1_valid;
  wire              _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_1_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_1_bits_writeData_groupCounter;
  wire              _maskedWrite_out_2_valid;
  wire              _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_2_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_2_bits_writeData_groupCounter;
  wire              _maskedWrite_out_3_valid;
  wire              _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_3_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_3_bits_writeData_groupCounter;
  wire              _maskedWrite_out_4_valid;
  wire              _maskedWrite_out_4_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_4_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_4_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_4_bits_writeData_groupCounter;
  wire              _maskedWrite_out_5_valid;
  wire              _maskedWrite_out_5_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_5_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_5_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_5_bits_writeData_groupCounter;
  wire              _maskedWrite_out_6_valid;
  wire              _maskedWrite_out_6_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_6_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_6_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_6_bits_writeData_groupCounter;
  wire              _maskedWrite_out_7_valid;
  wire              _maskedWrite_out_7_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_7_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_7_bits_writeData_mask;
  wire [5:0]        _maskedWrite_out_7_bits_writeData_groupCounter;
  wire              _maskedWrite_readChannel_0_valid;
  wire [4:0]        _maskedWrite_readChannel_0_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_0_bits_offset;
  wire              _maskedWrite_readChannel_1_valid;
  wire [4:0]        _maskedWrite_readChannel_1_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_1_bits_offset;
  wire              _maskedWrite_readChannel_2_valid;
  wire [4:0]        _maskedWrite_readChannel_2_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_2_bits_offset;
  wire              _maskedWrite_readChannel_3_valid;
  wire [4:0]        _maskedWrite_readChannel_3_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_3_bits_offset;
  wire              _maskedWrite_readChannel_4_valid;
  wire [4:0]        _maskedWrite_readChannel_4_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_4_bits_offset;
  wire              _maskedWrite_readChannel_5_valid;
  wire [4:0]        _maskedWrite_readChannel_5_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_5_bits_offset;
  wire              _maskedWrite_readChannel_6_valid;
  wire [4:0]        _maskedWrite_readChannel_6_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_6_bits_offset;
  wire              _maskedWrite_readChannel_7_valid;
  wire [4:0]        _maskedWrite_readChannel_7_bits_vs;
  wire [1:0]        _maskedWrite_readChannel_7_bits_offset;
  wire              _maskedWrite_stageClear;
  wire              writeQueue_7_almostFull;
  wire              writeQueue_7_almostEmpty;
  wire              writeQueue_6_almostFull;
  wire              writeQueue_6_almostEmpty;
  wire              writeQueue_5_almostFull;
  wire              writeQueue_5_almostEmpty;
  wire              writeQueue_4_almostFull;
  wire              writeQueue_4_almostEmpty;
  wire              writeQueue_3_almostFull;
  wire              writeQueue_3_almostEmpty;
  wire              writeQueue_2_almostFull;
  wire              writeQueue_2_almostEmpty;
  wire              writeQueue_1_almostFull;
  wire              writeQueue_1_almostEmpty;
  wire              writeQueue_0_almostFull;
  wire              writeQueue_0_almostEmpty;
  wire              readData_readDataQueue_7_almostFull;
  wire              readData_readDataQueue_7_almostEmpty;
  wire              readData_readDataQueue_6_almostFull;
  wire              readData_readDataQueue_6_almostEmpty;
  wire              readData_readDataQueue_5_almostFull;
  wire              readData_readDataQueue_5_almostEmpty;
  wire              readData_readDataQueue_4_almostFull;
  wire              readData_readDataQueue_4_almostEmpty;
  wire              readData_readDataQueue_3_almostFull;
  wire              readData_readDataQueue_3_almostEmpty;
  wire              readData_readDataQueue_2_almostFull;
  wire              readData_readDataQueue_2_almostEmpty;
  wire              readData_readDataQueue_1_almostFull;
  wire              readData_readDataQueue_1_almostEmpty;
  wire              readData_readDataQueue_almostFull;
  wire              readData_readDataQueue_almostEmpty;
  wire              readMessageQueue_7_almostFull;
  wire              readMessageQueue_7_almostEmpty;
  wire              readMessageQueue_6_almostFull;
  wire              readMessageQueue_6_almostEmpty;
  wire              readMessageQueue_5_almostFull;
  wire              readMessageQueue_5_almostEmpty;
  wire              readMessageQueue_4_almostFull;
  wire              readMessageQueue_4_almostEmpty;
  wire              readMessageQueue_3_almostFull;
  wire              readMessageQueue_3_almostEmpty;
  wire              readMessageQueue_2_almostFull;
  wire              readMessageQueue_2_almostEmpty;
  wire              readMessageQueue_1_almostFull;
  wire              readMessageQueue_1_almostEmpty;
  wire              readMessageQueue_almostFull;
  wire              readMessageQueue_almostEmpty;
  wire              reorderQueueVec_7_almostFull;
  wire              reorderQueueVec_7_almostEmpty;
  wire              reorderQueueVec_6_almostFull;
  wire              reorderQueueVec_6_almostEmpty;
  wire              reorderQueueVec_5_almostFull;
  wire              reorderQueueVec_5_almostEmpty;
  wire              reorderQueueVec_4_almostFull;
  wire              reorderQueueVec_4_almostEmpty;
  wire              reorderQueueVec_3_almostFull;
  wire              reorderQueueVec_3_almostEmpty;
  wire              reorderQueueVec_2_almostFull;
  wire              reorderQueueVec_2_almostEmpty;
  wire              reorderQueueVec_1_almostFull;
  wire              reorderQueueVec_1_almostEmpty;
  wire              reorderQueueVec_0_almostFull;
  wire              reorderQueueVec_0_almostEmpty;
  wire              compressUnitResultQueue_almostFull;
  wire              compressUnitResultQueue_almostEmpty;
  wire              readWaitQueue_almostFull;
  wire              readWaitQueue_almostEmpty;
  wire              accessCountQueue_almostFull;
  wire              accessCountQueue_almostEmpty;
  wire              exeRequestQueue_7_almostFull;
  wire              exeRequestQueue_7_almostEmpty;
  wire              exeRequestQueue_6_almostFull;
  wire              exeRequestQueue_6_almostEmpty;
  wire              exeRequestQueue_5_almostFull;
  wire              exeRequestQueue_5_almostEmpty;
  wire              exeRequestQueue_4_almostFull;
  wire              exeRequestQueue_4_almostEmpty;
  wire              exeRequestQueue_3_almostFull;
  wire              exeRequestQueue_3_almostEmpty;
  wire              exeRequestQueue_2_almostFull;
  wire              exeRequestQueue_2_almostEmpty;
  wire              exeRequestQueue_1_almostFull;
  wire              exeRequestQueue_1_almostEmpty;
  wire              exeRequestQueue_0_almostFull;
  wire              exeRequestQueue_0_almostEmpty;
  wire [31:0]       reorderQueueVec_7_deq_bits_data;
  wire [31:0]       reorderQueueVec_6_deq_bits_data;
  wire [31:0]       reorderQueueVec_5_deq_bits_data;
  wire [31:0]       reorderQueueVec_4_deq_bits_data;
  wire [31:0]       reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_deq_bits_data;
  wire [3:0]        accessCountEnq_7;
  wire [3:0]        accessCountEnq_6;
  wire [3:0]        accessCountEnq_5;
  wire [3:0]        accessCountEnq_4;
  wire [3:0]        accessCountEnq_3;
  wire [3:0]        accessCountEnq_2;
  wire [3:0]        accessCountEnq_1;
  wire [3:0]        accessCountEnq_0;
  wire              exeResp_0_ready_0 = exeResp_0_ready;
  wire              exeResp_1_ready_0 = exeResp_1_ready;
  wire              exeResp_2_ready_0 = exeResp_2_ready;
  wire              exeResp_3_ready_0 = exeResp_3_ready;
  wire              exeResp_4_ready_0 = exeResp_4_ready;
  wire              exeResp_5_ready_0 = exeResp_5_ready;
  wire              exeResp_6_ready_0 = exeResp_6_ready;
  wire              exeResp_7_ready_0 = exeResp_7_ready;
  wire              readChannel_0_ready_0 = readChannel_0_ready;
  wire              readChannel_1_ready_0 = readChannel_1_ready;
  wire              readChannel_2_ready_0 = readChannel_2_ready;
  wire              readChannel_3_ready_0 = readChannel_3_ready;
  wire              readChannel_4_ready_0 = readChannel_4_ready;
  wire              readChannel_5_ready_0 = readChannel_5_ready;
  wire              readChannel_6_ready_0 = readChannel_6_ready;
  wire              readChannel_7_ready_0 = readChannel_7_ready;
  wire              gatherData_ready_0 = gatherData_ready;
  wire              exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]       exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]       exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]        exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire              exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire              exeRequestQueue_0_enq_bits_fpReduceValid = exeReq_0_bits_fpReduceValid;
  wire              exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]       exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]       exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]        exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire              exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire              exeRequestQueue_1_enq_bits_fpReduceValid = exeReq_1_bits_fpReduceValid;
  wire              exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]       exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]       exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]        exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire              exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire              exeRequestQueue_2_enq_bits_fpReduceValid = exeReq_2_bits_fpReduceValid;
  wire              exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]       exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]       exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]        exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire              exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire              exeRequestQueue_3_enq_bits_fpReduceValid = exeReq_3_bits_fpReduceValid;
  wire              exeRequestQueue_4_enq_valid = exeReq_4_valid;
  wire [31:0]       exeRequestQueue_4_enq_bits_source1 = exeReq_4_bits_source1;
  wire [31:0]       exeRequestQueue_4_enq_bits_source2 = exeReq_4_bits_source2;
  wire [2:0]        exeRequestQueue_4_enq_bits_index = exeReq_4_bits_index;
  wire              exeRequestQueue_4_enq_bits_ffo = exeReq_4_bits_ffo;
  wire              exeRequestQueue_4_enq_bits_fpReduceValid = exeReq_4_bits_fpReduceValid;
  wire              exeRequestQueue_5_enq_valid = exeReq_5_valid;
  wire [31:0]       exeRequestQueue_5_enq_bits_source1 = exeReq_5_bits_source1;
  wire [31:0]       exeRequestQueue_5_enq_bits_source2 = exeReq_5_bits_source2;
  wire [2:0]        exeRequestQueue_5_enq_bits_index = exeReq_5_bits_index;
  wire              exeRequestQueue_5_enq_bits_ffo = exeReq_5_bits_ffo;
  wire              exeRequestQueue_5_enq_bits_fpReduceValid = exeReq_5_bits_fpReduceValid;
  wire              exeRequestQueue_6_enq_valid = exeReq_6_valid;
  wire [31:0]       exeRequestQueue_6_enq_bits_source1 = exeReq_6_bits_source1;
  wire [31:0]       exeRequestQueue_6_enq_bits_source2 = exeReq_6_bits_source2;
  wire [2:0]        exeRequestQueue_6_enq_bits_index = exeReq_6_bits_index;
  wire              exeRequestQueue_6_enq_bits_ffo = exeReq_6_bits_ffo;
  wire              exeRequestQueue_6_enq_bits_fpReduceValid = exeReq_6_bits_fpReduceValid;
  wire              exeRequestQueue_7_enq_valid = exeReq_7_valid;
  wire [31:0]       exeRequestQueue_7_enq_bits_source1 = exeReq_7_bits_source1;
  wire [31:0]       exeRequestQueue_7_enq_bits_source2 = exeReq_7_bits_source2;
  wire [2:0]        exeRequestQueue_7_enq_bits_index = exeReq_7_bits_index;
  wire              exeRequestQueue_7_enq_bits_ffo = exeReq_7_bits_ffo;
  wire              exeRequestQueue_7_enq_bits_fpReduceValid = exeReq_7_bits_fpReduceValid;
  wire              reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire              reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire              reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire              reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire              reorderQueueVec_4_enq_valid = readResult_4_valid;
  wire              reorderQueueVec_5_enq_valid = readResult_5_valid;
  wire              reorderQueueVec_6_enq_valid = readResult_6_valid;
  wire              reorderQueueVec_7_enq_valid = readResult_7_valid;
  wire              readMessageQueue_deq_ready = readResult_0_valid;
  wire              readMessageQueue_1_deq_ready = readResult_1_valid;
  wire              readMessageQueue_2_deq_ready = readResult_2_valid;
  wire              readMessageQueue_3_deq_ready = readResult_3_valid;
  wire              readMessageQueue_4_deq_ready = readResult_4_valid;
  wire              readMessageQueue_5_deq_ready = readResult_5_valid;
  wire              readMessageQueue_6_deq_ready = readResult_6_valid;
  wire              readMessageQueue_7_deq_ready = readResult_7_valid;
  wire [7:0]        checkVec_checkResult_lo_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_lo_hi_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_hi_14 = 8'hFF;
  wire [1:0]        checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_4_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_5_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_6_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_7_1_2 = 2'h0;
  wire [15:0]       checkVec_checkResult_lo_14 = 16'hFFFF;
  wire [15:0]       checkVec_checkResult_hi_14 = 16'hFFFF;
  wire [31:0]       checkVec_2_0 = 32'hFFFFFFFF;
  wire [3:0]        checkVec_checkResult_lo_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_lo_hi_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_hi_15 = 4'h0;
  wire [15:0]       checkVec_2_1 = 16'h0;
  wire [2:0]        readVS1Req_requestIndex = 3'h0;
  wire [2:0]        selectExecuteReq_0_bits_requestIndex = 3'h0;
  wire [2:0]        selectExecuteReq_1_bits_requestIndex = 3'h1;
  wire [2:0]        selectExecuteReq_2_bits_requestIndex = 3'h2;
  wire [2:0]        selectExecuteReq_3_bits_requestIndex = 3'h3;
  wire [2:0]        selectExecuteReq_4_bits_requestIndex = 3'h4;
  wire [2:0]        selectExecuteReq_5_bits_requestIndex = 3'h5;
  wire [2:0]        selectExecuteReq_6_bits_requestIndex = 3'h6;
  wire [2:0]        selectExecuteReq_7_bits_requestIndex = 3'h7;
  wire [7:0]        checkVec_checkResult_lo_15 = 8'h0;
  wire [7:0]        checkVec_checkResult_hi_15 = 8'h0;
  wire              vs1Split_0_2 = 1'h1;
  wire [1:0]        readChannel_0_bits_readSource = 2'h2;
  wire [1:0]        readChannel_1_bits_readSource = 2'h2;
  wire [1:0]        readChannel_2_bits_readSource = 2'h2;
  wire [1:0]        readChannel_3_bits_readSource = 2'h2;
  wire [1:0]        readChannel_4_bits_readSource = 2'h2;
  wire [1:0]        readChannel_5_bits_readSource = 2'h2;
  wire [1:0]        readChannel_6_bits_readSource = 2'h2;
  wire [1:0]        readChannel_7_bits_readSource = 2'h2;
  wire              exeResp_0_bits_last = 1'h0;
  wire              exeResp_1_bits_last = 1'h0;
  wire              exeResp_2_bits_last = 1'h0;
  wire              exeResp_3_bits_last = 1'h0;
  wire              exeResp_4_bits_last = 1'h0;
  wire              exeResp_5_bits_last = 1'h0;
  wire              exeResp_6_bits_last = 1'h0;
  wire              exeResp_7_bits_last = 1'h0;
  wire              writeRequest_0_ffoByOther = 1'h0;
  wire              writeRequest_1_ffoByOther = 1'h0;
  wire              writeRequest_2_ffoByOther = 1'h0;
  wire              writeRequest_3_ffoByOther = 1'h0;
  wire              writeRequest_4_ffoByOther = 1'h0;
  wire              writeRequest_5_ffoByOther = 1'h0;
  wire              writeRequest_6_ffoByOther = 1'h0;
  wire              writeRequest_7_ffoByOther = 1'h0;
  wire              writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire              writeQueue_0_deq_valid;
  wire [3:0]        writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_0_deq_bits_writeData_data;
  wire              writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire              writeQueue_1_deq_valid;
  wire [3:0]        writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_1_deq_bits_writeData_data;
  wire              writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire              writeQueue_2_deq_valid;
  wire [3:0]        writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_2_deq_bits_writeData_data;
  wire              writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire              writeQueue_3_deq_valid;
  wire [3:0]        writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_3_deq_bits_writeData_data;
  wire              writeQueue_4_deq_ready = exeResp_4_ready_0;
  wire              writeQueue_4_deq_valid;
  wire [3:0]        writeQueue_4_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_4_deq_bits_writeData_data;
  wire              writeQueue_5_deq_ready = exeResp_5_ready_0;
  wire              writeQueue_5_deq_valid;
  wire [3:0]        writeQueue_5_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_5_deq_bits_writeData_data;
  wire              writeQueue_6_deq_ready = exeResp_6_ready_0;
  wire              writeQueue_6_deq_valid;
  wire [3:0]        writeQueue_6_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_6_deq_bits_writeData_data;
  wire              writeQueue_7_deq_ready = exeResp_7_ready_0;
  wire              writeQueue_7_deq_valid;
  wire [3:0]        writeQueue_7_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_7_deq_bits_writeData_data;
  wire              gatherResponse;
  reg  [31:0]       v0_0;
  reg  [31:0]       v0_1;
  reg  [31:0]       v0_2;
  reg  [31:0]       v0_3;
  reg  [31:0]       v0_4;
  reg  [31:0]       v0_5;
  reg  [31:0]       v0_6;
  reg  [31:0]       v0_7;
  reg  [31:0]       v0_8;
  reg  [31:0]       v0_9;
  reg  [31:0]       v0_10;
  reg  [31:0]       v0_11;
  reg  [31:0]       v0_12;
  reg  [31:0]       v0_13;
  reg  [31:0]       v0_14;
  reg  [31:0]       v0_15;
  reg  [31:0]       v0_16;
  reg  [31:0]       v0_17;
  reg  [31:0]       v0_18;
  reg  [31:0]       v0_19;
  reg  [31:0]       v0_20;
  reg  [31:0]       v0_21;
  reg  [31:0]       v0_22;
  reg  [31:0]       v0_23;
  reg  [31:0]       v0_24;
  reg  [31:0]       v0_25;
  reg  [31:0]       v0_26;
  reg  [31:0]       v0_27;
  reg  [31:0]       v0_28;
  reg  [31:0]       v0_29;
  reg  [31:0]       v0_30;
  reg  [31:0]       v0_31;
  wire [15:0]       maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]       maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]       maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]       maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]       maskExt_lo_4 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_4 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]       maskExt_lo_5 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_5 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]       maskExt_lo_6 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_6 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]       maskExt_lo_7 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_7 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]       maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]       maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]       maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]       maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]       maskExt_lo_12 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_12 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]       maskExt_lo_13 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_13 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]       maskExt_lo_14 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_14 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]       maskExt_lo_15 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_15 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]       maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]       maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]       maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]       maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]       maskExt_lo_20 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_20 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]       maskExt_lo_21 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_21 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]       maskExt_lo_22 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_22 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]       maskExt_lo_23 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_23 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]       maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]       maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]       maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]       maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]       maskExt_lo_28 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_28 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]       maskExt_lo_29 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_29 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]       maskExt_lo_30 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_30 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]       maskExt_lo_31 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_31 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [63:0]       _GEN = {v0_1, v0_0};
  wire [63:0]       regroupV0_lo_lo_lo_lo;
  assign regroupV0_lo_lo_lo_lo = _GEN;
  wire [63:0]       regroupV0_lo_lo_lo_lo_9;
  assign regroupV0_lo_lo_lo_lo_9 = _GEN;
  wire [63:0]       regroupV0_lo_lo_lo_lo_18;
  assign regroupV0_lo_lo_lo_lo_18 = _GEN;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo = _GEN;
  wire [63:0]       selectReadStageMask_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]       maskForDestination_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_lo = _GEN;
  wire [63:0]       _GEN_0 = {v0_3, v0_2};
  wire [63:0]       regroupV0_lo_lo_lo_hi;
  assign regroupV0_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       regroupV0_lo_lo_lo_hi_9;
  assign regroupV0_lo_lo_lo_hi_9 = _GEN_0;
  wire [63:0]       regroupV0_lo_lo_lo_hi_18;
  assign regroupV0_lo_lo_lo_hi_18 = _GEN_0;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       selectReadStageMask_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]       maskForDestination_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_hi = _GEN_0;
  wire [127:0]      regroupV0_lo_lo_lo = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [63:0]       _GEN_1 = {v0_5, v0_4};
  wire [63:0]       regroupV0_lo_lo_hi_lo;
  assign regroupV0_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       regroupV0_lo_lo_hi_lo_9;
  assign regroupV0_lo_lo_hi_lo_9 = _GEN_1;
  wire [63:0]       regroupV0_lo_lo_hi_lo_18;
  assign regroupV0_lo_lo_hi_lo_18 = _GEN_1;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       selectReadStageMask_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]       maskForDestination_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       _GEN_2 = {v0_7, v0_6};
  wire [63:0]       regroupV0_lo_lo_hi_hi;
  assign regroupV0_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       regroupV0_lo_lo_hi_hi_9;
  assign regroupV0_lo_lo_hi_hi_9 = _GEN_2;
  wire [63:0]       regroupV0_lo_lo_hi_hi_18;
  assign regroupV0_lo_lo_hi_hi_18 = _GEN_2;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       selectReadStageMask_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]       maskForDestination_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_hi_hi = _GEN_2;
  wire [127:0]      regroupV0_lo_lo_hi = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [255:0]      regroupV0_lo_lo = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [63:0]       _GEN_3 = {v0_9, v0_8};
  wire [63:0]       regroupV0_lo_hi_lo_lo;
  assign regroupV0_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       regroupV0_lo_hi_lo_lo_9;
  assign regroupV0_lo_hi_lo_lo_9 = _GEN_3;
  wire [63:0]       regroupV0_lo_hi_lo_lo_18;
  assign regroupV0_lo_hi_lo_lo_18 = _GEN_3;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       selectReadStageMask_lo_hi_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]       maskForDestination_lo_hi_lo_lo;
  assign maskForDestination_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       _GEN_4 = {v0_11, v0_10};
  wire [63:0]       regroupV0_lo_hi_lo_hi;
  assign regroupV0_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       regroupV0_lo_hi_lo_hi_9;
  assign regroupV0_lo_hi_lo_hi_9 = _GEN_4;
  wire [63:0]       regroupV0_lo_hi_lo_hi_18;
  assign regroupV0_lo_hi_lo_hi_18 = _GEN_4;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       selectReadStageMask_lo_hi_lo_hi;
  assign selectReadStageMask_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]       maskForDestination_lo_hi_lo_hi;
  assign maskForDestination_lo_hi_lo_hi = _GEN_4;
  wire [127:0]      regroupV0_lo_hi_lo = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [63:0]       _GEN_5 = {v0_13, v0_12};
  wire [63:0]       regroupV0_lo_hi_hi_lo;
  assign regroupV0_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       regroupV0_lo_hi_hi_lo_9;
  assign regroupV0_lo_hi_hi_lo_9 = _GEN_5;
  wire [63:0]       regroupV0_lo_hi_hi_lo_18;
  assign regroupV0_lo_hi_hi_lo_18 = _GEN_5;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       selectReadStageMask_lo_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]       maskForDestination_lo_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       _GEN_6 = {v0_15, v0_14};
  wire [63:0]       regroupV0_lo_hi_hi_hi;
  assign regroupV0_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       regroupV0_lo_hi_hi_hi_9;
  assign regroupV0_lo_hi_hi_hi_9 = _GEN_6;
  wire [63:0]       regroupV0_lo_hi_hi_hi_18;
  assign regroupV0_lo_hi_hi_hi_18 = _GEN_6;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       selectReadStageMask_lo_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]       maskForDestination_lo_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_hi = _GEN_6;
  wire [127:0]      regroupV0_lo_hi_hi = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [255:0]      regroupV0_lo_hi = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [511:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]       _GEN_7 = {v0_17, v0_16};
  wire [63:0]       regroupV0_hi_lo_lo_lo;
  assign regroupV0_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       regroupV0_hi_lo_lo_lo_9;
  assign regroupV0_hi_lo_lo_lo_9 = _GEN_7;
  wire [63:0]       regroupV0_hi_lo_lo_lo_18;
  assign regroupV0_hi_lo_lo_lo_18 = _GEN_7;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       selectReadStageMask_hi_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]       maskForDestination_hi_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       _GEN_8 = {v0_19, v0_18};
  wire [63:0]       regroupV0_hi_lo_lo_hi;
  assign regroupV0_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       regroupV0_hi_lo_lo_hi_9;
  assign regroupV0_hi_lo_lo_hi_9 = _GEN_8;
  wire [63:0]       regroupV0_hi_lo_lo_hi_18;
  assign regroupV0_hi_lo_lo_hi_18 = _GEN_8;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       selectReadStageMask_hi_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]       maskForDestination_hi_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_hi = _GEN_8;
  wire [127:0]      regroupV0_hi_lo_lo = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [63:0]       _GEN_9 = {v0_21, v0_20};
  wire [63:0]       regroupV0_hi_lo_hi_lo;
  assign regroupV0_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       regroupV0_hi_lo_hi_lo_9;
  assign regroupV0_hi_lo_hi_lo_9 = _GEN_9;
  wire [63:0]       regroupV0_hi_lo_hi_lo_18;
  assign regroupV0_hi_lo_hi_lo_18 = _GEN_9;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       selectReadStageMask_hi_lo_hi_lo;
  assign selectReadStageMask_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]       maskForDestination_hi_lo_hi_lo;
  assign maskForDestination_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       _GEN_10 = {v0_23, v0_22};
  wire [63:0]       regroupV0_hi_lo_hi_hi;
  assign regroupV0_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       regroupV0_hi_lo_hi_hi_9;
  assign regroupV0_hi_lo_hi_hi_9 = _GEN_10;
  wire [63:0]       regroupV0_hi_lo_hi_hi_18;
  assign regroupV0_hi_lo_hi_hi_18 = _GEN_10;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       selectReadStageMask_hi_lo_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]       maskForDestination_hi_lo_hi_hi;
  assign maskForDestination_hi_lo_hi_hi = _GEN_10;
  wire [127:0]      regroupV0_hi_lo_hi = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [255:0]      regroupV0_hi_lo = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [63:0]       _GEN_11 = {v0_25, v0_24};
  wire [63:0]       regroupV0_hi_hi_lo_lo;
  assign regroupV0_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       regroupV0_hi_hi_lo_lo_9;
  assign regroupV0_hi_hi_lo_lo_9 = _GEN_11;
  wire [63:0]       regroupV0_hi_hi_lo_lo_18;
  assign regroupV0_hi_hi_lo_lo_18 = _GEN_11;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       selectReadStageMask_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]       maskForDestination_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       _GEN_12 = {v0_27, v0_26};
  wire [63:0]       regroupV0_hi_hi_lo_hi;
  assign regroupV0_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       regroupV0_hi_hi_lo_hi_9;
  assign regroupV0_hi_hi_lo_hi_9 = _GEN_12;
  wire [63:0]       regroupV0_hi_hi_lo_hi_18;
  assign regroupV0_hi_hi_lo_hi_18 = _GEN_12;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       selectReadStageMask_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]       maskForDestination_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_lo_hi = _GEN_12;
  wire [127:0]      regroupV0_hi_hi_lo = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [63:0]       _GEN_13 = {v0_29, v0_28};
  wire [63:0]       regroupV0_hi_hi_hi_lo;
  assign regroupV0_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       regroupV0_hi_hi_hi_lo_9;
  assign regroupV0_hi_hi_hi_lo_9 = _GEN_13;
  wire [63:0]       regroupV0_hi_hi_hi_lo_18;
  assign regroupV0_hi_hi_hi_lo_18 = _GEN_13;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       selectReadStageMask_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]       maskForDestination_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       _GEN_14 = {v0_31, v0_30};
  wire [63:0]       regroupV0_hi_hi_hi_hi;
  assign regroupV0_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       regroupV0_hi_hi_hi_hi_9;
  assign regroupV0_hi_hi_hi_hi_9 = _GEN_14;
  wire [63:0]       regroupV0_hi_hi_hi_hi_18;
  assign regroupV0_hi_hi_hi_hi_18 = _GEN_14;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       selectReadStageMask_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]       maskForDestination_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_hi = _GEN_14;
  wire [127:0]      regroupV0_hi_hi_hi = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [255:0]      regroupV0_hi_hi = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [511:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_lo_1 = {regroupV0_lo[35:32], regroupV0_lo[3:0]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_1 = {regroupV0_lo[99:96], regroupV0_lo[67:64]};
  wire [15:0]       regroupV0_lo_lo_lo_1 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [7:0]        regroupV0_lo_lo_hi_lo_1 = {regroupV0_lo[163:160], regroupV0_lo[131:128]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_1 = {regroupV0_lo[227:224], regroupV0_lo[195:192]};
  wire [15:0]       regroupV0_lo_lo_hi_1 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [31:0]       regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_lo_1 = {regroupV0_lo[291:288], regroupV0_lo[259:256]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_1 = {regroupV0_lo[355:352], regroupV0_lo[323:320]};
  wire [15:0]       regroupV0_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [7:0]        regroupV0_lo_hi_hi_lo_1 = {regroupV0_lo[419:416], regroupV0_lo[387:384]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_1 = {regroupV0_lo[483:480], regroupV0_lo[451:448]};
  wire [15:0]       regroupV0_lo_hi_hi_1 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [31:0]       regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [63:0]       regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_lo_1 = {regroupV0_hi[35:32], regroupV0_hi[3:0]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_1 = {regroupV0_hi[99:96], regroupV0_hi[67:64]};
  wire [15:0]       regroupV0_hi_lo_lo_1 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [7:0]        regroupV0_hi_lo_hi_lo_1 = {regroupV0_hi[163:160], regroupV0_hi[131:128]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_1 = {regroupV0_hi[227:224], regroupV0_hi[195:192]};
  wire [15:0]       regroupV0_hi_lo_hi_1 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [31:0]       regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_lo_1 = {regroupV0_hi[291:288], regroupV0_hi[259:256]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_1 = {regroupV0_hi[355:352], regroupV0_hi[323:320]};
  wire [15:0]       regroupV0_hi_hi_lo_1 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [7:0]        regroupV0_hi_hi_hi_lo_1 = {regroupV0_hi[419:416], regroupV0_hi[387:384]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_1 = {regroupV0_hi[483:480], regroupV0_hi[451:448]};
  wire [15:0]       regroupV0_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [31:0]       regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [63:0]       regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo[39:36], regroupV0_lo[7:4]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo[103:100], regroupV0_lo[71:68]};
  wire [15:0]       regroupV0_lo_lo_lo_2 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [7:0]        regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo[167:164], regroupV0_lo[135:132]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo[231:228], regroupV0_lo[199:196]};
  wire [15:0]       regroupV0_lo_lo_hi_2 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [31:0]       regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo[295:292], regroupV0_lo[263:260]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo[359:356], regroupV0_lo[327:324]};
  wire [15:0]       regroupV0_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [7:0]        regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo[423:420], regroupV0_lo[391:388]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo[487:484], regroupV0_lo[455:452]};
  wire [15:0]       regroupV0_lo_hi_hi_2 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [31:0]       regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [63:0]       regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi[39:36], regroupV0_hi[7:4]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi[103:100], regroupV0_hi[71:68]};
  wire [15:0]       regroupV0_hi_lo_lo_2 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [7:0]        regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi[167:164], regroupV0_hi[135:132]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi[231:228], regroupV0_hi[199:196]};
  wire [15:0]       regroupV0_hi_lo_hi_2 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [31:0]       regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi[295:292], regroupV0_hi[263:260]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi[359:356], regroupV0_hi[327:324]};
  wire [15:0]       regroupV0_hi_hi_lo_2 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [7:0]        regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi[423:420], regroupV0_hi[391:388]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi[487:484], regroupV0_hi[455:452]};
  wire [15:0]       regroupV0_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [31:0]       regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [63:0]       regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo[43:40], regroupV0_lo[11:8]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo[107:104], regroupV0_lo[75:72]};
  wire [15:0]       regroupV0_lo_lo_lo_3 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [7:0]        regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo[171:168], regroupV0_lo[139:136]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo[235:232], regroupV0_lo[203:200]};
  wire [15:0]       regroupV0_lo_lo_hi_3 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [31:0]       regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo[299:296], regroupV0_lo[267:264]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo[363:360], regroupV0_lo[331:328]};
  wire [15:0]       regroupV0_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [7:0]        regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo[427:424], regroupV0_lo[395:392]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo[491:488], regroupV0_lo[459:456]};
  wire [15:0]       regroupV0_lo_hi_hi_3 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [31:0]       regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [63:0]       regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi[43:40], regroupV0_hi[11:8]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi[107:104], regroupV0_hi[75:72]};
  wire [15:0]       regroupV0_hi_lo_lo_3 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [7:0]        regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi[171:168], regroupV0_hi[139:136]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi[235:232], regroupV0_hi[203:200]};
  wire [15:0]       regroupV0_hi_lo_hi_3 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [31:0]       regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi[299:296], regroupV0_hi[267:264]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi[363:360], regroupV0_hi[331:328]};
  wire [15:0]       regroupV0_hi_hi_lo_3 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [7:0]        regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi[427:424], regroupV0_hi[395:392]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi[491:488], regroupV0_hi[459:456]};
  wire [15:0]       regroupV0_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [31:0]       regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [63:0]       regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo[47:44], regroupV0_lo[15:12]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo[111:108], regroupV0_lo[79:76]};
  wire [15:0]       regroupV0_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [7:0]        regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo[175:172], regroupV0_lo[143:140]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo[239:236], regroupV0_lo[207:204]};
  wire [15:0]       regroupV0_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [31:0]       regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [7:0]        regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo[303:300], regroupV0_lo[271:268]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo[367:364], regroupV0_lo[335:332]};
  wire [15:0]       regroupV0_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [7:0]        regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo[431:428], regroupV0_lo[399:396]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo[495:492], regroupV0_lo[463:460]};
  wire [15:0]       regroupV0_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [31:0]       regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [63:0]       regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi[47:44], regroupV0_hi[15:12]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi[111:108], regroupV0_hi[79:76]};
  wire [15:0]       regroupV0_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [7:0]        regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi[175:172], regroupV0_hi[143:140]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi[239:236], regroupV0_hi[207:204]};
  wire [15:0]       regroupV0_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [31:0]       regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [7:0]        regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi[303:300], regroupV0_hi[271:268]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi[367:364], regroupV0_hi[335:332]};
  wire [15:0]       regroupV0_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [7:0]        regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi[431:428], regroupV0_hi[399:396]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi[495:492], regroupV0_hi[463:460]};
  wire [15:0]       regroupV0_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [31:0]       regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [63:0]       regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo[51:48], regroupV0_lo[19:16]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo[115:112], regroupV0_lo[83:80]};
  wire [15:0]       regroupV0_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [7:0]        regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo[179:176], regroupV0_lo[147:144]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo[243:240], regroupV0_lo[211:208]};
  wire [15:0]       regroupV0_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [31:0]       regroupV0_lo_lo_5 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [7:0]        regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo[307:304], regroupV0_lo[275:272]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo[371:368], regroupV0_lo[339:336]};
  wire [15:0]       regroupV0_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [7:0]        regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo[435:432], regroupV0_lo[403:400]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo[499:496], regroupV0_lo[467:464]};
  wire [15:0]       regroupV0_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [31:0]       regroupV0_lo_hi_5 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [63:0]       regroupV0_lo_5 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [7:0]        regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi[51:48], regroupV0_hi[19:16]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi[115:112], regroupV0_hi[83:80]};
  wire [15:0]       regroupV0_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [7:0]        regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi[179:176], regroupV0_hi[147:144]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi[243:240], regroupV0_hi[211:208]};
  wire [15:0]       regroupV0_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [31:0]       regroupV0_hi_lo_5 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [7:0]        regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi[307:304], regroupV0_hi[275:272]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi[371:368], regroupV0_hi[339:336]};
  wire [15:0]       regroupV0_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [7:0]        regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi[435:432], regroupV0_hi[403:400]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi[499:496], regroupV0_hi[467:464]};
  wire [15:0]       regroupV0_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [31:0]       regroupV0_hi_hi_5 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [63:0]       regroupV0_hi_5 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo[55:52], regroupV0_lo[23:20]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo[119:116], regroupV0_lo[87:84]};
  wire [15:0]       regroupV0_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [7:0]        regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo[183:180], regroupV0_lo[151:148]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo[247:244], regroupV0_lo[215:212]};
  wire [15:0]       regroupV0_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [31:0]       regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [7:0]        regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo[311:308], regroupV0_lo[279:276]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo[375:372], regroupV0_lo[343:340]};
  wire [15:0]       regroupV0_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [7:0]        regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo[439:436], regroupV0_lo[407:404]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo[503:500], regroupV0_lo[471:468]};
  wire [15:0]       regroupV0_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [31:0]       regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [63:0]       regroupV0_lo_6 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [7:0]        regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi[55:52], regroupV0_hi[23:20]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi[119:116], regroupV0_hi[87:84]};
  wire [15:0]       regroupV0_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [7:0]        regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi[183:180], regroupV0_hi[151:148]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi[247:244], regroupV0_hi[215:212]};
  wire [15:0]       regroupV0_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [31:0]       regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [7:0]        regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi[311:308], regroupV0_hi[279:276]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi[375:372], regroupV0_hi[343:340]};
  wire [15:0]       regroupV0_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [7:0]        regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi[439:436], regroupV0_hi[407:404]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi[503:500], regroupV0_hi[471:468]};
  wire [15:0]       regroupV0_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [31:0]       regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [63:0]       regroupV0_hi_6 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo[59:56], regroupV0_lo[27:24]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo[123:120], regroupV0_lo[91:88]};
  wire [15:0]       regroupV0_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [7:0]        regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo[187:184], regroupV0_lo[155:152]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo[251:248], regroupV0_lo[219:216]};
  wire [15:0]       regroupV0_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [31:0]       regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [7:0]        regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo[315:312], regroupV0_lo[283:280]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo[379:376], regroupV0_lo[347:344]};
  wire [15:0]       regroupV0_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [7:0]        regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo[443:440], regroupV0_lo[411:408]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo[507:504], regroupV0_lo[475:472]};
  wire [15:0]       regroupV0_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [31:0]       regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [63:0]       regroupV0_lo_7 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [7:0]        regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi[59:56], regroupV0_hi[27:24]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi[123:120], regroupV0_hi[91:88]};
  wire [15:0]       regroupV0_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [7:0]        regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi[187:184], regroupV0_hi[155:152]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi[251:248], regroupV0_hi[219:216]};
  wire [15:0]       regroupV0_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [31:0]       regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [7:0]        regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi[315:312], regroupV0_hi[283:280]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi[379:376], regroupV0_hi[347:344]};
  wire [15:0]       regroupV0_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [7:0]        regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi[443:440], regroupV0_hi[411:408]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi[507:504], regroupV0_hi[475:472]};
  wire [15:0]       regroupV0_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [31:0]       regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [63:0]       regroupV0_hi_7 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_lo_lo_8 = {regroupV0_lo[63:60], regroupV0_lo[31:28]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_8 = {regroupV0_lo[127:124], regroupV0_lo[95:92]};
  wire [15:0]       regroupV0_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_8};
  wire [7:0]        regroupV0_lo_lo_hi_lo_8 = {regroupV0_lo[191:188], regroupV0_lo[159:156]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_8 = {regroupV0_lo[255:252], regroupV0_lo[223:220]};
  wire [15:0]       regroupV0_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_8};
  wire [31:0]       regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [7:0]        regroupV0_lo_hi_lo_lo_8 = {regroupV0_lo[319:316], regroupV0_lo[287:284]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_8 = {regroupV0_lo[383:380], regroupV0_lo[351:348]};
  wire [15:0]       regroupV0_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_8};
  wire [7:0]        regroupV0_lo_hi_hi_lo_8 = {regroupV0_lo[447:444], regroupV0_lo[415:412]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_8 = {regroupV0_lo[511:508], regroupV0_lo[479:476]};
  wire [15:0]       regroupV0_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_8};
  wire [31:0]       regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [63:0]       regroupV0_lo_8 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [7:0]        regroupV0_hi_lo_lo_lo_8 = {regroupV0_hi[63:60], regroupV0_hi[31:28]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_8 = {regroupV0_hi[127:124], regroupV0_hi[95:92]};
  wire [15:0]       regroupV0_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_8};
  wire [7:0]        regroupV0_hi_lo_hi_lo_8 = {regroupV0_hi[191:188], regroupV0_hi[159:156]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_8 = {regroupV0_hi[255:252], regroupV0_hi[223:220]};
  wire [15:0]       regroupV0_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_8};
  wire [31:0]       regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [7:0]        regroupV0_hi_hi_lo_lo_8 = {regroupV0_hi[319:316], regroupV0_hi[287:284]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_8 = {regroupV0_hi[383:380], regroupV0_hi[351:348]};
  wire [15:0]       regroupV0_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_8};
  wire [7:0]        regroupV0_hi_hi_hi_lo_8 = {regroupV0_hi[447:444], regroupV0_hi[415:412]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_8 = {regroupV0_hi[511:508], regroupV0_hi[479:476]};
  wire [15:0]       regroupV0_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_8};
  wire [31:0]       regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [63:0]       regroupV0_hi_8 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [255:0]      regroupV0_lo_lo_9 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [255:0]      regroupV0_lo_hi_9 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [511:0]      regroupV0_lo_9 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [255:0]      regroupV0_hi_lo_9 = {regroupV0_hi_6, regroupV0_lo_6, regroupV0_hi_5, regroupV0_lo_5};
  wire [255:0]      regroupV0_hi_hi_9 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [511:0]      regroupV0_hi_9 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [1023:0]     regroupV0_0 = {regroupV0_hi_9, regroupV0_lo_9};
  wire [127:0]      regroupV0_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_9};
  wire [127:0]      regroupV0_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_9};
  wire [255:0]      regroupV0_lo_lo_10 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [127:0]      regroupV0_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_9};
  wire [127:0]      regroupV0_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_9};
  wire [255:0]      regroupV0_lo_hi_10 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [511:0]      regroupV0_lo_10 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [127:0]      regroupV0_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_9};
  wire [127:0]      regroupV0_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_9};
  wire [255:0]      regroupV0_hi_lo_10 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [127:0]      regroupV0_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_9};
  wire [127:0]      regroupV0_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_9};
  wire [255:0]      regroupV0_hi_hi_10 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [511:0]      regroupV0_hi_10 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo = {regroupV0_lo_10[17:16], regroupV0_lo_10[1:0]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi = {regroupV0_lo_10[49:48], regroupV0_lo_10[33:32]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo = {regroupV0_lo_10[81:80], regroupV0_lo_10[65:64]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi = {regroupV0_lo_10[113:112], regroupV0_lo_10[97:96]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [15:0]       regroupV0_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_10};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo = {regroupV0_lo_10[145:144], regroupV0_lo_10[129:128]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi = {regroupV0_lo_10[177:176], regroupV0_lo_10[161:160]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo = {regroupV0_lo_10[209:208], regroupV0_lo_10[193:192]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi = {regroupV0_lo_10[241:240], regroupV0_lo_10[225:224]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [15:0]       regroupV0_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_10};
  wire [31:0]       regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo = {regroupV0_lo_10[273:272], regroupV0_lo_10[257:256]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi = {regroupV0_lo_10[305:304], regroupV0_lo_10[289:288]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo = {regroupV0_lo_10[337:336], regroupV0_lo_10[321:320]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi = {regroupV0_lo_10[369:368], regroupV0_lo_10[353:352]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [15:0]       regroupV0_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_10};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo = {regroupV0_lo_10[401:400], regroupV0_lo_10[385:384]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi = {regroupV0_lo_10[433:432], regroupV0_lo_10[417:416]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo = {regroupV0_lo_10[465:464], regroupV0_lo_10[449:448]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi = {regroupV0_lo_10[497:496], regroupV0_lo_10[481:480]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [15:0]       regroupV0_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_10};
  wire [31:0]       regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [63:0]       regroupV0_lo_11 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo = {regroupV0_hi_10[17:16], regroupV0_hi_10[1:0]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi = {regroupV0_hi_10[49:48], regroupV0_hi_10[33:32]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo = {regroupV0_hi_10[81:80], regroupV0_hi_10[65:64]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi = {regroupV0_hi_10[113:112], regroupV0_hi_10[97:96]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_10 = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [15:0]       regroupV0_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_10};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo = {regroupV0_hi_10[145:144], regroupV0_hi_10[129:128]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi = {regroupV0_hi_10[177:176], regroupV0_hi_10[161:160]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo = {regroupV0_hi_10[209:208], regroupV0_hi_10[193:192]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi = {regroupV0_hi_10[241:240], regroupV0_hi_10[225:224]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [15:0]       regroupV0_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_10};
  wire [31:0]       regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo = {regroupV0_hi_10[273:272], regroupV0_hi_10[257:256]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi = {regroupV0_hi_10[305:304], regroupV0_hi_10[289:288]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_10 = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo = {regroupV0_hi_10[337:336], regroupV0_hi_10[321:320]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi = {regroupV0_hi_10[369:368], regroupV0_hi_10[353:352]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [15:0]       regroupV0_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_10};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo = {regroupV0_hi_10[401:400], regroupV0_hi_10[385:384]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi = {regroupV0_hi_10[433:432], regroupV0_hi_10[417:416]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo = {regroupV0_hi_10[465:464], regroupV0_hi_10[449:448]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi = {regroupV0_hi_10[497:496], regroupV0_hi_10[481:480]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [15:0]       regroupV0_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_10};
  wire [31:0]       regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [63:0]       regroupV0_hi_11 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_1 = {regroupV0_lo_10[19:18], regroupV0_lo_10[3:2]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_1 = {regroupV0_lo_10[51:50], regroupV0_lo_10[35:34]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_1 = {regroupV0_lo_10[83:82], regroupV0_lo_10[67:66]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_1 = {regroupV0_lo_10[115:114], regroupV0_lo_10[99:98]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [15:0]       regroupV0_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_11};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_1 = {regroupV0_lo_10[147:146], regroupV0_lo_10[131:130]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_1 = {regroupV0_lo_10[179:178], regroupV0_lo_10[163:162]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_1 = {regroupV0_lo_10[211:210], regroupV0_lo_10[195:194]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_1 = {regroupV0_lo_10[243:242], regroupV0_lo_10[227:226]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [15:0]       regroupV0_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_11};
  wire [31:0]       regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_1 = {regroupV0_lo_10[275:274], regroupV0_lo_10[259:258]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_1 = {regroupV0_lo_10[307:306], regroupV0_lo_10[291:290]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_1 = {regroupV0_lo_10[339:338], regroupV0_lo_10[323:322]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_1 = {regroupV0_lo_10[371:370], regroupV0_lo_10[355:354]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [15:0]       regroupV0_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_11};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_1 = {regroupV0_lo_10[403:402], regroupV0_lo_10[387:386]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_1 = {regroupV0_lo_10[435:434], regroupV0_lo_10[419:418]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_1 = {regroupV0_lo_10[467:466], regroupV0_lo_10[451:450]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_1 = {regroupV0_lo_10[499:498], regroupV0_lo_10[483:482]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [15:0]       regroupV0_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_11};
  wire [31:0]       regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [63:0]       regroupV0_lo_12 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_1 = {regroupV0_hi_10[19:18], regroupV0_hi_10[3:2]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_1 = {regroupV0_hi_10[51:50], regroupV0_hi_10[35:34]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_1 = {regroupV0_hi_10[83:82], regroupV0_hi_10[67:66]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_1 = {regroupV0_hi_10[115:114], regroupV0_hi_10[99:98]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [15:0]       regroupV0_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_11};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_1 = {regroupV0_hi_10[147:146], regroupV0_hi_10[131:130]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_1 = {regroupV0_hi_10[179:178], regroupV0_hi_10[163:162]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_1 = {regroupV0_hi_10[211:210], regroupV0_hi_10[195:194]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_1 = {regroupV0_hi_10[243:242], regroupV0_hi_10[227:226]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [15:0]       regroupV0_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_11};
  wire [31:0]       regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_1 = {regroupV0_hi_10[275:274], regroupV0_hi_10[259:258]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_1 = {regroupV0_hi_10[307:306], regroupV0_hi_10[291:290]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_1 = {regroupV0_hi_10[339:338], regroupV0_hi_10[323:322]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_1 = {regroupV0_hi_10[371:370], regroupV0_hi_10[355:354]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [15:0]       regroupV0_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_11};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_1 = {regroupV0_hi_10[403:402], regroupV0_hi_10[387:386]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_1 = {regroupV0_hi_10[435:434], regroupV0_hi_10[419:418]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_1 = {regroupV0_hi_10[467:466], regroupV0_hi_10[451:450]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_1 = {regroupV0_hi_10[499:498], regroupV0_hi_10[483:482]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [15:0]       regroupV0_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_11};
  wire [31:0]       regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [63:0]       regroupV0_hi_12 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_2 = {regroupV0_lo_10[21:20], regroupV0_lo_10[5:4]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_2 = {regroupV0_lo_10[53:52], regroupV0_lo_10[37:36]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_2 = {regroupV0_lo_10[85:84], regroupV0_lo_10[69:68]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_2 = {regroupV0_lo_10[117:116], regroupV0_lo_10[101:100]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [15:0]       regroupV0_lo_lo_lo_12 = {regroupV0_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_12};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_2 = {regroupV0_lo_10[149:148], regroupV0_lo_10[133:132]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_2 = {regroupV0_lo_10[181:180], regroupV0_lo_10[165:164]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_12 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_2 = {regroupV0_lo_10[213:212], regroupV0_lo_10[197:196]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_2 = {regroupV0_lo_10[245:244], regroupV0_lo_10[229:228]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [15:0]       regroupV0_lo_lo_hi_12 = {regroupV0_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_12};
  wire [31:0]       regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_12, regroupV0_lo_lo_lo_12};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_2 = {regroupV0_lo_10[277:276], regroupV0_lo_10[261:260]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_2 = {regroupV0_lo_10[309:308], regroupV0_lo_10[293:292]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_12 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_2 = {regroupV0_lo_10[341:340], regroupV0_lo_10[325:324]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_2 = {regroupV0_lo_10[373:372], regroupV0_lo_10[357:356]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_12 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [15:0]       regroupV0_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_12};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_2 = {regroupV0_lo_10[405:404], regroupV0_lo_10[389:388]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_2 = {regroupV0_lo_10[437:436], regroupV0_lo_10[421:420]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_12 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_2 = {regroupV0_lo_10[469:468], regroupV0_lo_10[453:452]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_2 = {regroupV0_lo_10[501:500], regroupV0_lo_10[485:484]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [15:0]       regroupV0_lo_hi_hi_12 = {regroupV0_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_12};
  wire [31:0]       regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_12, regroupV0_lo_hi_lo_12};
  wire [63:0]       regroupV0_lo_13 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_2 = {regroupV0_hi_10[21:20], regroupV0_hi_10[5:4]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_2 = {regroupV0_hi_10[53:52], regroupV0_hi_10[37:36]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_2 = {regroupV0_hi_10[85:84], regroupV0_hi_10[69:68]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_2 = {regroupV0_hi_10[117:116], regroupV0_hi_10[101:100]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_12 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [15:0]       regroupV0_hi_lo_lo_12 = {regroupV0_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_12};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_2 = {regroupV0_hi_10[149:148], regroupV0_hi_10[133:132]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_2 = {regroupV0_hi_10[181:180], regroupV0_hi_10[165:164]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_12 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_2 = {regroupV0_hi_10[213:212], regroupV0_hi_10[197:196]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_2 = {regroupV0_hi_10[245:244], regroupV0_hi_10[229:228]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [15:0]       regroupV0_hi_lo_hi_12 = {regroupV0_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_12};
  wire [31:0]       regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_12, regroupV0_hi_lo_lo_12};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_2 = {regroupV0_hi_10[277:276], regroupV0_hi_10[261:260]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_2 = {regroupV0_hi_10[309:308], regroupV0_hi_10[293:292]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_12 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_2 = {regroupV0_hi_10[341:340], regroupV0_hi_10[325:324]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_2 = {regroupV0_hi_10[373:372], regroupV0_hi_10[357:356]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_12 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [15:0]       regroupV0_hi_hi_lo_12 = {regroupV0_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_12};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_2 = {regroupV0_hi_10[405:404], regroupV0_hi_10[389:388]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_2 = {regroupV0_hi_10[437:436], regroupV0_hi_10[421:420]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_2 = {regroupV0_hi_10[469:468], regroupV0_hi_10[453:452]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_2 = {regroupV0_hi_10[501:500], regroupV0_hi_10[485:484]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [15:0]       regroupV0_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_12};
  wire [31:0]       regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_12, regroupV0_hi_hi_lo_12};
  wire [63:0]       regroupV0_hi_13 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_10[23:22], regroupV0_lo_10[7:6]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_10[55:54], regroupV0_lo_10[39:38]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_10[87:86], regroupV0_lo_10[71:70]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_10[119:118], regroupV0_lo_10[103:102]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [15:0]       regroupV0_lo_lo_lo_13 = {regroupV0_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_13};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_10[151:150], regroupV0_lo_10[135:134]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_10[183:182], regroupV0_lo_10[167:166]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_13 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_10[215:214], regroupV0_lo_10[199:198]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_10[247:246], regroupV0_lo_10[231:230]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [15:0]       regroupV0_lo_lo_hi_13 = {regroupV0_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_13};
  wire [31:0]       regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_13, regroupV0_lo_lo_lo_13};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_10[279:278], regroupV0_lo_10[263:262]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_10[311:310], regroupV0_lo_10[295:294]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_13 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_10[343:342], regroupV0_lo_10[327:326]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_10[375:374], regroupV0_lo_10[359:358]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_13 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [15:0]       regroupV0_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_13};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_10[407:406], regroupV0_lo_10[391:390]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_10[439:438], regroupV0_lo_10[423:422]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_13 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_10[471:470], regroupV0_lo_10[455:454]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_10[503:502], regroupV0_lo_10[487:486]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [15:0]       regroupV0_lo_hi_hi_13 = {regroupV0_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_13};
  wire [31:0]       regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_13, regroupV0_lo_hi_lo_13};
  wire [63:0]       regroupV0_lo_14 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_10[23:22], regroupV0_hi_10[7:6]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_10[55:54], regroupV0_hi_10[39:38]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_10[87:86], regroupV0_hi_10[71:70]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_10[119:118], regroupV0_hi_10[103:102]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_13 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [15:0]       regroupV0_hi_lo_lo_13 = {regroupV0_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_13};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_10[151:150], regroupV0_hi_10[135:134]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_10[183:182], regroupV0_hi_10[167:166]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_13 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_10[215:214], regroupV0_hi_10[199:198]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_10[247:246], regroupV0_hi_10[231:230]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [15:0]       regroupV0_hi_lo_hi_13 = {regroupV0_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_13};
  wire [31:0]       regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_13, regroupV0_hi_lo_lo_13};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_10[279:278], regroupV0_hi_10[263:262]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_10[311:310], regroupV0_hi_10[295:294]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_13 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_10[343:342], regroupV0_hi_10[327:326]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_10[375:374], regroupV0_hi_10[359:358]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_13 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [15:0]       regroupV0_hi_hi_lo_13 = {regroupV0_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_13};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_10[407:406], regroupV0_hi_10[391:390]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_10[439:438], regroupV0_hi_10[423:422]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_10[471:470], regroupV0_hi_10[455:454]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_10[503:502], regroupV0_hi_10[487:486]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [15:0]       regroupV0_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_13};
  wire [31:0]       regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_13, regroupV0_hi_hi_lo_13};
  wire [63:0]       regroupV0_hi_14 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_4 = {regroupV0_lo_10[25:24], regroupV0_lo_10[9:8]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_4 = {regroupV0_lo_10[57:56], regroupV0_lo_10[41:40]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_4};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_4 = {regroupV0_lo_10[89:88], regroupV0_lo_10[73:72]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_4 = {regroupV0_lo_10[121:120], regroupV0_lo_10[105:104]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_4};
  wire [15:0]       regroupV0_lo_lo_lo_14 = {regroupV0_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_14};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_4 = {regroupV0_lo_10[153:152], regroupV0_lo_10[137:136]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_4 = {regroupV0_lo_10[185:184], regroupV0_lo_10[169:168]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_14 = {regroupV0_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_4};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_4 = {regroupV0_lo_10[217:216], regroupV0_lo_10[201:200]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_4 = {regroupV0_lo_10[249:248], regroupV0_lo_10[233:232]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_4};
  wire [15:0]       regroupV0_lo_lo_hi_14 = {regroupV0_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_14};
  wire [31:0]       regroupV0_lo_lo_15 = {regroupV0_lo_lo_hi_14, regroupV0_lo_lo_lo_14};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_4 = {regroupV0_lo_10[281:280], regroupV0_lo_10[265:264]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_4 = {regroupV0_lo_10[313:312], regroupV0_lo_10[297:296]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_14 = {regroupV0_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_4};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_4 = {regroupV0_lo_10[345:344], regroupV0_lo_10[329:328]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_4 = {regroupV0_lo_10[377:376], regroupV0_lo_10[361:360]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_14 = {regroupV0_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_4};
  wire [15:0]       regroupV0_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_14};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_4 = {regroupV0_lo_10[409:408], regroupV0_lo_10[393:392]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_4 = {regroupV0_lo_10[441:440], regroupV0_lo_10[425:424]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_14 = {regroupV0_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_4};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_4 = {regroupV0_lo_10[473:472], regroupV0_lo_10[457:456]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_4 = {regroupV0_lo_10[505:504], regroupV0_lo_10[489:488]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_4};
  wire [15:0]       regroupV0_lo_hi_hi_14 = {regroupV0_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_14};
  wire [31:0]       regroupV0_lo_hi_15 = {regroupV0_lo_hi_hi_14, regroupV0_lo_hi_lo_14};
  wire [63:0]       regroupV0_lo_15 = {regroupV0_lo_hi_15, regroupV0_lo_lo_15};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_4 = {regroupV0_hi_10[25:24], regroupV0_hi_10[9:8]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_4 = {regroupV0_hi_10[57:56], regroupV0_hi_10[41:40]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_4};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_4 = {regroupV0_hi_10[89:88], regroupV0_hi_10[73:72]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_4 = {regroupV0_hi_10[121:120], regroupV0_hi_10[105:104]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_14 = {regroupV0_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_4};
  wire [15:0]       regroupV0_hi_lo_lo_14 = {regroupV0_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_14};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_4 = {regroupV0_hi_10[153:152], regroupV0_hi_10[137:136]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_4 = {regroupV0_hi_10[185:184], regroupV0_hi_10[169:168]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_14 = {regroupV0_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_4};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_4 = {regroupV0_hi_10[217:216], regroupV0_hi_10[201:200]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_4 = {regroupV0_hi_10[249:248], regroupV0_hi_10[233:232]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_4};
  wire [15:0]       regroupV0_hi_lo_hi_14 = {regroupV0_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_14};
  wire [31:0]       regroupV0_hi_lo_15 = {regroupV0_hi_lo_hi_14, regroupV0_hi_lo_lo_14};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_4 = {regroupV0_hi_10[281:280], regroupV0_hi_10[265:264]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_4 = {regroupV0_hi_10[313:312], regroupV0_hi_10[297:296]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_14 = {regroupV0_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_4};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_4 = {regroupV0_hi_10[345:344], regroupV0_hi_10[329:328]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_4 = {regroupV0_hi_10[377:376], regroupV0_hi_10[361:360]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_14 = {regroupV0_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_4};
  wire [15:0]       regroupV0_hi_hi_lo_14 = {regroupV0_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_14};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_4 = {regroupV0_hi_10[409:408], regroupV0_hi_10[393:392]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_4 = {regroupV0_hi_10[441:440], regroupV0_hi_10[425:424]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_4};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_4 = {regroupV0_hi_10[473:472], regroupV0_hi_10[457:456]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_4 = {regroupV0_hi_10[505:504], regroupV0_hi_10[489:488]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_4};
  wire [15:0]       regroupV0_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_14};
  wire [31:0]       regroupV0_hi_hi_15 = {regroupV0_hi_hi_hi_14, regroupV0_hi_hi_lo_14};
  wire [63:0]       regroupV0_hi_15 = {regroupV0_hi_hi_15, regroupV0_hi_lo_15};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_5 = {regroupV0_lo_10[27:26], regroupV0_lo_10[11:10]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_5 = {regroupV0_lo_10[59:58], regroupV0_lo_10[43:42]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_15 = {regroupV0_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_5};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_5 = {regroupV0_lo_10[91:90], regroupV0_lo_10[75:74]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_5 = {regroupV0_lo_10[123:122], regroupV0_lo_10[107:106]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_15 = {regroupV0_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_5};
  wire [15:0]       regroupV0_lo_lo_lo_15 = {regroupV0_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_15};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_5 = {regroupV0_lo_10[155:154], regroupV0_lo_10[139:138]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_5 = {regroupV0_lo_10[187:186], regroupV0_lo_10[171:170]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_15 = {regroupV0_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_5};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_5 = {regroupV0_lo_10[219:218], regroupV0_lo_10[203:202]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_5 = {regroupV0_lo_10[251:250], regroupV0_lo_10[235:234]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_15 = {regroupV0_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_5};
  wire [15:0]       regroupV0_lo_lo_hi_15 = {regroupV0_lo_lo_hi_hi_15, regroupV0_lo_lo_hi_lo_15};
  wire [31:0]       regroupV0_lo_lo_16 = {regroupV0_lo_lo_hi_15, regroupV0_lo_lo_lo_15};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_5 = {regroupV0_lo_10[283:282], regroupV0_lo_10[267:266]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_5 = {regroupV0_lo_10[315:314], regroupV0_lo_10[299:298]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_15 = {regroupV0_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_5};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_5 = {regroupV0_lo_10[347:346], regroupV0_lo_10[331:330]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_5 = {regroupV0_lo_10[379:378], regroupV0_lo_10[363:362]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_15 = {regroupV0_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_5};
  wire [15:0]       regroupV0_lo_hi_lo_15 = {regroupV0_lo_hi_lo_hi_15, regroupV0_lo_hi_lo_lo_15};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_5 = {regroupV0_lo_10[411:410], regroupV0_lo_10[395:394]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_5 = {regroupV0_lo_10[443:442], regroupV0_lo_10[427:426]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_15 = {regroupV0_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_5};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_5 = {regroupV0_lo_10[475:474], regroupV0_lo_10[459:458]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_5 = {regroupV0_lo_10[507:506], regroupV0_lo_10[491:490]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_15 = {regroupV0_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_5};
  wire [15:0]       regroupV0_lo_hi_hi_15 = {regroupV0_lo_hi_hi_hi_15, regroupV0_lo_hi_hi_lo_15};
  wire [31:0]       regroupV0_lo_hi_16 = {regroupV0_lo_hi_hi_15, regroupV0_lo_hi_lo_15};
  wire [63:0]       regroupV0_lo_16 = {regroupV0_lo_hi_16, regroupV0_lo_lo_16};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_5 = {regroupV0_hi_10[27:26], regroupV0_hi_10[11:10]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_5 = {regroupV0_hi_10[59:58], regroupV0_hi_10[43:42]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_15 = {regroupV0_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_5};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_5 = {regroupV0_hi_10[91:90], regroupV0_hi_10[75:74]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_5 = {regroupV0_hi_10[123:122], regroupV0_hi_10[107:106]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_15 = {regroupV0_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_5};
  wire [15:0]       regroupV0_hi_lo_lo_15 = {regroupV0_hi_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_15};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_5 = {regroupV0_hi_10[155:154], regroupV0_hi_10[139:138]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_5 = {regroupV0_hi_10[187:186], regroupV0_hi_10[171:170]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_15 = {regroupV0_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_5};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_5 = {regroupV0_hi_10[219:218], regroupV0_hi_10[203:202]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_5 = {regroupV0_hi_10[251:250], regroupV0_hi_10[235:234]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_15 = {regroupV0_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_5};
  wire [15:0]       regroupV0_hi_lo_hi_15 = {regroupV0_hi_lo_hi_hi_15, regroupV0_hi_lo_hi_lo_15};
  wire [31:0]       regroupV0_hi_lo_16 = {regroupV0_hi_lo_hi_15, regroupV0_hi_lo_lo_15};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_5 = {regroupV0_hi_10[283:282], regroupV0_hi_10[267:266]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_5 = {regroupV0_hi_10[315:314], regroupV0_hi_10[299:298]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_15 = {regroupV0_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_5};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_5 = {regroupV0_hi_10[347:346], regroupV0_hi_10[331:330]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_5 = {regroupV0_hi_10[379:378], regroupV0_hi_10[363:362]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_15 = {regroupV0_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_5};
  wire [15:0]       regroupV0_hi_hi_lo_15 = {regroupV0_hi_hi_lo_hi_15, regroupV0_hi_hi_lo_lo_15};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_5 = {regroupV0_hi_10[411:410], regroupV0_hi_10[395:394]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_5 = {regroupV0_hi_10[443:442], regroupV0_hi_10[427:426]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_15 = {regroupV0_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_5};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_5 = {regroupV0_hi_10[475:474], regroupV0_hi_10[459:458]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_5 = {regroupV0_hi_10[507:506], regroupV0_hi_10[491:490]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_15 = {regroupV0_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_5};
  wire [15:0]       regroupV0_hi_hi_hi_15 = {regroupV0_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_lo_15};
  wire [31:0]       regroupV0_hi_hi_16 = {regroupV0_hi_hi_hi_15, regroupV0_hi_hi_lo_15};
  wire [63:0]       regroupV0_hi_16 = {regroupV0_hi_hi_16, regroupV0_hi_lo_16};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_6 = {regroupV0_lo_10[29:28], regroupV0_lo_10[13:12]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_6 = {regroupV0_lo_10[61:60], regroupV0_lo_10[45:44]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_16 = {regroupV0_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_6};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_6 = {regroupV0_lo_10[93:92], regroupV0_lo_10[77:76]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_6 = {regroupV0_lo_10[125:124], regroupV0_lo_10[109:108]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_16 = {regroupV0_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_6};
  wire [15:0]       regroupV0_lo_lo_lo_16 = {regroupV0_lo_lo_lo_hi_16, regroupV0_lo_lo_lo_lo_16};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_6 = {regroupV0_lo_10[157:156], regroupV0_lo_10[141:140]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_6 = {regroupV0_lo_10[189:188], regroupV0_lo_10[173:172]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_16 = {regroupV0_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_6};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_6 = {regroupV0_lo_10[221:220], regroupV0_lo_10[205:204]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_6 = {regroupV0_lo_10[253:252], regroupV0_lo_10[237:236]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_16 = {regroupV0_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_6};
  wire [15:0]       regroupV0_lo_lo_hi_16 = {regroupV0_lo_lo_hi_hi_16, regroupV0_lo_lo_hi_lo_16};
  wire [31:0]       regroupV0_lo_lo_17 = {regroupV0_lo_lo_hi_16, regroupV0_lo_lo_lo_16};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_6 = {regroupV0_lo_10[285:284], regroupV0_lo_10[269:268]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_6 = {regroupV0_lo_10[317:316], regroupV0_lo_10[301:300]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_16 = {regroupV0_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_6};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_6 = {regroupV0_lo_10[349:348], regroupV0_lo_10[333:332]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_6 = {regroupV0_lo_10[381:380], regroupV0_lo_10[365:364]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_16 = {regroupV0_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_6};
  wire [15:0]       regroupV0_lo_hi_lo_16 = {regroupV0_lo_hi_lo_hi_16, regroupV0_lo_hi_lo_lo_16};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_6 = {regroupV0_lo_10[413:412], regroupV0_lo_10[397:396]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_6 = {regroupV0_lo_10[445:444], regroupV0_lo_10[429:428]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_16 = {regroupV0_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_6};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_6 = {regroupV0_lo_10[477:476], regroupV0_lo_10[461:460]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_6 = {regroupV0_lo_10[509:508], regroupV0_lo_10[493:492]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_16 = {regroupV0_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_6};
  wire [15:0]       regroupV0_lo_hi_hi_16 = {regroupV0_lo_hi_hi_hi_16, regroupV0_lo_hi_hi_lo_16};
  wire [31:0]       regroupV0_lo_hi_17 = {regroupV0_lo_hi_hi_16, regroupV0_lo_hi_lo_16};
  wire [63:0]       regroupV0_lo_17 = {regroupV0_lo_hi_17, regroupV0_lo_lo_17};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_6 = {regroupV0_hi_10[29:28], regroupV0_hi_10[13:12]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_6 = {regroupV0_hi_10[61:60], regroupV0_hi_10[45:44]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_16 = {regroupV0_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_6};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_6 = {regroupV0_hi_10[93:92], regroupV0_hi_10[77:76]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_6 = {regroupV0_hi_10[125:124], regroupV0_hi_10[109:108]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_16 = {regroupV0_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_6};
  wire [15:0]       regroupV0_hi_lo_lo_16 = {regroupV0_hi_lo_lo_hi_16, regroupV0_hi_lo_lo_lo_16};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_6 = {regroupV0_hi_10[157:156], regroupV0_hi_10[141:140]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_6 = {regroupV0_hi_10[189:188], regroupV0_hi_10[173:172]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_16 = {regroupV0_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_6};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_6 = {regroupV0_hi_10[221:220], regroupV0_hi_10[205:204]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_6 = {regroupV0_hi_10[253:252], regroupV0_hi_10[237:236]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_16 = {regroupV0_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_6};
  wire [15:0]       regroupV0_hi_lo_hi_16 = {regroupV0_hi_lo_hi_hi_16, regroupV0_hi_lo_hi_lo_16};
  wire [31:0]       regroupV0_hi_lo_17 = {regroupV0_hi_lo_hi_16, regroupV0_hi_lo_lo_16};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_6 = {regroupV0_hi_10[285:284], regroupV0_hi_10[269:268]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_6 = {regroupV0_hi_10[317:316], regroupV0_hi_10[301:300]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_16 = {regroupV0_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_6};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_6 = {regroupV0_hi_10[349:348], regroupV0_hi_10[333:332]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_6 = {regroupV0_hi_10[381:380], regroupV0_hi_10[365:364]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_16 = {regroupV0_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_6};
  wire [15:0]       regroupV0_hi_hi_lo_16 = {regroupV0_hi_hi_lo_hi_16, regroupV0_hi_hi_lo_lo_16};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_6 = {regroupV0_hi_10[413:412], regroupV0_hi_10[397:396]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_6 = {regroupV0_hi_10[445:444], regroupV0_hi_10[429:428]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_16 = {regroupV0_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_6};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_6 = {regroupV0_hi_10[477:476], regroupV0_hi_10[461:460]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_6 = {regroupV0_hi_10[509:508], regroupV0_hi_10[493:492]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_16 = {regroupV0_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_6};
  wire [15:0]       regroupV0_hi_hi_hi_16 = {regroupV0_hi_hi_hi_hi_16, regroupV0_hi_hi_hi_lo_16};
  wire [31:0]       regroupV0_hi_hi_17 = {regroupV0_hi_hi_hi_16, regroupV0_hi_hi_lo_16};
  wire [63:0]       regroupV0_hi_17 = {regroupV0_hi_hi_17, regroupV0_hi_lo_17};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_7 = {regroupV0_lo_10[31:30], regroupV0_lo_10[15:14]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_7 = {regroupV0_lo_10[63:62], regroupV0_lo_10[47:46]};
  wire [7:0]        regroupV0_lo_lo_lo_lo_17 = {regroupV0_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_7};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_7 = {regroupV0_lo_10[95:94], regroupV0_lo_10[79:78]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_7 = {regroupV0_lo_10[127:126], regroupV0_lo_10[111:110]};
  wire [7:0]        regroupV0_lo_lo_lo_hi_17 = {regroupV0_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_7};
  wire [15:0]       regroupV0_lo_lo_lo_17 = {regroupV0_lo_lo_lo_hi_17, regroupV0_lo_lo_lo_lo_17};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_7 = {regroupV0_lo_10[159:158], regroupV0_lo_10[143:142]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_7 = {regroupV0_lo_10[191:190], regroupV0_lo_10[175:174]};
  wire [7:0]        regroupV0_lo_lo_hi_lo_17 = {regroupV0_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_7};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_7 = {regroupV0_lo_10[223:222], regroupV0_lo_10[207:206]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_7 = {regroupV0_lo_10[255:254], regroupV0_lo_10[239:238]};
  wire [7:0]        regroupV0_lo_lo_hi_hi_17 = {regroupV0_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_7};
  wire [15:0]       regroupV0_lo_lo_hi_17 = {regroupV0_lo_lo_hi_hi_17, regroupV0_lo_lo_hi_lo_17};
  wire [31:0]       regroupV0_lo_lo_18 = {regroupV0_lo_lo_hi_17, regroupV0_lo_lo_lo_17};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_7 = {regroupV0_lo_10[287:286], regroupV0_lo_10[271:270]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_7 = {regroupV0_lo_10[319:318], regroupV0_lo_10[303:302]};
  wire [7:0]        regroupV0_lo_hi_lo_lo_17 = {regroupV0_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_7};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_7 = {regroupV0_lo_10[351:350], regroupV0_lo_10[335:334]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_7 = {regroupV0_lo_10[383:382], regroupV0_lo_10[367:366]};
  wire [7:0]        regroupV0_lo_hi_lo_hi_17 = {regroupV0_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_7};
  wire [15:0]       regroupV0_lo_hi_lo_17 = {regroupV0_lo_hi_lo_hi_17, regroupV0_lo_hi_lo_lo_17};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_7 = {regroupV0_lo_10[415:414], regroupV0_lo_10[399:398]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_7 = {regroupV0_lo_10[447:446], regroupV0_lo_10[431:430]};
  wire [7:0]        regroupV0_lo_hi_hi_lo_17 = {regroupV0_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_7};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_7 = {regroupV0_lo_10[479:478], regroupV0_lo_10[463:462]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_7 = {regroupV0_lo_10[511:510], regroupV0_lo_10[495:494]};
  wire [7:0]        regroupV0_lo_hi_hi_hi_17 = {regroupV0_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_7};
  wire [15:0]       regroupV0_lo_hi_hi_17 = {regroupV0_lo_hi_hi_hi_17, regroupV0_lo_hi_hi_lo_17};
  wire [31:0]       regroupV0_lo_hi_18 = {regroupV0_lo_hi_hi_17, regroupV0_lo_hi_lo_17};
  wire [63:0]       regroupV0_lo_18 = {regroupV0_lo_hi_18, regroupV0_lo_lo_18};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_7 = {regroupV0_hi_10[31:30], regroupV0_hi_10[15:14]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_7 = {regroupV0_hi_10[63:62], regroupV0_hi_10[47:46]};
  wire [7:0]        regroupV0_hi_lo_lo_lo_17 = {regroupV0_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_7};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_7 = {regroupV0_hi_10[95:94], regroupV0_hi_10[79:78]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_7 = {regroupV0_hi_10[127:126], regroupV0_hi_10[111:110]};
  wire [7:0]        regroupV0_hi_lo_lo_hi_17 = {regroupV0_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_7};
  wire [15:0]       regroupV0_hi_lo_lo_17 = {regroupV0_hi_lo_lo_hi_17, regroupV0_hi_lo_lo_lo_17};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_7 = {regroupV0_hi_10[159:158], regroupV0_hi_10[143:142]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_7 = {regroupV0_hi_10[191:190], regroupV0_hi_10[175:174]};
  wire [7:0]        regroupV0_hi_lo_hi_lo_17 = {regroupV0_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_7};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_7 = {regroupV0_hi_10[223:222], regroupV0_hi_10[207:206]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_7 = {regroupV0_hi_10[255:254], regroupV0_hi_10[239:238]};
  wire [7:0]        regroupV0_hi_lo_hi_hi_17 = {regroupV0_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_7};
  wire [15:0]       regroupV0_hi_lo_hi_17 = {regroupV0_hi_lo_hi_hi_17, regroupV0_hi_lo_hi_lo_17};
  wire [31:0]       regroupV0_hi_lo_18 = {regroupV0_hi_lo_hi_17, regroupV0_hi_lo_lo_17};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_7 = {regroupV0_hi_10[287:286], regroupV0_hi_10[271:270]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_7 = {regroupV0_hi_10[319:318], regroupV0_hi_10[303:302]};
  wire [7:0]        regroupV0_hi_hi_lo_lo_17 = {regroupV0_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_7};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_7 = {regroupV0_hi_10[351:350], regroupV0_hi_10[335:334]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_7 = {regroupV0_hi_10[383:382], regroupV0_hi_10[367:366]};
  wire [7:0]        regroupV0_hi_hi_lo_hi_17 = {regroupV0_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_7};
  wire [15:0]       regroupV0_hi_hi_lo_17 = {regroupV0_hi_hi_lo_hi_17, regroupV0_hi_hi_lo_lo_17};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_7 = {regroupV0_hi_10[415:414], regroupV0_hi_10[399:398]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_7 = {regroupV0_hi_10[447:446], regroupV0_hi_10[431:430]};
  wire [7:0]        regroupV0_hi_hi_hi_lo_17 = {regroupV0_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_7};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_7 = {regroupV0_hi_10[479:478], regroupV0_hi_10[463:462]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_7 = {regroupV0_hi_10[511:510], regroupV0_hi_10[495:494]};
  wire [7:0]        regroupV0_hi_hi_hi_hi_17 = {regroupV0_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_7};
  wire [15:0]       regroupV0_hi_hi_hi_17 = {regroupV0_hi_hi_hi_hi_17, regroupV0_hi_hi_hi_lo_17};
  wire [31:0]       regroupV0_hi_hi_18 = {regroupV0_hi_hi_hi_17, regroupV0_hi_hi_lo_17};
  wire [63:0]       regroupV0_hi_18 = {regroupV0_hi_hi_18, regroupV0_hi_lo_18};
  wire [255:0]      regroupV0_lo_lo_19 = {regroupV0_hi_12, regroupV0_lo_12, regroupV0_hi_11, regroupV0_lo_11};
  wire [255:0]      regroupV0_lo_hi_19 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [511:0]      regroupV0_lo_19 = {regroupV0_lo_hi_19, regroupV0_lo_lo_19};
  wire [255:0]      regroupV0_hi_lo_19 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [255:0]      regroupV0_hi_hi_19 = {regroupV0_hi_18, regroupV0_lo_18, regroupV0_hi_17, regroupV0_lo_17};
  wire [511:0]      regroupV0_hi_19 = {regroupV0_hi_hi_19, regroupV0_hi_lo_19};
  wire [1023:0]     regroupV0_1 = {regroupV0_hi_19, regroupV0_lo_19};
  wire [127:0]      regroupV0_lo_lo_lo_18 = {regroupV0_lo_lo_lo_hi_18, regroupV0_lo_lo_lo_lo_18};
  wire [127:0]      regroupV0_lo_lo_hi_18 = {regroupV0_lo_lo_hi_hi_18, regroupV0_lo_lo_hi_lo_18};
  wire [255:0]      regroupV0_lo_lo_20 = {regroupV0_lo_lo_hi_18, regroupV0_lo_lo_lo_18};
  wire [127:0]      regroupV0_lo_hi_lo_18 = {regroupV0_lo_hi_lo_hi_18, regroupV0_lo_hi_lo_lo_18};
  wire [127:0]      regroupV0_lo_hi_hi_18 = {regroupV0_lo_hi_hi_hi_18, regroupV0_lo_hi_hi_lo_18};
  wire [255:0]      regroupV0_lo_hi_20 = {regroupV0_lo_hi_hi_18, regroupV0_lo_hi_lo_18};
  wire [511:0]      regroupV0_lo_20 = {regroupV0_lo_hi_20, regroupV0_lo_lo_20};
  wire [127:0]      regroupV0_hi_lo_lo_18 = {regroupV0_hi_lo_lo_hi_18, regroupV0_hi_lo_lo_lo_18};
  wire [127:0]      regroupV0_hi_lo_hi_18 = {regroupV0_hi_lo_hi_hi_18, regroupV0_hi_lo_hi_lo_18};
  wire [255:0]      regroupV0_hi_lo_20 = {regroupV0_hi_lo_hi_18, regroupV0_hi_lo_lo_18};
  wire [127:0]      regroupV0_hi_hi_lo_18 = {regroupV0_hi_hi_lo_hi_18, regroupV0_hi_hi_lo_lo_18};
  wire [127:0]      regroupV0_hi_hi_hi_18 = {regroupV0_hi_hi_hi_hi_18, regroupV0_hi_hi_hi_lo_18};
  wire [255:0]      regroupV0_hi_hi_20 = {regroupV0_hi_hi_hi_18, regroupV0_hi_hi_lo_18};
  wire [511:0]      regroupV0_hi_20 = {regroupV0_hi_hi_20, regroupV0_hi_lo_20};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo = {regroupV0_lo_20[8], regroupV0_lo_20[0]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi = {regroupV0_lo_20[24], regroupV0_lo_20[16]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo = {regroupV0_lo_20[40], regroupV0_lo_20[32]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi = {regroupV0_lo_20[56], regroupV0_lo_20[48]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_lo_19 = {regroupV0_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_8};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo = {regroupV0_lo_20[72], regroupV0_lo_20[64]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi = {regroupV0_lo_20[88], regroupV0_lo_20[80]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo = {regroupV0_lo_20[104], regroupV0_lo_20[96]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi = {regroupV0_lo_20[120], regroupV0_lo_20[112]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_hi_19 = {regroupV0_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_8};
  wire [15:0]       regroupV0_lo_lo_lo_19 = {regroupV0_lo_lo_lo_hi_19, regroupV0_lo_lo_lo_lo_19};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo = {regroupV0_lo_20[136], regroupV0_lo_20[128]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi = {regroupV0_lo_20[152], regroupV0_lo_20[144]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo = {regroupV0_lo_20[168], regroupV0_lo_20[160]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi = {regroupV0_lo_20[184], regroupV0_lo_20[176]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo};
  wire [7:0]        regroupV0_lo_lo_hi_lo_19 = {regroupV0_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_8};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo = {regroupV0_lo_20[200], regroupV0_lo_20[192]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi = {regroupV0_lo_20[216], regroupV0_lo_20[208]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo = {regroupV0_lo_20[232], regroupV0_lo_20[224]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi = {regroupV0_lo_20[248], regroupV0_lo_20[240]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo};
  wire [7:0]        regroupV0_lo_lo_hi_hi_19 = {regroupV0_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_8};
  wire [15:0]       regroupV0_lo_lo_hi_19 = {regroupV0_lo_lo_hi_hi_19, regroupV0_lo_lo_hi_lo_19};
  wire [31:0]       regroupV0_lo_lo_21 = {regroupV0_lo_lo_hi_19, regroupV0_lo_lo_lo_19};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo = {regroupV0_lo_20[264], regroupV0_lo_20[256]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi = {regroupV0_lo_20[280], regroupV0_lo_20[272]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo = {regroupV0_lo_20[296], regroupV0_lo_20[288]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi = {regroupV0_lo_20[312], regroupV0_lo_20[304]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo};
  wire [7:0]        regroupV0_lo_hi_lo_lo_19 = {regroupV0_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_8};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo = {regroupV0_lo_20[328], regroupV0_lo_20[320]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi = {regroupV0_lo_20[344], regroupV0_lo_20[336]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo = {regroupV0_lo_20[360], regroupV0_lo_20[352]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi = {regroupV0_lo_20[376], regroupV0_lo_20[368]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo};
  wire [7:0]        regroupV0_lo_hi_lo_hi_19 = {regroupV0_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_8};
  wire [15:0]       regroupV0_lo_hi_lo_19 = {regroupV0_lo_hi_lo_hi_19, regroupV0_lo_hi_lo_lo_19};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo = {regroupV0_lo_20[392], regroupV0_lo_20[384]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi = {regroupV0_lo_20[408], regroupV0_lo_20[400]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo = {regroupV0_lo_20[424], regroupV0_lo_20[416]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi = {regroupV0_lo_20[440], regroupV0_lo_20[432]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo};
  wire [7:0]        regroupV0_lo_hi_hi_lo_19 = {regroupV0_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_8};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo = {regroupV0_lo_20[456], regroupV0_lo_20[448]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi = {regroupV0_lo_20[472], regroupV0_lo_20[464]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo = {regroupV0_lo_20[488], regroupV0_lo_20[480]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi = {regroupV0_lo_20[504], regroupV0_lo_20[496]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo};
  wire [7:0]        regroupV0_lo_hi_hi_hi_19 = {regroupV0_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_8};
  wire [15:0]       regroupV0_lo_hi_hi_19 = {regroupV0_lo_hi_hi_hi_19, regroupV0_lo_hi_hi_lo_19};
  wire [31:0]       regroupV0_lo_hi_21 = {regroupV0_lo_hi_hi_19, regroupV0_lo_hi_lo_19};
  wire [63:0]       regroupV0_lo_21 = {regroupV0_lo_hi_21, regroupV0_lo_lo_21};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo = {regroupV0_hi_20[8], regroupV0_hi_20[0]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi = {regroupV0_hi_20[24], regroupV0_hi_20[16]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo = {regroupV0_hi_20[40], regroupV0_hi_20[32]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi = {regroupV0_hi_20[56], regroupV0_hi_20[48]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo};
  wire [7:0]        regroupV0_hi_lo_lo_lo_19 = {regroupV0_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_8};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo = {regroupV0_hi_20[72], regroupV0_hi_20[64]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi = {regroupV0_hi_20[88], regroupV0_hi_20[80]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo = {regroupV0_hi_20[104], regroupV0_hi_20[96]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi = {regroupV0_hi_20[120], regroupV0_hi_20[112]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo};
  wire [7:0]        regroupV0_hi_lo_lo_hi_19 = {regroupV0_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_8};
  wire [15:0]       regroupV0_hi_lo_lo_19 = {regroupV0_hi_lo_lo_hi_19, regroupV0_hi_lo_lo_lo_19};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo = {regroupV0_hi_20[136], regroupV0_hi_20[128]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi = {regroupV0_hi_20[152], regroupV0_hi_20[144]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo = {regroupV0_hi_20[168], regroupV0_hi_20[160]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi = {regroupV0_hi_20[184], regroupV0_hi_20[176]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo};
  wire [7:0]        regroupV0_hi_lo_hi_lo_19 = {regroupV0_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_8};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo = {regroupV0_hi_20[200], regroupV0_hi_20[192]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi = {regroupV0_hi_20[216], regroupV0_hi_20[208]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo = {regroupV0_hi_20[232], regroupV0_hi_20[224]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi = {regroupV0_hi_20[248], regroupV0_hi_20[240]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo};
  wire [7:0]        regroupV0_hi_lo_hi_hi_19 = {regroupV0_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_8};
  wire [15:0]       regroupV0_hi_lo_hi_19 = {regroupV0_hi_lo_hi_hi_19, regroupV0_hi_lo_hi_lo_19};
  wire [31:0]       regroupV0_hi_lo_21 = {regroupV0_hi_lo_hi_19, regroupV0_hi_lo_lo_19};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo = {regroupV0_hi_20[264], regroupV0_hi_20[256]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi = {regroupV0_hi_20[280], regroupV0_hi_20[272]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo = {regroupV0_hi_20[296], regroupV0_hi_20[288]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi = {regroupV0_hi_20[312], regroupV0_hi_20[304]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo};
  wire [7:0]        regroupV0_hi_hi_lo_lo_19 = {regroupV0_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_8};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo = {regroupV0_hi_20[328], regroupV0_hi_20[320]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi = {regroupV0_hi_20[344], regroupV0_hi_20[336]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo = {regroupV0_hi_20[360], regroupV0_hi_20[352]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi = {regroupV0_hi_20[376], regroupV0_hi_20[368]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo};
  wire [7:0]        regroupV0_hi_hi_lo_hi_19 = {regroupV0_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_8};
  wire [15:0]       regroupV0_hi_hi_lo_19 = {regroupV0_hi_hi_lo_hi_19, regroupV0_hi_hi_lo_lo_19};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo = {regroupV0_hi_20[392], regroupV0_hi_20[384]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi = {regroupV0_hi_20[408], regroupV0_hi_20[400]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo = {regroupV0_hi_20[424], regroupV0_hi_20[416]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi = {regroupV0_hi_20[440], regroupV0_hi_20[432]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo};
  wire [7:0]        regroupV0_hi_hi_hi_lo_19 = {regroupV0_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_8};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo = {regroupV0_hi_20[456], regroupV0_hi_20[448]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi = {regroupV0_hi_20[472], regroupV0_hi_20[464]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo = {regroupV0_hi_20[488], regroupV0_hi_20[480]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi = {regroupV0_hi_20[504], regroupV0_hi_20[496]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo};
  wire [7:0]        regroupV0_hi_hi_hi_hi_19 = {regroupV0_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_8};
  wire [15:0]       regroupV0_hi_hi_hi_19 = {regroupV0_hi_hi_hi_hi_19, regroupV0_hi_hi_hi_lo_19};
  wire [31:0]       regroupV0_hi_hi_21 = {regroupV0_hi_hi_hi_19, regroupV0_hi_hi_lo_19};
  wire [63:0]       regroupV0_hi_21 = {regroupV0_hi_hi_21, regroupV0_hi_lo_21};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_20[9], regroupV0_lo_20[1]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_20[25], regroupV0_lo_20[17]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_20[41], regroupV0_lo_20[33]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_20[57], regroupV0_lo_20[49]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_lo_20 = {regroupV0_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_9};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_20[73], regroupV0_lo_20[65]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_20[89], regroupV0_lo_20[81]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_20[105], regroupV0_lo_20[97]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_20[121], regroupV0_lo_20[113]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_hi_20 = {regroupV0_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_9};
  wire [15:0]       regroupV0_lo_lo_lo_20 = {regroupV0_lo_lo_lo_hi_20, regroupV0_lo_lo_lo_lo_20};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_20[137], regroupV0_lo_20[129]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_20[153], regroupV0_lo_20[145]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_20[169], regroupV0_lo_20[161]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_20[185], regroupV0_lo_20[177]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_hi_lo_20 = {regroupV0_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_9};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_20[201], regroupV0_lo_20[193]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_20[217], regroupV0_lo_20[209]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_20[233], regroupV0_lo_20[225]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_20[249], regroupV0_lo_20[241]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_hi_hi_20 = {regroupV0_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_9};
  wire [15:0]       regroupV0_lo_lo_hi_20 = {regroupV0_lo_lo_hi_hi_20, regroupV0_lo_lo_hi_lo_20};
  wire [31:0]       regroupV0_lo_lo_22 = {regroupV0_lo_lo_hi_20, regroupV0_lo_lo_lo_20};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_20[265], regroupV0_lo_20[257]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_20[281], regroupV0_lo_20[273]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_20[297], regroupV0_lo_20[289]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_20[313], regroupV0_lo_20[305]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_lo_20 = {regroupV0_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_9};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_20[329], regroupV0_lo_20[321]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_20[345], regroupV0_lo_20[337]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_20[361], regroupV0_lo_20[353]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_20[377], regroupV0_lo_20[369]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_hi_20 = {regroupV0_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_9};
  wire [15:0]       regroupV0_lo_hi_lo_20 = {regroupV0_lo_hi_lo_hi_20, regroupV0_lo_hi_lo_lo_20};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_20[393], regroupV0_lo_20[385]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_20[409], regroupV0_lo_20[401]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_20[425], regroupV0_lo_20[417]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_20[441], regroupV0_lo_20[433]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_hi_lo_20 = {regroupV0_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_9};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_20[457], regroupV0_lo_20[449]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_20[473], regroupV0_lo_20[465]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_20[489], regroupV0_lo_20[481]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_20[505], regroupV0_lo_20[497]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_hi_hi_20 = {regroupV0_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_9};
  wire [15:0]       regroupV0_lo_hi_hi_20 = {regroupV0_lo_hi_hi_hi_20, regroupV0_lo_hi_hi_lo_20};
  wire [31:0]       regroupV0_lo_hi_22 = {regroupV0_lo_hi_hi_20, regroupV0_lo_hi_lo_20};
  wire [63:0]       regroupV0_lo_22 = {regroupV0_lo_hi_22, regroupV0_lo_lo_22};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_20[9], regroupV0_hi_20[1]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_20[25], regroupV0_hi_20[17]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_20[41], regroupV0_hi_20[33]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_20[57], regroupV0_hi_20[49]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_lo_20 = {regroupV0_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_9};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_20[73], regroupV0_hi_20[65]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_20[89], regroupV0_hi_20[81]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_20[105], regroupV0_hi_20[97]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_20[121], regroupV0_hi_20[113]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_hi_20 = {regroupV0_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_9};
  wire [15:0]       regroupV0_hi_lo_lo_20 = {regroupV0_hi_lo_lo_hi_20, regroupV0_hi_lo_lo_lo_20};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_20[137], regroupV0_hi_20[129]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_20[153], regroupV0_hi_20[145]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_20[169], regroupV0_hi_20[161]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_20[185], regroupV0_hi_20[177]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_hi_lo_20 = {regroupV0_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_9};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_20[201], regroupV0_hi_20[193]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_20[217], regroupV0_hi_20[209]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_20[233], regroupV0_hi_20[225]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_20[249], regroupV0_hi_20[241]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_hi_hi_20 = {regroupV0_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_9};
  wire [15:0]       regroupV0_hi_lo_hi_20 = {regroupV0_hi_lo_hi_hi_20, regroupV0_hi_lo_hi_lo_20};
  wire [31:0]       regroupV0_hi_lo_22 = {regroupV0_hi_lo_hi_20, regroupV0_hi_lo_lo_20};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_20[265], regroupV0_hi_20[257]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_20[281], regroupV0_hi_20[273]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_20[297], regroupV0_hi_20[289]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_20[313], regroupV0_hi_20[305]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_lo_20 = {regroupV0_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_9};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_20[329], regroupV0_hi_20[321]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_20[345], regroupV0_hi_20[337]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_20[361], regroupV0_hi_20[353]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_20[377], regroupV0_hi_20[369]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_hi_20 = {regroupV0_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_9};
  wire [15:0]       regroupV0_hi_hi_lo_20 = {regroupV0_hi_hi_lo_hi_20, regroupV0_hi_hi_lo_lo_20};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_20[393], regroupV0_hi_20[385]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_20[409], regroupV0_hi_20[401]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_20[425], regroupV0_hi_20[417]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_20[441], regroupV0_hi_20[433]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_hi_lo_20 = {regroupV0_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_9};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_20[457], regroupV0_hi_20[449]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_20[473], regroupV0_hi_20[465]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_20[489], regroupV0_hi_20[481]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_20[505], regroupV0_hi_20[497]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_hi_hi_20 = {regroupV0_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_9};
  wire [15:0]       regroupV0_hi_hi_hi_20 = {regroupV0_hi_hi_hi_hi_20, regroupV0_hi_hi_hi_lo_20};
  wire [31:0]       regroupV0_hi_hi_22 = {regroupV0_hi_hi_hi_20, regroupV0_hi_hi_lo_20};
  wire [63:0]       regroupV0_hi_22 = {regroupV0_hi_hi_22, regroupV0_hi_lo_22};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_20[10], regroupV0_lo_20[2]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_20[26], regroupV0_lo_20[18]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_20[42], regroupV0_lo_20[34]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_20[58], regroupV0_lo_20[50]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_lo_21 = {regroupV0_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_10};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_20[74], regroupV0_lo_20[66]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_20[90], regroupV0_lo_20[82]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_20[106], regroupV0_lo_20[98]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_20[122], regroupV0_lo_20[114]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_hi_21 = {regroupV0_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_10};
  wire [15:0]       regroupV0_lo_lo_lo_21 = {regroupV0_lo_lo_lo_hi_21, regroupV0_lo_lo_lo_lo_21};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_20[138], regroupV0_lo_20[130]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_20[154], regroupV0_lo_20[146]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_20[170], regroupV0_lo_20[162]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_20[186], regroupV0_lo_20[178]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_hi_lo_21 = {regroupV0_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_10};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_20[202], regroupV0_lo_20[194]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_20[218], regroupV0_lo_20[210]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_20[234], regroupV0_lo_20[226]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_20[250], regroupV0_lo_20[242]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_hi_hi_21 = {regroupV0_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_10};
  wire [15:0]       regroupV0_lo_lo_hi_21 = {regroupV0_lo_lo_hi_hi_21, regroupV0_lo_lo_hi_lo_21};
  wire [31:0]       regroupV0_lo_lo_23 = {regroupV0_lo_lo_hi_21, regroupV0_lo_lo_lo_21};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_20[266], regroupV0_lo_20[258]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_20[282], regroupV0_lo_20[274]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_20[298], regroupV0_lo_20[290]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_20[314], regroupV0_lo_20[306]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_lo_21 = {regroupV0_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_10};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_20[330], regroupV0_lo_20[322]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_20[346], regroupV0_lo_20[338]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_20[362], regroupV0_lo_20[354]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_20[378], regroupV0_lo_20[370]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_hi_21 = {regroupV0_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_10};
  wire [15:0]       regroupV0_lo_hi_lo_21 = {regroupV0_lo_hi_lo_hi_21, regroupV0_lo_hi_lo_lo_21};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_20[394], regroupV0_lo_20[386]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_20[410], regroupV0_lo_20[402]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_20[426], regroupV0_lo_20[418]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_20[442], regroupV0_lo_20[434]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_hi_lo_21 = {regroupV0_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_10};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_20[458], regroupV0_lo_20[450]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_20[474], regroupV0_lo_20[466]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_20[490], regroupV0_lo_20[482]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_20[506], regroupV0_lo_20[498]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_hi_hi_21 = {regroupV0_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_10};
  wire [15:0]       regroupV0_lo_hi_hi_21 = {regroupV0_lo_hi_hi_hi_21, regroupV0_lo_hi_hi_lo_21};
  wire [31:0]       regroupV0_lo_hi_23 = {regroupV0_lo_hi_hi_21, regroupV0_lo_hi_lo_21};
  wire [63:0]       regroupV0_lo_23 = {regroupV0_lo_hi_23, regroupV0_lo_lo_23};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_20[10], regroupV0_hi_20[2]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_20[26], regroupV0_hi_20[18]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_20[42], regroupV0_hi_20[34]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_20[58], regroupV0_hi_20[50]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_lo_21 = {regroupV0_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_10};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_20[74], regroupV0_hi_20[66]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_20[90], regroupV0_hi_20[82]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_20[106], regroupV0_hi_20[98]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_20[122], regroupV0_hi_20[114]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_hi_21 = {regroupV0_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_10};
  wire [15:0]       regroupV0_hi_lo_lo_21 = {regroupV0_hi_lo_lo_hi_21, regroupV0_hi_lo_lo_lo_21};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_20[138], regroupV0_hi_20[130]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_20[154], regroupV0_hi_20[146]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_20[170], regroupV0_hi_20[162]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_20[186], regroupV0_hi_20[178]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_hi_lo_21 = {regroupV0_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_10};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_20[202], regroupV0_hi_20[194]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_20[218], regroupV0_hi_20[210]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_20[234], regroupV0_hi_20[226]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_20[250], regroupV0_hi_20[242]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_hi_hi_21 = {regroupV0_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_10};
  wire [15:0]       regroupV0_hi_lo_hi_21 = {regroupV0_hi_lo_hi_hi_21, regroupV0_hi_lo_hi_lo_21};
  wire [31:0]       regroupV0_hi_lo_23 = {regroupV0_hi_lo_hi_21, regroupV0_hi_lo_lo_21};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_20[266], regroupV0_hi_20[258]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_20[282], regroupV0_hi_20[274]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_20[298], regroupV0_hi_20[290]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_20[314], regroupV0_hi_20[306]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_lo_21 = {regroupV0_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_10};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_20[330], regroupV0_hi_20[322]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_20[346], regroupV0_hi_20[338]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_20[362], regroupV0_hi_20[354]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_20[378], regroupV0_hi_20[370]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_hi_21 = {regroupV0_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_10};
  wire [15:0]       regroupV0_hi_hi_lo_21 = {regroupV0_hi_hi_lo_hi_21, regroupV0_hi_hi_lo_lo_21};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_20[394], regroupV0_hi_20[386]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_20[410], regroupV0_hi_20[402]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_20[426], regroupV0_hi_20[418]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_20[442], regroupV0_hi_20[434]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_hi_lo_21 = {regroupV0_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_10};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_20[458], regroupV0_hi_20[450]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_20[474], regroupV0_hi_20[466]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_20[490], regroupV0_hi_20[482]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_20[506], regroupV0_hi_20[498]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_hi_hi_21 = {regroupV0_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_10};
  wire [15:0]       regroupV0_hi_hi_hi_21 = {regroupV0_hi_hi_hi_hi_21, regroupV0_hi_hi_hi_lo_21};
  wire [31:0]       regroupV0_hi_hi_23 = {regroupV0_hi_hi_hi_21, regroupV0_hi_hi_lo_21};
  wire [63:0]       regroupV0_hi_23 = {regroupV0_hi_hi_23, regroupV0_hi_lo_23};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_20[11], regroupV0_lo_20[3]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_20[27], regroupV0_lo_20[19]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_20[43], regroupV0_lo_20[35]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_20[59], regroupV0_lo_20[51]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_lo_22 = {regroupV0_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_11};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_20[75], regroupV0_lo_20[67]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_20[91], regroupV0_lo_20[83]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_20[107], regroupV0_lo_20[99]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_20[123], regroupV0_lo_20[115]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_hi_22 = {regroupV0_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_11};
  wire [15:0]       regroupV0_lo_lo_lo_22 = {regroupV0_lo_lo_lo_hi_22, regroupV0_lo_lo_lo_lo_22};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_20[139], regroupV0_lo_20[131]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_20[155], regroupV0_lo_20[147]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_20[171], regroupV0_lo_20[163]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_20[187], regroupV0_lo_20[179]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_hi_lo_22 = {regroupV0_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_11};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_20[203], regroupV0_lo_20[195]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_20[219], regroupV0_lo_20[211]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_20[235], regroupV0_lo_20[227]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_20[251], regroupV0_lo_20[243]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_hi_hi_22 = {regroupV0_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_11};
  wire [15:0]       regroupV0_lo_lo_hi_22 = {regroupV0_lo_lo_hi_hi_22, regroupV0_lo_lo_hi_lo_22};
  wire [31:0]       regroupV0_lo_lo_24 = {regroupV0_lo_lo_hi_22, regroupV0_lo_lo_lo_22};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_20[267], regroupV0_lo_20[259]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_20[283], regroupV0_lo_20[275]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_20[299], regroupV0_lo_20[291]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_20[315], regroupV0_lo_20[307]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_lo_22 = {regroupV0_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_11};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_20[331], regroupV0_lo_20[323]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_20[347], regroupV0_lo_20[339]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_20[363], regroupV0_lo_20[355]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_20[379], regroupV0_lo_20[371]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_hi_22 = {regroupV0_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_11};
  wire [15:0]       regroupV0_lo_hi_lo_22 = {regroupV0_lo_hi_lo_hi_22, regroupV0_lo_hi_lo_lo_22};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_20[395], regroupV0_lo_20[387]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_20[411], regroupV0_lo_20[403]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_20[427], regroupV0_lo_20[419]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_20[443], regroupV0_lo_20[435]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_hi_lo_22 = {regroupV0_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_11};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_20[459], regroupV0_lo_20[451]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_20[475], regroupV0_lo_20[467]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_20[491], regroupV0_lo_20[483]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_20[507], regroupV0_lo_20[499]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_hi_hi_22 = {regroupV0_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_11};
  wire [15:0]       regroupV0_lo_hi_hi_22 = {regroupV0_lo_hi_hi_hi_22, regroupV0_lo_hi_hi_lo_22};
  wire [31:0]       regroupV0_lo_hi_24 = {regroupV0_lo_hi_hi_22, regroupV0_lo_hi_lo_22};
  wire [63:0]       regroupV0_lo_24 = {regroupV0_lo_hi_24, regroupV0_lo_lo_24};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_20[11], regroupV0_hi_20[3]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_20[27], regroupV0_hi_20[19]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_20[43], regroupV0_hi_20[35]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_20[59], regroupV0_hi_20[51]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_lo_22 = {regroupV0_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_11};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_20[75], regroupV0_hi_20[67]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_20[91], regroupV0_hi_20[83]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_20[107], regroupV0_hi_20[99]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_20[123], regroupV0_hi_20[115]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_hi_22 = {regroupV0_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_11};
  wire [15:0]       regroupV0_hi_lo_lo_22 = {regroupV0_hi_lo_lo_hi_22, regroupV0_hi_lo_lo_lo_22};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_20[139], regroupV0_hi_20[131]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_20[155], regroupV0_hi_20[147]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_20[171], regroupV0_hi_20[163]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_20[187], regroupV0_hi_20[179]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_hi_lo_22 = {regroupV0_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_11};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_20[203], regroupV0_hi_20[195]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_20[219], regroupV0_hi_20[211]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_20[235], regroupV0_hi_20[227]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_20[251], regroupV0_hi_20[243]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_hi_hi_22 = {regroupV0_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_11};
  wire [15:0]       regroupV0_hi_lo_hi_22 = {regroupV0_hi_lo_hi_hi_22, regroupV0_hi_lo_hi_lo_22};
  wire [31:0]       regroupV0_hi_lo_24 = {regroupV0_hi_lo_hi_22, regroupV0_hi_lo_lo_22};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_20[267], regroupV0_hi_20[259]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_20[283], regroupV0_hi_20[275]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_20[299], regroupV0_hi_20[291]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_20[315], regroupV0_hi_20[307]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_lo_22 = {regroupV0_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_11};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_20[331], regroupV0_hi_20[323]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_20[347], regroupV0_hi_20[339]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_20[363], regroupV0_hi_20[355]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_20[379], regroupV0_hi_20[371]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_hi_22 = {regroupV0_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_11};
  wire [15:0]       regroupV0_hi_hi_lo_22 = {regroupV0_hi_hi_lo_hi_22, regroupV0_hi_hi_lo_lo_22};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_20[395], regroupV0_hi_20[387]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_20[411], regroupV0_hi_20[403]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_20[427], regroupV0_hi_20[419]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_20[443], regroupV0_hi_20[435]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_hi_lo_22 = {regroupV0_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_11};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_20[459], regroupV0_hi_20[451]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_20[475], regroupV0_hi_20[467]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_20[491], regroupV0_hi_20[483]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_20[507], regroupV0_hi_20[499]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_hi_hi_22 = {regroupV0_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_11};
  wire [15:0]       regroupV0_hi_hi_hi_22 = {regroupV0_hi_hi_hi_hi_22, regroupV0_hi_hi_hi_lo_22};
  wire [31:0]       regroupV0_hi_hi_24 = {regroupV0_hi_hi_hi_22, regroupV0_hi_hi_lo_22};
  wire [63:0]       regroupV0_hi_24 = {regroupV0_hi_hi_24, regroupV0_hi_lo_24};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_20[12], regroupV0_lo_20[4]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_20[28], regroupV0_lo_20[20]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_20[44], regroupV0_lo_20[36]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_20[60], regroupV0_lo_20[52]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_lo_lo_23 = {regroupV0_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_12};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_20[76], regroupV0_lo_20[68]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_20[92], regroupV0_lo_20[84]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_12 = {regroupV0_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_20[108], regroupV0_lo_20[100]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_20[124], regroupV0_lo_20[116]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_12 = {regroupV0_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_lo_hi_23 = {regroupV0_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_12};
  wire [15:0]       regroupV0_lo_lo_lo_23 = {regroupV0_lo_lo_lo_hi_23, regroupV0_lo_lo_lo_lo_23};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_20[140], regroupV0_lo_20[132]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_20[156], regroupV0_lo_20[148]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_12 = {regroupV0_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_20[172], regroupV0_lo_20[164]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_20[188], regroupV0_lo_20[180]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_12 = {regroupV0_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_hi_lo_23 = {regroupV0_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_12};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_20[204], regroupV0_lo_20[196]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_20[220], regroupV0_lo_20[212]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_12 = {regroupV0_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_20[236], regroupV0_lo_20[228]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_20[252], regroupV0_lo_20[244]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_hi_hi_23 = {regroupV0_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_12};
  wire [15:0]       regroupV0_lo_lo_hi_23 = {regroupV0_lo_lo_hi_hi_23, regroupV0_lo_lo_hi_lo_23};
  wire [31:0]       regroupV0_lo_lo_25 = {regroupV0_lo_lo_hi_23, regroupV0_lo_lo_lo_23};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_20[268], regroupV0_lo_20[260]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_20[284], regroupV0_lo_20[276]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_12 = {regroupV0_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_20[300], regroupV0_lo_20[292]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_20[316], regroupV0_lo_20[308]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_12 = {regroupV0_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_lo_lo_23 = {regroupV0_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_12};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_20[332], regroupV0_lo_20[324]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_20[348], regroupV0_lo_20[340]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_20[364], regroupV0_lo_20[356]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_20[380], regroupV0_lo_20[372]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_12 = {regroupV0_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_lo_hi_23 = {regroupV0_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_12};
  wire [15:0]       regroupV0_lo_hi_lo_23 = {regroupV0_lo_hi_lo_hi_23, regroupV0_lo_hi_lo_lo_23};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_20[396], regroupV0_lo_20[388]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_20[412], regroupV0_lo_20[404]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_12 = {regroupV0_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_20[428], regroupV0_lo_20[420]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_20[444], regroupV0_lo_20[436]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_12 = {regroupV0_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_hi_lo_23 = {regroupV0_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_12};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_20[460], regroupV0_lo_20[452]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_20[476], regroupV0_lo_20[468]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_12 = {regroupV0_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_20[492], regroupV0_lo_20[484]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_20[508], regroupV0_lo_20[500]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_hi_hi_23 = {regroupV0_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_12};
  wire [15:0]       regroupV0_lo_hi_hi_23 = {regroupV0_lo_hi_hi_hi_23, regroupV0_lo_hi_hi_lo_23};
  wire [31:0]       regroupV0_lo_hi_25 = {regroupV0_lo_hi_hi_23, regroupV0_lo_hi_lo_23};
  wire [63:0]       regroupV0_lo_25 = {regroupV0_lo_hi_25, regroupV0_lo_lo_25};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_20[12], regroupV0_hi_20[4]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_20[28], regroupV0_hi_20[20]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_20[44], regroupV0_hi_20[36]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_20[60], regroupV0_hi_20[52]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_12 = {regroupV0_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_lo_23 = {regroupV0_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_12};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_20[76], regroupV0_hi_20[68]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_20[92], regroupV0_hi_20[84]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_12 = {regroupV0_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_20[108], regroupV0_hi_20[100]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_20[124], regroupV0_hi_20[116]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_12 = {regroupV0_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_hi_23 = {regroupV0_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_12};
  wire [15:0]       regroupV0_hi_lo_lo_23 = {regroupV0_hi_lo_lo_hi_23, regroupV0_hi_lo_lo_lo_23};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_20[140], regroupV0_hi_20[132]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_20[156], regroupV0_hi_20[148]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_12 = {regroupV0_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_20[172], regroupV0_hi_20[164]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_20[188], regroupV0_hi_20[180]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_12 = {regroupV0_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_hi_lo_23 = {regroupV0_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_12};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_20[204], regroupV0_hi_20[196]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_20[220], regroupV0_hi_20[212]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_12 = {regroupV0_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_20[236], regroupV0_hi_20[228]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_20[252], regroupV0_hi_20[244]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_hi_hi_23 = {regroupV0_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_12};
  wire [15:0]       regroupV0_hi_lo_hi_23 = {regroupV0_hi_lo_hi_hi_23, regroupV0_hi_lo_hi_lo_23};
  wire [31:0]       regroupV0_hi_lo_25 = {regroupV0_hi_lo_hi_23, regroupV0_hi_lo_lo_23};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_20[268], regroupV0_hi_20[260]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_20[284], regroupV0_hi_20[276]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_12 = {regroupV0_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_20[300], regroupV0_hi_20[292]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_20[316], regroupV0_hi_20[308]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_12 = {regroupV0_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_lo_lo_23 = {regroupV0_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_12};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_20[332], regroupV0_hi_20[324]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_20[348], regroupV0_hi_20[340]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_12 = {regroupV0_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_20[364], regroupV0_hi_20[356]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_20[380], regroupV0_hi_20[372]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_12 = {regroupV0_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_lo_hi_23 = {regroupV0_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_12};
  wire [15:0]       regroupV0_hi_hi_lo_23 = {regroupV0_hi_hi_lo_hi_23, regroupV0_hi_hi_lo_lo_23};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_20[396], regroupV0_hi_20[388]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_20[412], regroupV0_hi_20[404]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_12 = {regroupV0_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_20[428], regroupV0_hi_20[420]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_20[444], regroupV0_hi_20[436]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_12 = {regroupV0_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_hi_lo_23 = {regroupV0_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_12};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_20[460], regroupV0_hi_20[452]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_20[476], regroupV0_hi_20[468]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_20[492], regroupV0_hi_20[484]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_20[508], regroupV0_hi_20[500]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_hi_hi_23 = {regroupV0_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_12};
  wire [15:0]       regroupV0_hi_hi_hi_23 = {regroupV0_hi_hi_hi_hi_23, regroupV0_hi_hi_hi_lo_23};
  wire [31:0]       regroupV0_hi_hi_25 = {regroupV0_hi_hi_hi_23, regroupV0_hi_hi_lo_23};
  wire [63:0]       regroupV0_hi_25 = {regroupV0_hi_hi_25, regroupV0_hi_lo_25};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_20[13], regroupV0_lo_20[5]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_20[29], regroupV0_lo_20[21]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_20[45], regroupV0_lo_20[37]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_20[61], regroupV0_lo_20[53]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_lo_lo_24 = {regroupV0_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_13};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_20[77], regroupV0_lo_20[69]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_20[93], regroupV0_lo_20[85]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_13 = {regroupV0_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_20[109], regroupV0_lo_20[101]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_20[125], regroupV0_lo_20[117]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_13 = {regroupV0_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_lo_hi_24 = {regroupV0_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_13};
  wire [15:0]       regroupV0_lo_lo_lo_24 = {regroupV0_lo_lo_lo_hi_24, regroupV0_lo_lo_lo_lo_24};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_20[141], regroupV0_lo_20[133]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_20[157], regroupV0_lo_20[149]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_13 = {regroupV0_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_20[173], regroupV0_lo_20[165]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_20[189], regroupV0_lo_20[181]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_13 = {regroupV0_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_hi_lo_24 = {regroupV0_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_13};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_20[205], regroupV0_lo_20[197]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_20[221], regroupV0_lo_20[213]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_13 = {regroupV0_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_20[237], regroupV0_lo_20[229]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_20[253], regroupV0_lo_20[245]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_hi_hi_24 = {regroupV0_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_13};
  wire [15:0]       regroupV0_lo_lo_hi_24 = {regroupV0_lo_lo_hi_hi_24, regroupV0_lo_lo_hi_lo_24};
  wire [31:0]       regroupV0_lo_lo_26 = {regroupV0_lo_lo_hi_24, regroupV0_lo_lo_lo_24};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_20[269], regroupV0_lo_20[261]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_20[285], regroupV0_lo_20[277]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_13 = {regroupV0_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_20[301], regroupV0_lo_20[293]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_20[317], regroupV0_lo_20[309]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_13 = {regroupV0_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_lo_lo_24 = {regroupV0_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_13};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_20[333], regroupV0_lo_20[325]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_20[349], regroupV0_lo_20[341]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_20[365], regroupV0_lo_20[357]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_20[381], regroupV0_lo_20[373]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_13 = {regroupV0_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_lo_hi_24 = {regroupV0_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_13};
  wire [15:0]       regroupV0_lo_hi_lo_24 = {regroupV0_lo_hi_lo_hi_24, regroupV0_lo_hi_lo_lo_24};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_20[397], regroupV0_lo_20[389]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_20[413], regroupV0_lo_20[405]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_13 = {regroupV0_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_20[429], regroupV0_lo_20[421]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_20[445], regroupV0_lo_20[437]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_13 = {regroupV0_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_hi_lo_24 = {regroupV0_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_13};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_20[461], regroupV0_lo_20[453]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_20[477], regroupV0_lo_20[469]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_13 = {regroupV0_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_20[493], regroupV0_lo_20[485]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_20[509], regroupV0_lo_20[501]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_hi_hi_24 = {regroupV0_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_13};
  wire [15:0]       regroupV0_lo_hi_hi_24 = {regroupV0_lo_hi_hi_hi_24, regroupV0_lo_hi_hi_lo_24};
  wire [31:0]       regroupV0_lo_hi_26 = {regroupV0_lo_hi_hi_24, regroupV0_lo_hi_lo_24};
  wire [63:0]       regroupV0_lo_26 = {regroupV0_lo_hi_26, regroupV0_lo_lo_26};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_20[13], regroupV0_hi_20[5]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_20[29], regroupV0_hi_20[21]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_20[45], regroupV0_hi_20[37]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_20[61], regroupV0_hi_20[53]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_13 = {regroupV0_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_lo_lo_24 = {regroupV0_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_13};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_20[77], regroupV0_hi_20[69]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_20[93], regroupV0_hi_20[85]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_13 = {regroupV0_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_20[109], regroupV0_hi_20[101]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_20[125], regroupV0_hi_20[117]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_13 = {regroupV0_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_lo_hi_24 = {regroupV0_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_13};
  wire [15:0]       regroupV0_hi_lo_lo_24 = {regroupV0_hi_lo_lo_hi_24, regroupV0_hi_lo_lo_lo_24};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_20[141], regroupV0_hi_20[133]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_20[157], regroupV0_hi_20[149]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_13 = {regroupV0_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_20[173], regroupV0_hi_20[165]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_20[189], regroupV0_hi_20[181]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_13 = {regroupV0_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_hi_lo_24 = {regroupV0_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_13};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_20[205], regroupV0_hi_20[197]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_20[221], regroupV0_hi_20[213]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_13 = {regroupV0_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_20[237], regroupV0_hi_20[229]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_20[253], regroupV0_hi_20[245]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_hi_hi_24 = {regroupV0_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_13};
  wire [15:0]       regroupV0_hi_lo_hi_24 = {regroupV0_hi_lo_hi_hi_24, regroupV0_hi_lo_hi_lo_24};
  wire [31:0]       regroupV0_hi_lo_26 = {regroupV0_hi_lo_hi_24, regroupV0_hi_lo_lo_24};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_20[269], regroupV0_hi_20[261]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_20[285], regroupV0_hi_20[277]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_13 = {regroupV0_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_20[301], regroupV0_hi_20[293]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_20[317], regroupV0_hi_20[309]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_13 = {regroupV0_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_lo_lo_24 = {regroupV0_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_13};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_20[333], regroupV0_hi_20[325]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_20[349], regroupV0_hi_20[341]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_13 = {regroupV0_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_20[365], regroupV0_hi_20[357]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_20[381], regroupV0_hi_20[373]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_13 = {regroupV0_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_lo_hi_24 = {regroupV0_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_13};
  wire [15:0]       regroupV0_hi_hi_lo_24 = {regroupV0_hi_hi_lo_hi_24, regroupV0_hi_hi_lo_lo_24};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_20[397], regroupV0_hi_20[389]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_20[413], regroupV0_hi_20[405]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_13 = {regroupV0_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_20[429], regroupV0_hi_20[421]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_20[445], regroupV0_hi_20[437]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_13 = {regroupV0_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_hi_lo_24 = {regroupV0_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_13};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_20[461], regroupV0_hi_20[453]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_20[477], regroupV0_hi_20[469]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_20[493], regroupV0_hi_20[485]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_20[509], regroupV0_hi_20[501]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_hi_hi_24 = {regroupV0_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_13};
  wire [15:0]       regroupV0_hi_hi_hi_24 = {regroupV0_hi_hi_hi_hi_24, regroupV0_hi_hi_hi_lo_24};
  wire [31:0]       regroupV0_hi_hi_26 = {regroupV0_hi_hi_hi_24, regroupV0_hi_hi_lo_24};
  wire [63:0]       regroupV0_hi_26 = {regroupV0_hi_hi_26, regroupV0_hi_lo_26};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_20[14], regroupV0_lo_20[6]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_20[30], regroupV0_lo_20[22]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_20[46], regroupV0_lo_20[38]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_20[62], regroupV0_lo_20[54]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_lo_lo_25 = {regroupV0_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_14};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_20[78], regroupV0_lo_20[70]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_20[94], regroupV0_lo_20[86]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_14 = {regroupV0_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_20[110], regroupV0_lo_20[102]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_20[126], regroupV0_lo_20[118]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_14 = {regroupV0_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_lo_hi_25 = {regroupV0_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_14};
  wire [15:0]       regroupV0_lo_lo_lo_25 = {regroupV0_lo_lo_lo_hi_25, regroupV0_lo_lo_lo_lo_25};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_20[142], regroupV0_lo_20[134]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_20[158], regroupV0_lo_20[150]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_14 = {regroupV0_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_20[174], regroupV0_lo_20[166]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_20[190], regroupV0_lo_20[182]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_14 = {regroupV0_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_hi_lo_25 = {regroupV0_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_14};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_20[206], regroupV0_lo_20[198]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_20[222], regroupV0_lo_20[214]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_14 = {regroupV0_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_20[238], regroupV0_lo_20[230]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_20[254], regroupV0_lo_20[246]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_hi_hi_25 = {regroupV0_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_14};
  wire [15:0]       regroupV0_lo_lo_hi_25 = {regroupV0_lo_lo_hi_hi_25, regroupV0_lo_lo_hi_lo_25};
  wire [31:0]       regroupV0_lo_lo_27 = {regroupV0_lo_lo_hi_25, regroupV0_lo_lo_lo_25};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_20[270], regroupV0_lo_20[262]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_20[286], regroupV0_lo_20[278]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_14 = {regroupV0_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_20[302], regroupV0_lo_20[294]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_20[318], regroupV0_lo_20[310]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_14 = {regroupV0_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_lo_lo_25 = {regroupV0_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_14};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_20[334], regroupV0_lo_20[326]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_20[350], regroupV0_lo_20[342]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_20[366], regroupV0_lo_20[358]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_20[382], regroupV0_lo_20[374]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_14 = {regroupV0_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_lo_hi_25 = {regroupV0_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_14};
  wire [15:0]       regroupV0_lo_hi_lo_25 = {regroupV0_lo_hi_lo_hi_25, regroupV0_lo_hi_lo_lo_25};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_20[398], regroupV0_lo_20[390]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_20[414], regroupV0_lo_20[406]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_14 = {regroupV0_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_20[430], regroupV0_lo_20[422]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_20[446], regroupV0_lo_20[438]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_14 = {regroupV0_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_hi_lo_25 = {regroupV0_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_14};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_20[462], regroupV0_lo_20[454]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_20[478], regroupV0_lo_20[470]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_14 = {regroupV0_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_20[494], regroupV0_lo_20[486]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_20[510], regroupV0_lo_20[502]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_hi_hi_25 = {regroupV0_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_14};
  wire [15:0]       regroupV0_lo_hi_hi_25 = {regroupV0_lo_hi_hi_hi_25, regroupV0_lo_hi_hi_lo_25};
  wire [31:0]       regroupV0_lo_hi_27 = {regroupV0_lo_hi_hi_25, regroupV0_lo_hi_lo_25};
  wire [63:0]       regroupV0_lo_27 = {regroupV0_lo_hi_27, regroupV0_lo_lo_27};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_20[14], regroupV0_hi_20[6]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_20[30], regroupV0_hi_20[22]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_20[46], regroupV0_hi_20[38]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_20[62], regroupV0_hi_20[54]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_14 = {regroupV0_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_lo_lo_25 = {regroupV0_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_14};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_20[78], regroupV0_hi_20[70]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_20[94], regroupV0_hi_20[86]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_14 = {regroupV0_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_20[110], regroupV0_hi_20[102]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_20[126], regroupV0_hi_20[118]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_14 = {regroupV0_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_lo_hi_25 = {regroupV0_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_14};
  wire [15:0]       regroupV0_hi_lo_lo_25 = {regroupV0_hi_lo_lo_hi_25, regroupV0_hi_lo_lo_lo_25};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_20[142], regroupV0_hi_20[134]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_20[158], regroupV0_hi_20[150]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_14 = {regroupV0_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_20[174], regroupV0_hi_20[166]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_20[190], regroupV0_hi_20[182]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_14 = {regroupV0_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_hi_lo_25 = {regroupV0_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_14};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_20[206], regroupV0_hi_20[198]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_20[222], regroupV0_hi_20[214]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_14 = {regroupV0_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_20[238], regroupV0_hi_20[230]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_20[254], regroupV0_hi_20[246]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_hi_hi_25 = {regroupV0_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_14};
  wire [15:0]       regroupV0_hi_lo_hi_25 = {regroupV0_hi_lo_hi_hi_25, regroupV0_hi_lo_hi_lo_25};
  wire [31:0]       regroupV0_hi_lo_27 = {regroupV0_hi_lo_hi_25, regroupV0_hi_lo_lo_25};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_20[270], regroupV0_hi_20[262]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_20[286], regroupV0_hi_20[278]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_14 = {regroupV0_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_20[302], regroupV0_hi_20[294]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_20[318], regroupV0_hi_20[310]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_14 = {regroupV0_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_lo_lo_25 = {regroupV0_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_14};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_20[334], regroupV0_hi_20[326]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_20[350], regroupV0_hi_20[342]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_14 = {regroupV0_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_20[366], regroupV0_hi_20[358]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_20[382], regroupV0_hi_20[374]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_14 = {regroupV0_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_lo_hi_25 = {regroupV0_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_14};
  wire [15:0]       regroupV0_hi_hi_lo_25 = {regroupV0_hi_hi_lo_hi_25, regroupV0_hi_hi_lo_lo_25};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_20[398], regroupV0_hi_20[390]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_20[414], regroupV0_hi_20[406]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_14 = {regroupV0_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_20[430], regroupV0_hi_20[422]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_20[446], regroupV0_hi_20[438]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_14 = {regroupV0_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_hi_lo_25 = {regroupV0_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_14};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_20[462], regroupV0_hi_20[454]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_20[478], regroupV0_hi_20[470]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_20[494], regroupV0_hi_20[486]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_20[510], regroupV0_hi_20[502]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_hi_hi_25 = {regroupV0_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_14};
  wire [15:0]       regroupV0_hi_hi_hi_25 = {regroupV0_hi_hi_hi_hi_25, regroupV0_hi_hi_hi_lo_25};
  wire [31:0]       regroupV0_hi_hi_27 = {regroupV0_hi_hi_hi_25, regroupV0_hi_hi_lo_25};
  wire [63:0]       regroupV0_hi_27 = {regroupV0_hi_hi_27, regroupV0_hi_lo_27};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_20[15], regroupV0_lo_20[7]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_20[31], regroupV0_lo_20[23]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_lo_15 = {regroupV0_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_20[47], regroupV0_lo_20[39]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_20[63], regroupV0_lo_20[55]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_hi_15 = {regroupV0_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_lo_lo_26 = {regroupV0_lo_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_lo_15};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_20[79], regroupV0_lo_20[71]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_20[95], regroupV0_lo_20[87]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_lo_15 = {regroupV0_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_20[111], regroupV0_lo_20[103]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_20[127], regroupV0_lo_20[119]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_hi_15 = {regroupV0_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_lo_hi_26 = {regroupV0_lo_lo_lo_hi_hi_15, regroupV0_lo_lo_lo_hi_lo_15};
  wire [15:0]       regroupV0_lo_lo_lo_26 = {regroupV0_lo_lo_lo_hi_26, regroupV0_lo_lo_lo_lo_26};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_20[143], regroupV0_lo_20[135]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_20[159], regroupV0_lo_20[151]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_lo_15 = {regroupV0_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_20[175], regroupV0_lo_20[167]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_20[191], regroupV0_lo_20[183]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_hi_15 = {regroupV0_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_hi_lo_26 = {regroupV0_lo_lo_hi_lo_hi_15, regroupV0_lo_lo_hi_lo_lo_15};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_20[207], regroupV0_lo_20[199]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_20[223], regroupV0_lo_20[215]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_lo_15 = {regroupV0_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_20[239], regroupV0_lo_20[231]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_20[255], regroupV0_lo_20[247]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_hi_15 = {regroupV0_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_hi_hi_26 = {regroupV0_lo_lo_hi_hi_hi_15, regroupV0_lo_lo_hi_hi_lo_15};
  wire [15:0]       regroupV0_lo_lo_hi_26 = {regroupV0_lo_lo_hi_hi_26, regroupV0_lo_lo_hi_lo_26};
  wire [31:0]       regroupV0_lo_lo_28 = {regroupV0_lo_lo_hi_26, regroupV0_lo_lo_lo_26};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_20[271], regroupV0_lo_20[263]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_20[287], regroupV0_lo_20[279]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_lo_15 = {regroupV0_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_20[303], regroupV0_lo_20[295]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_20[319], regroupV0_lo_20[311]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_hi_15 = {regroupV0_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_lo_lo_26 = {regroupV0_lo_hi_lo_lo_hi_15, regroupV0_lo_hi_lo_lo_lo_15};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_20[335], regroupV0_lo_20[327]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_20[351], regroupV0_lo_20[343]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_lo_15 = {regroupV0_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_20[367], regroupV0_lo_20[359]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_20[383], regroupV0_lo_20[375]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_hi_15 = {regroupV0_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_lo_hi_26 = {regroupV0_lo_hi_lo_hi_hi_15, regroupV0_lo_hi_lo_hi_lo_15};
  wire [15:0]       regroupV0_lo_hi_lo_26 = {regroupV0_lo_hi_lo_hi_26, regroupV0_lo_hi_lo_lo_26};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_20[399], regroupV0_lo_20[391]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_20[415], regroupV0_lo_20[407]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_lo_15 = {regroupV0_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_20[431], regroupV0_lo_20[423]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_20[447], regroupV0_lo_20[439]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_hi_15 = {regroupV0_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_hi_lo_26 = {regroupV0_lo_hi_hi_lo_hi_15, regroupV0_lo_hi_hi_lo_lo_15};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_20[463], regroupV0_lo_20[455]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_20[479], regroupV0_lo_20[471]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_lo_15 = {regroupV0_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_20[495], regroupV0_lo_20[487]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_20[511], regroupV0_lo_20[503]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_hi_15 = {regroupV0_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_hi_hi_26 = {regroupV0_lo_hi_hi_hi_hi_15, regroupV0_lo_hi_hi_hi_lo_15};
  wire [15:0]       regroupV0_lo_hi_hi_26 = {regroupV0_lo_hi_hi_hi_26, regroupV0_lo_hi_hi_lo_26};
  wire [31:0]       regroupV0_lo_hi_28 = {regroupV0_lo_hi_hi_26, regroupV0_lo_hi_lo_26};
  wire [63:0]       regroupV0_lo_28 = {regroupV0_lo_hi_28, regroupV0_lo_lo_28};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_20[15], regroupV0_hi_20[7]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_20[31], regroupV0_hi_20[23]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_lo_15 = {regroupV0_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_20[47], regroupV0_hi_20[39]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_20[63], regroupV0_hi_20[55]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_hi_15 = {regroupV0_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_lo_lo_26 = {regroupV0_hi_lo_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_lo_15};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_20[79], regroupV0_hi_20[71]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_20[95], regroupV0_hi_20[87]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_lo_15 = {regroupV0_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_20[111], regroupV0_hi_20[103]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_20[127], regroupV0_hi_20[119]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_hi_15 = {regroupV0_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_lo_hi_26 = {regroupV0_hi_lo_lo_hi_hi_15, regroupV0_hi_lo_lo_hi_lo_15};
  wire [15:0]       regroupV0_hi_lo_lo_26 = {regroupV0_hi_lo_lo_hi_26, regroupV0_hi_lo_lo_lo_26};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_20[143], regroupV0_hi_20[135]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_20[159], regroupV0_hi_20[151]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_lo_15 = {regroupV0_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_20[175], regroupV0_hi_20[167]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_20[191], regroupV0_hi_20[183]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_hi_15 = {regroupV0_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_hi_lo_26 = {regroupV0_hi_lo_hi_lo_hi_15, regroupV0_hi_lo_hi_lo_lo_15};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_20[207], regroupV0_hi_20[199]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_20[223], regroupV0_hi_20[215]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_lo_15 = {regroupV0_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_20[239], regroupV0_hi_20[231]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_20[255], regroupV0_hi_20[247]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_hi_15 = {regroupV0_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_hi_hi_26 = {regroupV0_hi_lo_hi_hi_hi_15, regroupV0_hi_lo_hi_hi_lo_15};
  wire [15:0]       regroupV0_hi_lo_hi_26 = {regroupV0_hi_lo_hi_hi_26, regroupV0_hi_lo_hi_lo_26};
  wire [31:0]       regroupV0_hi_lo_28 = {regroupV0_hi_lo_hi_26, regroupV0_hi_lo_lo_26};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_20[271], regroupV0_hi_20[263]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_20[287], regroupV0_hi_20[279]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_lo_15 = {regroupV0_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_20[303], regroupV0_hi_20[295]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_20[319], regroupV0_hi_20[311]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_hi_15 = {regroupV0_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_lo_lo_26 = {regroupV0_hi_hi_lo_lo_hi_15, regroupV0_hi_hi_lo_lo_lo_15};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_20[335], regroupV0_hi_20[327]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_20[351], regroupV0_hi_20[343]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_lo_15 = {regroupV0_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_20[367], regroupV0_hi_20[359]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_20[383], regroupV0_hi_20[375]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_hi_15 = {regroupV0_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_lo_hi_26 = {regroupV0_hi_hi_lo_hi_hi_15, regroupV0_hi_hi_lo_hi_lo_15};
  wire [15:0]       regroupV0_hi_hi_lo_26 = {regroupV0_hi_hi_lo_hi_26, regroupV0_hi_hi_lo_lo_26};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_20[399], regroupV0_hi_20[391]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_20[415], regroupV0_hi_20[407]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_lo_15 = {regroupV0_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_20[431], regroupV0_hi_20[423]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_20[447], regroupV0_hi_20[439]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_hi_15 = {regroupV0_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_hi_lo_26 = {regroupV0_hi_hi_hi_lo_hi_15, regroupV0_hi_hi_hi_lo_lo_15};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_20[463], regroupV0_hi_20[455]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_20[479], regroupV0_hi_20[471]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_lo_15 = {regroupV0_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_20[495], regroupV0_hi_20[487]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_20[511], regroupV0_hi_20[503]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_hi_15 = {regroupV0_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_hi_hi_26 = {regroupV0_hi_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_hi_lo_15};
  wire [15:0]       regroupV0_hi_hi_hi_26 = {regroupV0_hi_hi_hi_hi_26, regroupV0_hi_hi_hi_lo_26};
  wire [31:0]       regroupV0_hi_hi_28 = {regroupV0_hi_hi_hi_26, regroupV0_hi_hi_lo_26};
  wire [63:0]       regroupV0_hi_28 = {regroupV0_hi_hi_28, regroupV0_hi_lo_28};
  wire [255:0]      regroupV0_lo_lo_29 = {regroupV0_hi_22, regroupV0_lo_22, regroupV0_hi_21, regroupV0_lo_21};
  wire [255:0]      regroupV0_lo_hi_29 = {regroupV0_hi_24, regroupV0_lo_24, regroupV0_hi_23, regroupV0_lo_23};
  wire [511:0]      regroupV0_lo_29 = {regroupV0_lo_hi_29, regroupV0_lo_lo_29};
  wire [255:0]      regroupV0_hi_lo_29 = {regroupV0_hi_26, regroupV0_lo_26, regroupV0_hi_25, regroupV0_lo_25};
  wire [255:0]      regroupV0_hi_hi_29 = {regroupV0_hi_28, regroupV0_lo_28, regroupV0_hi_27, regroupV0_lo_27};
  wire [511:0]      regroupV0_hi_29 = {regroupV0_hi_hi_29, regroupV0_hi_lo_29};
  wire [1023:0]     regroupV0_2 = {regroupV0_hi_29, regroupV0_lo_29};
  wire [3:0]        _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [127:0]      v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[127:0] : 128'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[127:0] : 128'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[127:0] : 128'h0);
  wire [3:0][31:0]  _GEN_15 = {{v0SelectBySew[127:96]}, {v0SelectBySew[95:64]}, {v0SelectBySew[63:32]}, {v0SelectBySew[31:0]}};
  wire [3:0]        _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [127:0]      v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[255:128] : 128'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[255:128] : 128'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[255:128] : 128'h0);
  wire [3:0][31:0]  _GEN_16 = {{v0SelectBySew_1[127:96]}, {v0SelectBySew_1[95:64]}, {v0SelectBySew_1[63:32]}, {v0SelectBySew_1[31:0]}};
  wire [3:0]        _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [127:0]      v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[383:256] : 128'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[383:256] : 128'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[383:256] : 128'h0);
  wire [3:0][31:0]  _GEN_17 = {{v0SelectBySew_2[127:96]}, {v0SelectBySew_2[95:64]}, {v0SelectBySew_2[63:32]}, {v0SelectBySew_2[31:0]}};
  wire [3:0]        _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [127:0]      v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[511:384] : 128'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[511:384] : 128'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[511:384] : 128'h0);
  wire [3:0][31:0]  _GEN_18 = {{v0SelectBySew_3[127:96]}, {v0SelectBySew_3[95:64]}, {v0SelectBySew_3[63:32]}, {v0SelectBySew_3[31:0]}};
  wire [3:0]        _v0SelectBySew_T_36 = 4'h1 << laneMaskSewSelect_4;
  wire [127:0]      v0SelectBySew_4 = (_v0SelectBySew_T_36[0] ? regroupV0_0[639:512] : 128'h0) | (_v0SelectBySew_T_36[1] ? regroupV0_1[639:512] : 128'h0) | (_v0SelectBySew_T_36[2] ? regroupV0_2[639:512] : 128'h0);
  wire [3:0][31:0]  _GEN_19 = {{v0SelectBySew_4[127:96]}, {v0SelectBySew_4[95:64]}, {v0SelectBySew_4[63:32]}, {v0SelectBySew_4[31:0]}};
  wire [3:0]        _v0SelectBySew_T_45 = 4'h1 << laneMaskSewSelect_5;
  wire [127:0]      v0SelectBySew_5 = (_v0SelectBySew_T_45[0] ? regroupV0_0[767:640] : 128'h0) | (_v0SelectBySew_T_45[1] ? regroupV0_1[767:640] : 128'h0) | (_v0SelectBySew_T_45[2] ? regroupV0_2[767:640] : 128'h0);
  wire [3:0][31:0]  _GEN_20 = {{v0SelectBySew_5[127:96]}, {v0SelectBySew_5[95:64]}, {v0SelectBySew_5[63:32]}, {v0SelectBySew_5[31:0]}};
  wire [3:0]        _v0SelectBySew_T_54 = 4'h1 << laneMaskSewSelect_6;
  wire [127:0]      v0SelectBySew_6 = (_v0SelectBySew_T_54[0] ? regroupV0_0[895:768] : 128'h0) | (_v0SelectBySew_T_54[1] ? regroupV0_1[895:768] : 128'h0) | (_v0SelectBySew_T_54[2] ? regroupV0_2[895:768] : 128'h0);
  wire [3:0][31:0]  _GEN_21 = {{v0SelectBySew_6[127:96]}, {v0SelectBySew_6[95:64]}, {v0SelectBySew_6[63:32]}, {v0SelectBySew_6[31:0]}};
  wire [3:0]        _v0SelectBySew_T_63 = 4'h1 << laneMaskSewSelect_7;
  wire [127:0]      v0SelectBySew_7 = (_v0SelectBySew_T_63[0] ? regroupV0_0[1023:896] : 128'h0) | (_v0SelectBySew_T_63[1] ? regroupV0_1[1023:896] : 128'h0) | (_v0SelectBySew_T_63[2] ? regroupV0_2[1023:896] : 128'h0);
  wire [3:0][31:0]  _GEN_22 = {{v0SelectBySew_7[127:96]}, {v0SelectBySew_7[95:64]}, {v0SelectBySew_7[63:32]}, {v0SelectBySew_7[31:0]}};
  wire [3:0]        intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [12:0]       _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[9:0]} << instReq_bits_sew;
  wire [9:0]        dataPosition = _dataPosition_T_1[9:0];
  wire [3:0]        _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]        sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]        dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [2:0]        accessLane = dataPosition[4:2];
  wire [4:0]        dataGroup = dataPosition[9:5];
  wire [1:0]        offset = dataGroup[1:0];
  wire [2:0]        accessRegGrowth = dataGroup[4:2];
  wire [2:0]        reallyGrowth = accessRegGrowth;
  wire [4:0]        decimalProportion = {offset, accessLane};
  wire [2:0]        decimal = decimalProportion[4:2];
  wire              notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:10]};
  reg  [1:0]        gatherReadState;
  wire              gatherSRead = gatherReadState == 2'h1;
  wire              gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire              gatherData_valid_0 = gatherResponse;
  reg  [1:0]        gatherDatOffset;
  reg  [2:0]        gatherLane;
  reg  [1:0]        gatherOffset;
  reg  [2:0]        gatherGrowth;
  reg  [2:0]        instReg_instructionIndex;
  wire [2:0]        exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_4_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_5_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_6_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_7_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_3_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_4_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_5_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_6_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_7_enq_bits_index = instReg_instructionIndex;
  reg               instReg_decodeResult_orderReduce;
  reg               instReg_decodeResult_floatMul;
  reg  [1:0]        instReg_decodeResult_fpExecutionType;
  reg               instReg_decodeResult_float;
  reg               instReg_decodeResult_specialSlot;
  reg  [4:0]        instReg_decodeResult_topUop;
  reg               instReg_decodeResult_popCount;
  reg               instReg_decodeResult_ffo;
  reg               instReg_decodeResult_average;
  reg               instReg_decodeResult_reverse;
  reg               instReg_decodeResult_dontNeedExecuteInLane;
  reg               instReg_decodeResult_scheduler;
  reg               instReg_decodeResult_sReadVD;
  reg               instReg_decodeResult_vtype;
  reg               instReg_decodeResult_sWrite;
  reg               instReg_decodeResult_crossRead;
  reg               instReg_decodeResult_crossWrite;
  reg               instReg_decodeResult_maskUnit;
  reg               instReg_decodeResult_special;
  reg               instReg_decodeResult_saturate;
  reg               instReg_decodeResult_vwmacc;
  reg               instReg_decodeResult_readOnly;
  reg               instReg_decodeResult_maskSource;
  reg               instReg_decodeResult_maskDestination;
  reg               instReg_decodeResult_maskLogic;
  reg  [3:0]        instReg_decodeResult_uop;
  reg               instReg_decodeResult_iota;
  reg               instReg_decodeResult_mv;
  reg               instReg_decodeResult_extend;
  reg               instReg_decodeResult_unOrderWrite;
  reg               instReg_decodeResult_compress;
  reg               instReg_decodeResult_gather16;
  reg               instReg_decodeResult_gather;
  reg               instReg_decodeResult_slid;
  reg               instReg_decodeResult_targetRd;
  reg               instReg_decodeResult_widenReduce;
  reg               instReg_decodeResult_red;
  reg               instReg_decodeResult_nr;
  reg               instReg_decodeResult_itype;
  reg               instReg_decodeResult_unsigned1;
  reg               instReg_decodeResult_unsigned0;
  reg               instReg_decodeResult_other;
  reg               instReg_decodeResult_multiCycle;
  reg               instReg_decodeResult_divider;
  reg               instReg_decodeResult_multiplier;
  reg               instReg_decodeResult_shift;
  reg               instReg_decodeResult_adder;
  reg               instReg_decodeResult_logic;
  reg  [31:0]       instReg_readFromScala;
  reg  [1:0]        instReg_sew;
  reg  [2:0]        instReg_vlmul;
  reg               instReg_maskType;
  reg  [2:0]        instReg_vxrm;
  reg  [4:0]        instReg_vs2;
  reg  [4:0]        instReg_vs1;
  reg  [4:0]        instReg_vd;
  wire [4:0]        writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_3_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_4_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_5_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_6_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_7_writeData_vd = instReg_vd;
  reg  [10:0]       instReg_vl;
  wire [10:0]       reduceLastDataNeed_byteForVl = instReg_vl;
  wire              enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg               instVlValid;
  wire              gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire              viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg               readVS1Reg_dataValid;
  reg               readVS1Reg_requestSend;
  reg               readVS1Reg_sendToExecution;
  reg  [31:0]       readVS1Reg_data;
  reg  [4:0]        readVS1Reg_readIndex;
  wire [3:0]        _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]        sew1H = _sew1H_T[2:0];
  wire [3:0]        unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]        subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire              readType = unitType[0];
  wire              gather16 = instReg_decodeResult_topUop == 5'h5;
  wire              maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire              compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire              viota = instReg_decodeResult_topUop == 5'h8;
  wire              mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire              mvRd = instReg_decodeResult_topUop == 5'hB;
  wire              mvVd = instReg_decodeResult_topUop == 5'hA;
  wire              orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire              ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire              extendType = unitType[3] & (subType[2] | subType[1]);
  wire              readValid = readType & instVlValid;
  wire              noSource = mv | viota;
  wire              allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire              useDefaultSew = readType & ~gather16;
  wire [1:0]        _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]        dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire              sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]        _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]        sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]        executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]        lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]        _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]        sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [9:0]        lastElementIndex = instReg_vl[9:0] - {9'h0, |instReg_vl};
  wire [9:0]        processingVl_lastByteIndex = lastElementIndex;
  wire              maskFormatSource = ffo | maskDestinationType;
  wire [4:0]        processingVl_lastGroupRemaining = processingVl_lastByteIndex[4:0];
  wire [4:0]        processingVl_0_1 = processingVl_lastByteIndex[9:5];
  wire [2:0]        processingVl_lastLaneIndex = processingVl_lastGroupRemaining[4:2];
  wire [7:0]        _processingVl_lastGroupDataNeed_T = 8'h1 << processingVl_lastLaneIndex;
  wire [6:0]        _GEN_23 = _processingVl_lastGroupDataNeed_T[6:0] | _processingVl_lastGroupDataNeed_T[7:1];
  wire [5:0]        _GEN_24 = _GEN_23[5:0] | {_processingVl_lastGroupDataNeed_T[7], _GEN_23[6:2]};
  wire [7:0]        processingVl_0_2 = {_processingVl_lastGroupDataNeed_T[7], _GEN_23[6], _GEN_24[5:4], _GEN_24[3:0] | {_processingVl_lastGroupDataNeed_T[7], _GEN_23[6], _GEN_24[5:4]}};
  wire [10:0]       processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [4:0]        processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[4:0];
  wire [5:0]        processingVl_1_1 = processingVl_lastByteIndex_1[10:5];
  wire [2:0]        processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[4:2];
  wire [7:0]        _processingVl_lastGroupDataNeed_T_7 = 8'h1 << processingVl_lastLaneIndex_1;
  wire [6:0]        _GEN_25 = _processingVl_lastGroupDataNeed_T_7[6:0] | _processingVl_lastGroupDataNeed_T_7[7:1];
  wire [5:0]        _GEN_26 = _GEN_25[5:0] | {_processingVl_lastGroupDataNeed_T_7[7], _GEN_25[6:2]};
  wire [7:0]        processingVl_1_2 = {_processingVl_lastGroupDataNeed_T_7[7], _GEN_25[6], _GEN_26[5:4], _GEN_26[3:0] | {_processingVl_lastGroupDataNeed_T_7[7], _GEN_25[6], _GEN_26[5:4]}};
  wire [11:0]       processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [4:0]        processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[4:0];
  wire [6:0]        processingVl_2_1 = processingVl_lastByteIndex_2[11:5];
  wire [2:0]        processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[4:2];
  wire [7:0]        _processingVl_lastGroupDataNeed_T_14 = 8'h1 << processingVl_lastLaneIndex_2;
  wire [6:0]        _GEN_27 = _processingVl_lastGroupDataNeed_T_14[6:0] | _processingVl_lastGroupDataNeed_T_14[7:1];
  wire [5:0]        _GEN_28 = _GEN_27[5:0] | {_processingVl_lastGroupDataNeed_T_14[7], _GEN_27[6:2]};
  wire [7:0]        processingVl_2_2 = {_processingVl_lastGroupDataNeed_T_14[7], _GEN_27[6], _GEN_28[5:4], _GEN_28[3:0] | {_processingVl_lastGroupDataNeed_T_14[7], _GEN_27[6], _GEN_28[5:4]}};
  wire [7:0]        processingMaskVl_lastGroupRemaining = lastElementIndex[7:0];
  wire [7:0]        elementTailForMaskDestination = lastElementIndex[7:0];
  wire              processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire [1:0]        processingMaskVl_0_1 = lastElementIndex[9:8];
  wire [2:0]        processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[7:5] - {2'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [7:0]        _processingMaskVl_dataNeedForPL_T = 8'h1 << processingMaskVl_lastLaneIndex;
  wire [6:0]        _GEN_29 = _processingMaskVl_dataNeedForPL_T[6:0] | _processingMaskVl_dataNeedForPL_T[7:1];
  wire [5:0]        _GEN_30 = _GEN_29[5:0] | {_processingMaskVl_dataNeedForPL_T[7], _GEN_29[6:2]};
  wire [7:0]        processingMaskVl_dataNeedForPL = {_processingMaskVl_dataNeedForPL_T[7], _GEN_29[6], _GEN_30[5:4], _GEN_30[3:0] | {_processingMaskVl_dataNeedForPL_T[7], _GEN_29[6], _GEN_30[5:4]}};
  wire              processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [6:0]        processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[7:2]} + {6'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire              processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[6:3]);
  wire [2:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[2:0];
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T = 8'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[6:0], 1'h0};
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_6 = _processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[5:0], 2'h0};
  wire [7:0]        processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_6 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_6[3:0], 4'h0}) | {8{processingMaskVl_dataNeedForNPL_allNeed}};
  wire              processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [7:0]        processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[7:1]} + {7'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire              processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[7:3]);
  wire [2:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[2:0];
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_13 = 8'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_16 = _processingMaskVl_dataNeedForNPL_dataNeed_T_13 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_13[6:0], 1'h0};
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_19 = _processingMaskVl_dataNeedForNPL_dataNeed_T_16 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_16[5:0], 2'h0};
  wire [7:0]        processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_19 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_19[3:0], 4'h0}) | {8{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [8:0]        processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire              processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[8:3]);
  wire [2:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[2:0];
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_26 = 8'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_29 = _processingMaskVl_dataNeedForNPL_dataNeed_T_26 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_26[6:0], 1'h0};
  wire [7:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_32 = _processingMaskVl_dataNeedForNPL_dataNeed_T_29 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_29[5:0], 2'h0};
  wire [7:0]        processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_32 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_32[3:0], 4'h0}) | {8{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [7:0]        processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 8'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 8'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 8'h0);
  wire [7:0]        processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire              reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[10:5]);
  wire [4:0]        reduceLastDataNeed_vlLSB = instReg_vl[4:0];
  wire [4:0]        reduceLastDataNeed_vlLSB_1 = instReg_vl[4:0];
  wire [4:0]        reduceLastDataNeed_vlLSB_2 = instReg_vl[4:0];
  wire [2:0]        reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[4:2] - {2'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [7:0]        _reduceLastDataNeed_T = 8'h1 << reduceLastDataNeed_lsbDSize;
  wire [6:0]        _GEN_31 = _reduceLastDataNeed_T[6:0] | _reduceLastDataNeed_T[7:1];
  wire [5:0]        _GEN_32 = _GEN_31[5:0] | {_reduceLastDataNeed_T[7], _GEN_31[6:2]};
  wire [11:0]       reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire              reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[11:5]);
  wire [2:0]        reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[4:2] - {2'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [7:0]        _reduceLastDataNeed_T_10 = 8'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [6:0]        _GEN_33 = _reduceLastDataNeed_T_10[6:0] | _reduceLastDataNeed_T_10[7:1];
  wire [5:0]        _GEN_34 = _GEN_33[5:0] | {_reduceLastDataNeed_T_10[7], _GEN_33[6:2]};
  wire [12:0]       reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire              reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[12:5]);
  wire [2:0]        reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[4:2] - {2'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [7:0]        _reduceLastDataNeed_T_20 = 8'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [6:0]        _GEN_35 = _reduceLastDataNeed_T_20[6:0] | _reduceLastDataNeed_T_20[7:1];
  wire [5:0]        _GEN_36 = _GEN_35[5:0] | {_reduceLastDataNeed_T_20[7], _GEN_35[6:2]};
  wire [7:0]        reduceLastDataNeed =
    (sew1H[0] ? {_reduceLastDataNeed_T[7], _GEN_31[6], _GEN_32[5:4], _GEN_32[3:0] | {_reduceLastDataNeed_T[7], _GEN_31[6], _GEN_32[5:4]}} | {8{reduceLastDataNeed_vlMSB}} : 8'h0)
    | (sew1H[1] ? {_reduceLastDataNeed_T_10[7], _GEN_33[6], _GEN_34[5:4], _GEN_34[3:0] | {_reduceLastDataNeed_T_10[7], _GEN_33[6], _GEN_34[5:4]}} | {8{reduceLastDataNeed_vlMSB_1}} : 8'h0)
    | (sew1H[2] ? {_reduceLastDataNeed_T_20[7], _GEN_35[6], _GEN_36[5:4], _GEN_36[3:0] | {_reduceLastDataNeed_T_20[7], _GEN_35[6], _GEN_36[5:4]}} | {8{reduceLastDataNeed_vlMSB_2}} : 8'h0);
  wire [1:0]        dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]        _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]        dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire              unorderReduce = ~orderReduce & unitType[2];
  wire              normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [6:0]        lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource ? processingMaskVl_0_1 : 2'h0} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 5'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 6'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 7'h0);
  wire [4:0]        popDataNeed_dataPathGroups = lastElementIndex[9:5];
  wire [2:0]        popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[2:0];
  wire              popDataNeed_lagerThanDLen = |(popDataNeed_dataPathGroups[4:3]);
  wire [7:0]        _popDataNeed_T = 8'h1 << popDataNeed_lastLaneIndex;
  wire [6:0]        _GEN_37 = _popDataNeed_T[6:0] | _popDataNeed_T[7:1];
  wire [5:0]        _GEN_38 = _GEN_37[5:0] | {_popDataNeed_T[7], _GEN_37[6:2]};
  wire [7:0]        popDataNeed = {_popDataNeed_T[7], _GEN_37[6], _GEN_38[5:4], _GEN_38[3:0] | {_popDataNeed_T[7], _GEN_37[6], _GEN_38[5:4]}} | {8{popDataNeed_lagerThanDLen}};
  wire [7:0]        lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 8'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 8'h0) | (maskFormatSource ? processingMaskVl_0_2 : 8'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 8'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 8'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 8'h0);
  wire [1:0]        exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_ffo, exeRequestQueue_0_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_queue_dataIn_hi_hi, exeRequestQueue_0_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire              exeRequestQueue_queue_dataOut_fpReduceValid = _exeRequestQueue_queue_fifo_data_out[0];
  wire              exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[68:37];
  wire              exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_0_deq_ready;
  wire              exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]       exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]       exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]        exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire              exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire              exeRequestQueue_0_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_fpReduceValid;
  wire              tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_ffo, exeRequestQueue_1_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_queue_dataIn_hi_hi_1, exeRequestQueue_1_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire              exeRequestQueue_queue_dataOut_1_fpReduceValid = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire              exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[68:37];
  wire              exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_1_deq_ready;
  wire              exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]       exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]       exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]        exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire              exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire              exeRequestQueue_1_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_1_fpReduceValid;
  wire              tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_ffo, exeRequestQueue_2_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_queue_dataIn_hi_hi_2, exeRequestQueue_2_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire              exeRequestQueue_queue_dataOut_2_fpReduceValid = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire              exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[68:37];
  wire              exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_2_deq_ready;
  wire              exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]       exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]       exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]        exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire              exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire              exeRequestQueue_2_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_2_fpReduceValid;
  wire              tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_ffo, exeRequestQueue_3_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_queue_dataIn_hi_hi_3, exeRequestQueue_3_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire              exeRequestQueue_queue_dataOut_3_fpReduceValid = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire              exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[68:37];
  wire              exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire              exeRequestQueue_3_deq_ready;
  wire              exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]       exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]       exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]        exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire              exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire              exeRequestQueue_3_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_3_fpReduceValid;
  wire              tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_4 = {exeRequestQueue_4_enq_bits_ffo, exeRequestQueue_4_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_4 = {exeRequestQueue_4_enq_bits_source1, exeRequestQueue_4_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_4 = {exeRequestQueue_queue_dataIn_hi_hi_4, exeRequestQueue_4_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_4 = {exeRequestQueue_queue_dataIn_hi_4, exeRequestQueue_queue_dataIn_lo_4};
  wire              exeRequestQueue_queue_dataOut_4_fpReduceValid = _exeRequestQueue_queue_fifo_4_data_out[0];
  wire              exeRequestQueue_queue_dataOut_4_ffo = _exeRequestQueue_queue_fifo_4_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_4_index = _exeRequestQueue_queue_fifo_4_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_4_source2 = _exeRequestQueue_queue_fifo_4_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_4_source1 = _exeRequestQueue_queue_fifo_4_data_out[68:37];
  wire              exeRequestQueue_4_enq_ready = ~_exeRequestQueue_queue_fifo_4_full;
  wire              exeRequestQueue_4_deq_ready;
  wire              exeRequestQueue_4_deq_valid = ~_exeRequestQueue_queue_fifo_4_empty | exeRequestQueue_4_enq_valid;
  wire [31:0]       exeRequestQueue_4_deq_bits_source1 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source1 : exeRequestQueue_queue_dataOut_4_source1;
  wire [31:0]       exeRequestQueue_4_deq_bits_source2 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source2 : exeRequestQueue_queue_dataOut_4_source2;
  wire [2:0]        exeRequestQueue_4_deq_bits_index = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_index : exeRequestQueue_queue_dataOut_4_index;
  wire              exeRequestQueue_4_deq_bits_ffo = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_ffo : exeRequestQueue_queue_dataOut_4_ffo;
  wire              exeRequestQueue_4_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_4_fpReduceValid;
  wire              tokenIO_4_maskRequestRelease_0 = exeRequestQueue_4_deq_ready & exeRequestQueue_4_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_5 = {exeRequestQueue_5_enq_bits_ffo, exeRequestQueue_5_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_5 = {exeRequestQueue_5_enq_bits_source1, exeRequestQueue_5_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_5 = {exeRequestQueue_queue_dataIn_hi_hi_5, exeRequestQueue_5_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_5 = {exeRequestQueue_queue_dataIn_hi_5, exeRequestQueue_queue_dataIn_lo_5};
  wire              exeRequestQueue_queue_dataOut_5_fpReduceValid = _exeRequestQueue_queue_fifo_5_data_out[0];
  wire              exeRequestQueue_queue_dataOut_5_ffo = _exeRequestQueue_queue_fifo_5_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_5_index = _exeRequestQueue_queue_fifo_5_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_5_source2 = _exeRequestQueue_queue_fifo_5_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_5_source1 = _exeRequestQueue_queue_fifo_5_data_out[68:37];
  wire              exeRequestQueue_5_enq_ready = ~_exeRequestQueue_queue_fifo_5_full;
  wire              exeRequestQueue_5_deq_ready;
  wire              exeRequestQueue_5_deq_valid = ~_exeRequestQueue_queue_fifo_5_empty | exeRequestQueue_5_enq_valid;
  wire [31:0]       exeRequestQueue_5_deq_bits_source1 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source1 : exeRequestQueue_queue_dataOut_5_source1;
  wire [31:0]       exeRequestQueue_5_deq_bits_source2 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source2 : exeRequestQueue_queue_dataOut_5_source2;
  wire [2:0]        exeRequestQueue_5_deq_bits_index = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_index : exeRequestQueue_queue_dataOut_5_index;
  wire              exeRequestQueue_5_deq_bits_ffo = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_ffo : exeRequestQueue_queue_dataOut_5_ffo;
  wire              exeRequestQueue_5_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_5_fpReduceValid;
  wire              tokenIO_5_maskRequestRelease_0 = exeRequestQueue_5_deq_ready & exeRequestQueue_5_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_6 = {exeRequestQueue_6_enq_bits_ffo, exeRequestQueue_6_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_6 = {exeRequestQueue_6_enq_bits_source1, exeRequestQueue_6_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_6 = {exeRequestQueue_queue_dataIn_hi_hi_6, exeRequestQueue_6_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_6 = {exeRequestQueue_queue_dataIn_hi_6, exeRequestQueue_queue_dataIn_lo_6};
  wire              exeRequestQueue_queue_dataOut_6_fpReduceValid = _exeRequestQueue_queue_fifo_6_data_out[0];
  wire              exeRequestQueue_queue_dataOut_6_ffo = _exeRequestQueue_queue_fifo_6_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_6_index = _exeRequestQueue_queue_fifo_6_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_6_source2 = _exeRequestQueue_queue_fifo_6_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_6_source1 = _exeRequestQueue_queue_fifo_6_data_out[68:37];
  wire              exeRequestQueue_6_enq_ready = ~_exeRequestQueue_queue_fifo_6_full;
  wire              exeRequestQueue_6_deq_ready;
  wire              exeRequestQueue_6_deq_valid = ~_exeRequestQueue_queue_fifo_6_empty | exeRequestQueue_6_enq_valid;
  wire [31:0]       exeRequestQueue_6_deq_bits_source1 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source1 : exeRequestQueue_queue_dataOut_6_source1;
  wire [31:0]       exeRequestQueue_6_deq_bits_source2 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source2 : exeRequestQueue_queue_dataOut_6_source2;
  wire [2:0]        exeRequestQueue_6_deq_bits_index = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_index : exeRequestQueue_queue_dataOut_6_index;
  wire              exeRequestQueue_6_deq_bits_ffo = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_ffo : exeRequestQueue_queue_dataOut_6_ffo;
  wire              exeRequestQueue_6_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_6_fpReduceValid;
  wire              tokenIO_6_maskRequestRelease_0 = exeRequestQueue_6_deq_ready & exeRequestQueue_6_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_7 = {exeRequestQueue_7_enq_bits_ffo, exeRequestQueue_7_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_7 = {exeRequestQueue_7_enq_bits_source1, exeRequestQueue_7_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_7 = {exeRequestQueue_queue_dataIn_hi_hi_7, exeRequestQueue_7_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_7 = {exeRequestQueue_queue_dataIn_hi_7, exeRequestQueue_queue_dataIn_lo_7};
  wire              exeRequestQueue_queue_dataOut_7_fpReduceValid = _exeRequestQueue_queue_fifo_7_data_out[0];
  wire              exeRequestQueue_queue_dataOut_7_ffo = _exeRequestQueue_queue_fifo_7_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_7_index = _exeRequestQueue_queue_fifo_7_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_7_source2 = _exeRequestQueue_queue_fifo_7_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_7_source1 = _exeRequestQueue_queue_fifo_7_data_out[68:37];
  wire              exeRequestQueue_7_enq_ready = ~_exeRequestQueue_queue_fifo_7_full;
  wire              exeRequestQueue_7_deq_ready;
  wire              exeRequestQueue_7_deq_valid = ~_exeRequestQueue_queue_fifo_7_empty | exeRequestQueue_7_enq_valid;
  wire [31:0]       exeRequestQueue_7_deq_bits_source1 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source1 : exeRequestQueue_queue_dataOut_7_source1;
  wire [31:0]       exeRequestQueue_7_deq_bits_source2 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source2 : exeRequestQueue_queue_dataOut_7_source2;
  wire [2:0]        exeRequestQueue_7_deq_bits_index = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_index : exeRequestQueue_queue_dataOut_7_index;
  wire              exeRequestQueue_7_deq_bits_ffo = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_ffo : exeRequestQueue_queue_dataOut_7_ffo;
  wire              exeRequestQueue_7_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_7_fpReduceValid;
  wire              tokenIO_7_maskRequestRelease_0 = exeRequestQueue_7_deq_ready & exeRequestQueue_7_deq_valid;
  reg               exeReqReg_0_valid;
  reg  [31:0]       exeReqReg_0_bits_source1;
  reg  [31:0]       exeReqReg_0_bits_source2;
  reg  [2:0]        exeReqReg_0_bits_index;
  reg               exeReqReg_0_bits_ffo;
  reg               exeReqReg_0_bits_fpReduceValid;
  reg               exeReqReg_1_valid;
  reg  [31:0]       exeReqReg_1_bits_source1;
  reg  [31:0]       exeReqReg_1_bits_source2;
  reg  [2:0]        exeReqReg_1_bits_index;
  reg               exeReqReg_1_bits_ffo;
  reg               exeReqReg_1_bits_fpReduceValid;
  reg               exeReqReg_2_valid;
  reg  [31:0]       exeReqReg_2_bits_source1;
  reg  [31:0]       exeReqReg_2_bits_source2;
  reg  [2:0]        exeReqReg_2_bits_index;
  reg               exeReqReg_2_bits_ffo;
  reg               exeReqReg_2_bits_fpReduceValid;
  reg               exeReqReg_3_valid;
  reg  [31:0]       exeReqReg_3_bits_source1;
  reg  [31:0]       exeReqReg_3_bits_source2;
  reg  [2:0]        exeReqReg_3_bits_index;
  reg               exeReqReg_3_bits_ffo;
  reg               exeReqReg_3_bits_fpReduceValid;
  reg               exeReqReg_4_valid;
  reg  [31:0]       exeReqReg_4_bits_source1;
  reg  [31:0]       exeReqReg_4_bits_source2;
  reg  [2:0]        exeReqReg_4_bits_index;
  reg               exeReqReg_4_bits_ffo;
  reg               exeReqReg_4_bits_fpReduceValid;
  reg               exeReqReg_5_valid;
  reg  [31:0]       exeReqReg_5_bits_source1;
  reg  [31:0]       exeReqReg_5_bits_source2;
  reg  [2:0]        exeReqReg_5_bits_index;
  reg               exeReqReg_5_bits_ffo;
  reg               exeReqReg_5_bits_fpReduceValid;
  reg               exeReqReg_6_valid;
  reg  [31:0]       exeReqReg_6_bits_source1;
  reg  [31:0]       exeReqReg_6_bits_source2;
  reg  [2:0]        exeReqReg_6_bits_index;
  reg               exeReqReg_6_bits_ffo;
  reg               exeReqReg_6_bits_fpReduceValid;
  reg               exeReqReg_7_valid;
  reg  [31:0]       exeReqReg_7_bits_source1;
  reg  [31:0]       exeReqReg_7_bits_source2;
  reg  [2:0]        exeReqReg_7_bits_index;
  reg               exeReqReg_7_bits_ffo;
  reg               exeReqReg_7_bits_fpReduceValid;
  reg  [5:0]        requestCounter;
  wire [6:0]        _GEN_39 = {1'h0, requestCounter};
  wire              counterValid = _GEN_39 <= lastGroupForInstruction;
  wire              lastGroup = _GEN_39 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]      slideAddressGen_slideMaskInput_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo};
  wire [511:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo};
  wire [511:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [127:0][7:0] _GEN_40 =
    {{slideAddressGen_slideMaskInput_hi[511:504]},
     {slideAddressGen_slideMaskInput_hi[503:496]},
     {slideAddressGen_slideMaskInput_hi[495:488]},
     {slideAddressGen_slideMaskInput_hi[487:480]},
     {slideAddressGen_slideMaskInput_hi[479:472]},
     {slideAddressGen_slideMaskInput_hi[471:464]},
     {slideAddressGen_slideMaskInput_hi[463:456]},
     {slideAddressGen_slideMaskInput_hi[455:448]},
     {slideAddressGen_slideMaskInput_hi[447:440]},
     {slideAddressGen_slideMaskInput_hi[439:432]},
     {slideAddressGen_slideMaskInput_hi[431:424]},
     {slideAddressGen_slideMaskInput_hi[423:416]},
     {slideAddressGen_slideMaskInput_hi[415:408]},
     {slideAddressGen_slideMaskInput_hi[407:400]},
     {slideAddressGen_slideMaskInput_hi[399:392]},
     {slideAddressGen_slideMaskInput_hi[391:384]},
     {slideAddressGen_slideMaskInput_hi[383:376]},
     {slideAddressGen_slideMaskInput_hi[375:368]},
     {slideAddressGen_slideMaskInput_hi[367:360]},
     {slideAddressGen_slideMaskInput_hi[359:352]},
     {slideAddressGen_slideMaskInput_hi[351:344]},
     {slideAddressGen_slideMaskInput_hi[343:336]},
     {slideAddressGen_slideMaskInput_hi[335:328]},
     {slideAddressGen_slideMaskInput_hi[327:320]},
     {slideAddressGen_slideMaskInput_hi[319:312]},
     {slideAddressGen_slideMaskInput_hi[311:304]},
     {slideAddressGen_slideMaskInput_hi[303:296]},
     {slideAddressGen_slideMaskInput_hi[295:288]},
     {slideAddressGen_slideMaskInput_hi[287:280]},
     {slideAddressGen_slideMaskInput_hi[279:272]},
     {slideAddressGen_slideMaskInput_hi[271:264]},
     {slideAddressGen_slideMaskInput_hi[263:256]},
     {slideAddressGen_slideMaskInput_hi[255:248]},
     {slideAddressGen_slideMaskInput_hi[247:240]},
     {slideAddressGen_slideMaskInput_hi[239:232]},
     {slideAddressGen_slideMaskInput_hi[231:224]},
     {slideAddressGen_slideMaskInput_hi[223:216]},
     {slideAddressGen_slideMaskInput_hi[215:208]},
     {slideAddressGen_slideMaskInput_hi[207:200]},
     {slideAddressGen_slideMaskInput_hi[199:192]},
     {slideAddressGen_slideMaskInput_hi[191:184]},
     {slideAddressGen_slideMaskInput_hi[183:176]},
     {slideAddressGen_slideMaskInput_hi[175:168]},
     {slideAddressGen_slideMaskInput_hi[167:160]},
     {slideAddressGen_slideMaskInput_hi[159:152]},
     {slideAddressGen_slideMaskInput_hi[151:144]},
     {slideAddressGen_slideMaskInput_hi[143:136]},
     {slideAddressGen_slideMaskInput_hi[135:128]},
     {slideAddressGen_slideMaskInput_hi[127:120]},
     {slideAddressGen_slideMaskInput_hi[119:112]},
     {slideAddressGen_slideMaskInput_hi[111:104]},
     {slideAddressGen_slideMaskInput_hi[103:96]},
     {slideAddressGen_slideMaskInput_hi[95:88]},
     {slideAddressGen_slideMaskInput_hi[87:80]},
     {slideAddressGen_slideMaskInput_hi[79:72]},
     {slideAddressGen_slideMaskInput_hi[71:64]},
     {slideAddressGen_slideMaskInput_hi[63:56]},
     {slideAddressGen_slideMaskInput_hi[55:48]},
     {slideAddressGen_slideMaskInput_hi[47:40]},
     {slideAddressGen_slideMaskInput_hi[39:32]},
     {slideAddressGen_slideMaskInput_hi[31:24]},
     {slideAddressGen_slideMaskInput_hi[23:16]},
     {slideAddressGen_slideMaskInput_hi[15:8]},
     {slideAddressGen_slideMaskInput_hi[7:0]},
     {slideAddressGen_slideMaskInput_lo[511:504]},
     {slideAddressGen_slideMaskInput_lo[503:496]},
     {slideAddressGen_slideMaskInput_lo[495:488]},
     {slideAddressGen_slideMaskInput_lo[487:480]},
     {slideAddressGen_slideMaskInput_lo[479:472]},
     {slideAddressGen_slideMaskInput_lo[471:464]},
     {slideAddressGen_slideMaskInput_lo[463:456]},
     {slideAddressGen_slideMaskInput_lo[455:448]},
     {slideAddressGen_slideMaskInput_lo[447:440]},
     {slideAddressGen_slideMaskInput_lo[439:432]},
     {slideAddressGen_slideMaskInput_lo[431:424]},
     {slideAddressGen_slideMaskInput_lo[423:416]},
     {slideAddressGen_slideMaskInput_lo[415:408]},
     {slideAddressGen_slideMaskInput_lo[407:400]},
     {slideAddressGen_slideMaskInput_lo[399:392]},
     {slideAddressGen_slideMaskInput_lo[391:384]},
     {slideAddressGen_slideMaskInput_lo[383:376]},
     {slideAddressGen_slideMaskInput_lo[375:368]},
     {slideAddressGen_slideMaskInput_lo[367:360]},
     {slideAddressGen_slideMaskInput_lo[359:352]},
     {slideAddressGen_slideMaskInput_lo[351:344]},
     {slideAddressGen_slideMaskInput_lo[343:336]},
     {slideAddressGen_slideMaskInput_lo[335:328]},
     {slideAddressGen_slideMaskInput_lo[327:320]},
     {slideAddressGen_slideMaskInput_lo[319:312]},
     {slideAddressGen_slideMaskInput_lo[311:304]},
     {slideAddressGen_slideMaskInput_lo[303:296]},
     {slideAddressGen_slideMaskInput_lo[295:288]},
     {slideAddressGen_slideMaskInput_lo[287:280]},
     {slideAddressGen_slideMaskInput_lo[279:272]},
     {slideAddressGen_slideMaskInput_lo[271:264]},
     {slideAddressGen_slideMaskInput_lo[263:256]},
     {slideAddressGen_slideMaskInput_lo[255:248]},
     {slideAddressGen_slideMaskInput_lo[247:240]},
     {slideAddressGen_slideMaskInput_lo[239:232]},
     {slideAddressGen_slideMaskInput_lo[231:224]},
     {slideAddressGen_slideMaskInput_lo[223:216]},
     {slideAddressGen_slideMaskInput_lo[215:208]},
     {slideAddressGen_slideMaskInput_lo[207:200]},
     {slideAddressGen_slideMaskInput_lo[199:192]},
     {slideAddressGen_slideMaskInput_lo[191:184]},
     {slideAddressGen_slideMaskInput_lo[183:176]},
     {slideAddressGen_slideMaskInput_lo[175:168]},
     {slideAddressGen_slideMaskInput_lo[167:160]},
     {slideAddressGen_slideMaskInput_lo[159:152]},
     {slideAddressGen_slideMaskInput_lo[151:144]},
     {slideAddressGen_slideMaskInput_lo[143:136]},
     {slideAddressGen_slideMaskInput_lo[135:128]},
     {slideAddressGen_slideMaskInput_lo[127:120]},
     {slideAddressGen_slideMaskInput_lo[119:112]},
     {slideAddressGen_slideMaskInput_lo[111:104]},
     {slideAddressGen_slideMaskInput_lo[103:96]},
     {slideAddressGen_slideMaskInput_lo[95:88]},
     {slideAddressGen_slideMaskInput_lo[87:80]},
     {slideAddressGen_slideMaskInput_lo[79:72]},
     {slideAddressGen_slideMaskInput_lo[71:64]},
     {slideAddressGen_slideMaskInput_lo[63:56]},
     {slideAddressGen_slideMaskInput_lo[55:48]},
     {slideAddressGen_slideMaskInput_lo[47:40]},
     {slideAddressGen_slideMaskInput_lo[39:32]},
     {slideAddressGen_slideMaskInput_lo[31:24]},
     {slideAddressGen_slideMaskInput_lo[23:16]},
     {slideAddressGen_slideMaskInput_lo[15:8]},
     {slideAddressGen_slideMaskInput_lo[7:0]}};
  wire              lastExecuteGroupDeq;
  wire              viotaCounterAdd;
  wire              groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [7:0]        groupDataNeed = lastGroup ? lastGroupDataNeed : 8'hFF;
  reg  [1:0]        executeIndex;
  reg  [7:0]        readIssueStageState_groupReadState;
  reg  [7:0]        readIssueStageState_needRead;
  wire [7:0]        readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [7:0]        readIssueStageState_elementValid;
  wire [7:0]        readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [7:0]        readIssueStageState_replaceVs1;
  wire [7:0]        readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [15:0]       readIssueStageState_readOffset;
  reg  [2:0]        readIssueStageState_accessLane_0;
  reg  [2:0]        readIssueStageState_accessLane_1;
  wire [2:0]        selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [2:0]        readIssueStageState_accessLane_2;
  wire [2:0]        selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [2:0]        readIssueStageState_accessLane_3;
  wire [2:0]        selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [2:0]        readIssueStageState_accessLane_4;
  wire [2:0]        selectExecuteReq_4_bits_readLane = readIssueStageState_accessLane_4;
  reg  [2:0]        readIssueStageState_accessLane_5;
  wire [2:0]        selectExecuteReq_5_bits_readLane = readIssueStageState_accessLane_5;
  reg  [2:0]        readIssueStageState_accessLane_6;
  wire [2:0]        selectExecuteReq_6_bits_readLane = readIssueStageState_accessLane_6;
  reg  [2:0]        readIssueStageState_accessLane_7;
  wire [2:0]        selectExecuteReq_7_bits_readLane = readIssueStageState_accessLane_7;
  reg  [2:0]        readIssueStageState_vsGrowth_0;
  reg  [2:0]        readIssueStageState_vsGrowth_1;
  reg  [2:0]        readIssueStageState_vsGrowth_2;
  reg  [2:0]        readIssueStageState_vsGrowth_3;
  reg  [2:0]        readIssueStageState_vsGrowth_4;
  reg  [2:0]        readIssueStageState_vsGrowth_5;
  reg  [2:0]        readIssueStageState_vsGrowth_6;
  reg  [2:0]        readIssueStageState_vsGrowth_7;
  reg  [7:0]        readIssueStageState_executeGroup;
  wire [7:0]        readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [15:0]       readIssueStageState_readDataOffset;
  reg               readIssueStageState_last;
  wire              readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg               readIssueStageValid;
  wire [3:0]        accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [3:0]        accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [3:0]        accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [3:0]        accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire [3:0]        accessCountQueue_enq_bits_4 = accessCountEnq_4;
  wire [3:0]        accessCountQueue_enq_bits_5 = accessCountEnq_5;
  wire [3:0]        accessCountQueue_enq_bits_6 = accessCountEnq_6;
  wire [3:0]        accessCountQueue_enq_bits_7 = accessCountEnq_7;
  wire              readIssueStageEnq;
  wire              accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [3:0]        accessCountQueue_dataOut_0;
  wire [3:0]        accessCountQueue_dataOut_1;
  wire [3:0]        accessCountQueue_dataOut_2;
  wire [3:0]        accessCountQueue_dataOut_3;
  wire [3:0]        accessCountQueue_dataOut_4;
  wire [3:0]        accessCountQueue_dataOut_5;
  wire [3:0]        accessCountQueue_dataOut_6;
  wire [3:0]        accessCountQueue_dataOut_7;
  wire [7:0]        accessCountQueue_dataIn_lo_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [7:0]        accessCountQueue_dataIn_lo_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [15:0]       accessCountQueue_dataIn_lo = {accessCountQueue_dataIn_lo_hi, accessCountQueue_dataIn_lo_lo};
  wire [7:0]        accessCountQueue_dataIn_hi_lo = {accessCountQueue_enq_bits_5, accessCountQueue_enq_bits_4};
  wire [7:0]        accessCountQueue_dataIn_hi_hi = {accessCountQueue_enq_bits_7, accessCountQueue_enq_bits_6};
  wire [15:0]       accessCountQueue_dataIn_hi = {accessCountQueue_dataIn_hi_hi, accessCountQueue_dataIn_hi_lo};
  wire [31:0]       accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[3:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[7:4];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[11:8];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[15:12];
  assign accessCountQueue_dataOut_4 = _accessCountQueue_fifo_data_out[19:16];
  assign accessCountQueue_dataOut_5 = _accessCountQueue_fifo_data_out[23:20];
  assign accessCountQueue_dataOut_6 = _accessCountQueue_fifo_data_out[27:24];
  assign accessCountQueue_dataOut_7 = _accessCountQueue_fifo_data_out[31:28];
  wire [3:0]        accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [3:0]        accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [3:0]        accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [3:0]        accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire [3:0]        accessCountQueue_deq_bits_4 = accessCountQueue_dataOut_4;
  wire [3:0]        accessCountQueue_deq_bits_5 = accessCountQueue_dataOut_5;
  wire [3:0]        accessCountQueue_deq_bits_6 = accessCountQueue_dataOut_6;
  wire [3:0]        accessCountQueue_deq_bits_7 = accessCountQueue_dataOut_7;
  wire              accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire              accessCountQueue_enq_valid;
  wire              accessCountQueue_deq_ready;
  wire [7:0]        _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [7:0]        _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 8'h0;
  wire [6:0]        _GEN_41 = _executeGroup_T_8[6:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 7'h0);
  wire [7:0]        executeGroup = {_executeGroup_T_8[7], _GEN_41[6], _GEN_41[5:0] | (executeIndexGrowth[2] ? requestCounter : 6'h0)};
  wire              vlMisAlign;
  assign vlMisAlign = |(instReg_vl[2:0]);
  wire [7:0]        lastexecuteGroup = instReg_vl[10:3] - {7'h0, ~vlMisAlign};
  wire              isVlBoundary = executeGroup == lastexecuteGroup;
  wire              validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_43 = 8'h1 << instReg_vl[2:0];
  wire [7:0]        _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_43 | {_maskSplit_vlBoundaryCorrection_T_43[6:0], 1'h0};
  wire [7:0]        _vlBoundaryCorrection_T_8 = _vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[5:0], 2'h0};
  wire [7:0]        vlBoundaryCorrection = ~({8{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_8 | {_vlBoundaryCorrection_T_8[3:0], 4'h0})) & {8{validExecuteGroup}};
  wire [127:0]      selectReadStageMask_lo_lo_lo = {selectReadStageMask_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo};
  wire [127:0]      selectReadStageMask_lo_lo_hi = {selectReadStageMask_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo};
  wire [255:0]      selectReadStageMask_lo_lo = {selectReadStageMask_lo_lo_hi, selectReadStageMask_lo_lo_lo};
  wire [127:0]      selectReadStageMask_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo};
  wire [127:0]      selectReadStageMask_lo_hi_hi = {selectReadStageMask_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo};
  wire [255:0]      selectReadStageMask_lo_hi = {selectReadStageMask_lo_hi_hi, selectReadStageMask_lo_hi_lo};
  wire [511:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]      selectReadStageMask_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo};
  wire [127:0]      selectReadStageMask_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo};
  wire [255:0]      selectReadStageMask_hi_lo = {selectReadStageMask_hi_lo_hi, selectReadStageMask_hi_lo_lo};
  wire [127:0]      selectReadStageMask_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo};
  wire [127:0]      selectReadStageMask_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo};
  wire [255:0]      selectReadStageMask_hi_hi = {selectReadStageMask_hi_hi_hi, selectReadStageMask_hi_hi_lo};
  wire [511:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [127:0][7:0] _GEN_42 =
    {{selectReadStageMask_hi[511:504]},
     {selectReadStageMask_hi[503:496]},
     {selectReadStageMask_hi[495:488]},
     {selectReadStageMask_hi[487:480]},
     {selectReadStageMask_hi[479:472]},
     {selectReadStageMask_hi[471:464]},
     {selectReadStageMask_hi[463:456]},
     {selectReadStageMask_hi[455:448]},
     {selectReadStageMask_hi[447:440]},
     {selectReadStageMask_hi[439:432]},
     {selectReadStageMask_hi[431:424]},
     {selectReadStageMask_hi[423:416]},
     {selectReadStageMask_hi[415:408]},
     {selectReadStageMask_hi[407:400]},
     {selectReadStageMask_hi[399:392]},
     {selectReadStageMask_hi[391:384]},
     {selectReadStageMask_hi[383:376]},
     {selectReadStageMask_hi[375:368]},
     {selectReadStageMask_hi[367:360]},
     {selectReadStageMask_hi[359:352]},
     {selectReadStageMask_hi[351:344]},
     {selectReadStageMask_hi[343:336]},
     {selectReadStageMask_hi[335:328]},
     {selectReadStageMask_hi[327:320]},
     {selectReadStageMask_hi[319:312]},
     {selectReadStageMask_hi[311:304]},
     {selectReadStageMask_hi[303:296]},
     {selectReadStageMask_hi[295:288]},
     {selectReadStageMask_hi[287:280]},
     {selectReadStageMask_hi[279:272]},
     {selectReadStageMask_hi[271:264]},
     {selectReadStageMask_hi[263:256]},
     {selectReadStageMask_hi[255:248]},
     {selectReadStageMask_hi[247:240]},
     {selectReadStageMask_hi[239:232]},
     {selectReadStageMask_hi[231:224]},
     {selectReadStageMask_hi[223:216]},
     {selectReadStageMask_hi[215:208]},
     {selectReadStageMask_hi[207:200]},
     {selectReadStageMask_hi[199:192]},
     {selectReadStageMask_hi[191:184]},
     {selectReadStageMask_hi[183:176]},
     {selectReadStageMask_hi[175:168]},
     {selectReadStageMask_hi[167:160]},
     {selectReadStageMask_hi[159:152]},
     {selectReadStageMask_hi[151:144]},
     {selectReadStageMask_hi[143:136]},
     {selectReadStageMask_hi[135:128]},
     {selectReadStageMask_hi[127:120]},
     {selectReadStageMask_hi[119:112]},
     {selectReadStageMask_hi[111:104]},
     {selectReadStageMask_hi[103:96]},
     {selectReadStageMask_hi[95:88]},
     {selectReadStageMask_hi[87:80]},
     {selectReadStageMask_hi[79:72]},
     {selectReadStageMask_hi[71:64]},
     {selectReadStageMask_hi[63:56]},
     {selectReadStageMask_hi[55:48]},
     {selectReadStageMask_hi[47:40]},
     {selectReadStageMask_hi[39:32]},
     {selectReadStageMask_hi[31:24]},
     {selectReadStageMask_hi[23:16]},
     {selectReadStageMask_hi[15:8]},
     {selectReadStageMask_hi[7:0]},
     {selectReadStageMask_lo[511:504]},
     {selectReadStageMask_lo[503:496]},
     {selectReadStageMask_lo[495:488]},
     {selectReadStageMask_lo[487:480]},
     {selectReadStageMask_lo[479:472]},
     {selectReadStageMask_lo[471:464]},
     {selectReadStageMask_lo[463:456]},
     {selectReadStageMask_lo[455:448]},
     {selectReadStageMask_lo[447:440]},
     {selectReadStageMask_lo[439:432]},
     {selectReadStageMask_lo[431:424]},
     {selectReadStageMask_lo[423:416]},
     {selectReadStageMask_lo[415:408]},
     {selectReadStageMask_lo[407:400]},
     {selectReadStageMask_lo[399:392]},
     {selectReadStageMask_lo[391:384]},
     {selectReadStageMask_lo[383:376]},
     {selectReadStageMask_lo[375:368]},
     {selectReadStageMask_lo[367:360]},
     {selectReadStageMask_lo[359:352]},
     {selectReadStageMask_lo[351:344]},
     {selectReadStageMask_lo[343:336]},
     {selectReadStageMask_lo[335:328]},
     {selectReadStageMask_lo[327:320]},
     {selectReadStageMask_lo[319:312]},
     {selectReadStageMask_lo[311:304]},
     {selectReadStageMask_lo[303:296]},
     {selectReadStageMask_lo[295:288]},
     {selectReadStageMask_lo[287:280]},
     {selectReadStageMask_lo[279:272]},
     {selectReadStageMask_lo[271:264]},
     {selectReadStageMask_lo[263:256]},
     {selectReadStageMask_lo[255:248]},
     {selectReadStageMask_lo[247:240]},
     {selectReadStageMask_lo[239:232]},
     {selectReadStageMask_lo[231:224]},
     {selectReadStageMask_lo[223:216]},
     {selectReadStageMask_lo[215:208]},
     {selectReadStageMask_lo[207:200]},
     {selectReadStageMask_lo[199:192]},
     {selectReadStageMask_lo[191:184]},
     {selectReadStageMask_lo[183:176]},
     {selectReadStageMask_lo[175:168]},
     {selectReadStageMask_lo[167:160]},
     {selectReadStageMask_lo[159:152]},
     {selectReadStageMask_lo[151:144]},
     {selectReadStageMask_lo[143:136]},
     {selectReadStageMask_lo[135:128]},
     {selectReadStageMask_lo[127:120]},
     {selectReadStageMask_lo[119:112]},
     {selectReadStageMask_lo[111:104]},
     {selectReadStageMask_lo[103:96]},
     {selectReadStageMask_lo[95:88]},
     {selectReadStageMask_lo[87:80]},
     {selectReadStageMask_lo[79:72]},
     {selectReadStageMask_lo[71:64]},
     {selectReadStageMask_lo[63:56]},
     {selectReadStageMask_lo[55:48]},
     {selectReadStageMask_lo[47:40]},
     {selectReadStageMask_lo[39:32]},
     {selectReadStageMask_lo[31:24]},
     {selectReadStageMask_lo[23:16]},
     {selectReadStageMask_lo[15:8]},
     {selectReadStageMask_lo[7:0]}};
  wire [7:0]        readMaskCorrection = (instReg_maskType ? _GEN_42[executeGroup[6:0]] : 8'hFF) & vlBoundaryCorrection;
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo};
  wire [255:0]      maskSplit_maskSelect_lo_lo = {maskSplit_maskSelect_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo};
  wire [255:0]      maskSplit_maskSelect_lo_hi = {maskSplit_maskSelect_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo};
  wire [511:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo};
  wire [255:0]      maskSplit_maskSelect_hi_lo = {maskSplit_maskSelect_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo};
  wire [255:0]      maskSplit_maskSelect_hi_hi = {maskSplit_maskSelect_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo};
  wire [511:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [5:0]        executeGroupCounter;
  wire              maskSplit_vlMisAlign = |(instReg_vl[4:0]);
  wire [5:0]        maskSplit_lastexecuteGroup = instReg_vl[10:5] - {5'h0, ~maskSplit_vlMisAlign};
  wire              maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire              maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_2 = 32'h1 << instReg_vl[4:0];
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[30:0], 1'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[29:0], 2'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[27:0], 4'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_14 = _maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[23:0], 8'h0};
  wire [31:0]       maskSplit_vlBoundaryCorrection = ~({32{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_14 | {_maskSplit_vlBoundaryCorrection_T_14[15:0], 16'h0})) & {32{maskSplit_validExecuteGroup}};
  wire [31:0][31:0] _GEN_43 =
    {{maskSplit_maskSelect_hi[511:480]},
     {maskSplit_maskSelect_hi[479:448]},
     {maskSplit_maskSelect_hi[447:416]},
     {maskSplit_maskSelect_hi[415:384]},
     {maskSplit_maskSelect_hi[383:352]},
     {maskSplit_maskSelect_hi[351:320]},
     {maskSplit_maskSelect_hi[319:288]},
     {maskSplit_maskSelect_hi[287:256]},
     {maskSplit_maskSelect_hi[255:224]},
     {maskSplit_maskSelect_hi[223:192]},
     {maskSplit_maskSelect_hi[191:160]},
     {maskSplit_maskSelect_hi[159:128]},
     {maskSplit_maskSelect_hi[127:96]},
     {maskSplit_maskSelect_hi[95:64]},
     {maskSplit_maskSelect_hi[63:32]},
     {maskSplit_maskSelect_hi[31:0]},
     {maskSplit_maskSelect_lo[511:480]},
     {maskSplit_maskSelect_lo[479:448]},
     {maskSplit_maskSelect_lo[447:416]},
     {maskSplit_maskSelect_lo[415:384]},
     {maskSplit_maskSelect_lo[383:352]},
     {maskSplit_maskSelect_lo[351:320]},
     {maskSplit_maskSelect_lo[319:288]},
     {maskSplit_maskSelect_lo[287:256]},
     {maskSplit_maskSelect_lo[255:224]},
     {maskSplit_maskSelect_lo[223:192]},
     {maskSplit_maskSelect_lo[191:160]},
     {maskSplit_maskSelect_lo[159:128]},
     {maskSplit_maskSelect_lo[127:96]},
     {maskSplit_maskSelect_lo[95:64]},
     {maskSplit_maskSelect_lo[63:32]},
     {maskSplit_maskSelect_lo[31:0]}};
  wire [31:0]       maskSplit_0_2 = (instReg_maskType ? _GEN_43[executeGroupCounter[4:0]] : 32'hFFFFFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]        maskSplit_byteMask_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]        maskSplit_byteMask_lo_lo_hi = {maskSplit_byteMask_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]        maskSplit_byteMask_lo_hi_lo = {maskSplit_byteMask_lo_hi_lo_hi, maskSplit_byteMask_lo_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]        maskSplit_byteMask_lo_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [15:0]       maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_lo = maskSplit_0_2[17:16];
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_hi = maskSplit_0_2[19:18];
  wire [3:0]        maskSplit_byteMask_hi_lo_lo = {maskSplit_byteMask_hi_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_lo = maskSplit_0_2[21:20];
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_hi = maskSplit_0_2[23:22];
  wire [3:0]        maskSplit_byteMask_hi_lo_hi = {maskSplit_byteMask_hi_lo_hi_hi, maskSplit_byteMask_hi_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_lo = maskSplit_0_2[25:24];
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_hi = maskSplit_0_2[27:26];
  wire [3:0]        maskSplit_byteMask_hi_hi_lo = {maskSplit_byteMask_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_lo = maskSplit_0_2[29:28];
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_hi = maskSplit_0_2[31:30];
  wire [3:0]        maskSplit_byteMask_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [15:0]       maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [31:0]       maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_1};
  wire [511:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_1};
  wire [511:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire              maskSplit_vlMisAlign_1 = |(instReg_vl[3:0]);
  wire [6:0]        maskSplit_lastexecuteGroup_1 = instReg_vl[10:4] - {6'h0, ~maskSplit_vlMisAlign_1};
  wire [6:0]        _GEN_44 = {1'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_1 = _GEN_44 == maskSplit_lastexecuteGroup_1;
  wire              maskSplit_validExecuteGroup_1 = _GEN_44 <= maskSplit_lastexecuteGroup_1;
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_24 = 16'h1 << instReg_vl[3:0];
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_27 = _maskSplit_vlBoundaryCorrection_T_24 | {_maskSplit_vlBoundaryCorrection_T_24[14:0], 1'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_30 = _maskSplit_vlBoundaryCorrection_T_27 | {_maskSplit_vlBoundaryCorrection_T_27[13:0], 2'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_33 = _maskSplit_vlBoundaryCorrection_T_30 | {_maskSplit_vlBoundaryCorrection_T_30[11:0], 4'h0};
  wire [15:0]       maskSplit_vlBoundaryCorrection_1 =
    ~({16{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_33 | {_maskSplit_vlBoundaryCorrection_T_33[7:0], 8'h0})) & {16{maskSplit_validExecuteGroup_1}};
  wire [63:0][15:0] _GEN_45 =
    {{maskSplit_maskSelect_hi_1[511:496]},
     {maskSplit_maskSelect_hi_1[495:480]},
     {maskSplit_maskSelect_hi_1[479:464]},
     {maskSplit_maskSelect_hi_1[463:448]},
     {maskSplit_maskSelect_hi_1[447:432]},
     {maskSplit_maskSelect_hi_1[431:416]},
     {maskSplit_maskSelect_hi_1[415:400]},
     {maskSplit_maskSelect_hi_1[399:384]},
     {maskSplit_maskSelect_hi_1[383:368]},
     {maskSplit_maskSelect_hi_1[367:352]},
     {maskSplit_maskSelect_hi_1[351:336]},
     {maskSplit_maskSelect_hi_1[335:320]},
     {maskSplit_maskSelect_hi_1[319:304]},
     {maskSplit_maskSelect_hi_1[303:288]},
     {maskSplit_maskSelect_hi_1[287:272]},
     {maskSplit_maskSelect_hi_1[271:256]},
     {maskSplit_maskSelect_hi_1[255:240]},
     {maskSplit_maskSelect_hi_1[239:224]},
     {maskSplit_maskSelect_hi_1[223:208]},
     {maskSplit_maskSelect_hi_1[207:192]},
     {maskSplit_maskSelect_hi_1[191:176]},
     {maskSplit_maskSelect_hi_1[175:160]},
     {maskSplit_maskSelect_hi_1[159:144]},
     {maskSplit_maskSelect_hi_1[143:128]},
     {maskSplit_maskSelect_hi_1[127:112]},
     {maskSplit_maskSelect_hi_1[111:96]},
     {maskSplit_maskSelect_hi_1[95:80]},
     {maskSplit_maskSelect_hi_1[79:64]},
     {maskSplit_maskSelect_hi_1[63:48]},
     {maskSplit_maskSelect_hi_1[47:32]},
     {maskSplit_maskSelect_hi_1[31:16]},
     {maskSplit_maskSelect_hi_1[15:0]},
     {maskSplit_maskSelect_lo_1[511:496]},
     {maskSplit_maskSelect_lo_1[495:480]},
     {maskSplit_maskSelect_lo_1[479:464]},
     {maskSplit_maskSelect_lo_1[463:448]},
     {maskSplit_maskSelect_lo_1[447:432]},
     {maskSplit_maskSelect_lo_1[431:416]},
     {maskSplit_maskSelect_lo_1[415:400]},
     {maskSplit_maskSelect_lo_1[399:384]},
     {maskSplit_maskSelect_lo_1[383:368]},
     {maskSplit_maskSelect_lo_1[367:352]},
     {maskSplit_maskSelect_lo_1[351:336]},
     {maskSplit_maskSelect_lo_1[335:320]},
     {maskSplit_maskSelect_lo_1[319:304]},
     {maskSplit_maskSelect_lo_1[303:288]},
     {maskSplit_maskSelect_lo_1[287:272]},
     {maskSplit_maskSelect_lo_1[271:256]},
     {maskSplit_maskSelect_lo_1[255:240]},
     {maskSplit_maskSelect_lo_1[239:224]},
     {maskSplit_maskSelect_lo_1[223:208]},
     {maskSplit_maskSelect_lo_1[207:192]},
     {maskSplit_maskSelect_lo_1[191:176]},
     {maskSplit_maskSelect_lo_1[175:160]},
     {maskSplit_maskSelect_lo_1[159:144]},
     {maskSplit_maskSelect_lo_1[143:128]},
     {maskSplit_maskSelect_lo_1[127:112]},
     {maskSplit_maskSelect_lo_1[111:96]},
     {maskSplit_maskSelect_lo_1[95:80]},
     {maskSplit_maskSelect_lo_1[79:64]},
     {maskSplit_maskSelect_lo_1[63:48]},
     {maskSplit_maskSelect_lo_1[47:32]},
     {maskSplit_maskSelect_lo_1[31:16]},
     {maskSplit_maskSelect_lo_1[15:0]}};
  wire [15:0]       maskSplit_1_2 = (instReg_maskType ? _GEN_45[executeGroupCounter] : 16'hFFFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]        maskSplit_byteMask_lo_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]        maskSplit_byteMask_lo_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]        maskSplit_byteMask_lo_lo_1 = {maskSplit_byteMask_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_lo_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]        maskSplit_byteMask_lo_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]        maskSplit_byteMask_lo_hi_1 = {maskSplit_byteMask_lo_hi_hi_1, maskSplit_byteMask_lo_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_lo_lo_1 = {{2{maskSplit_1_2[9]}}, {2{maskSplit_1_2[8]}}};
  wire [3:0]        maskSplit_byteMask_hi_lo_hi_1 = {{2{maskSplit_1_2[11]}}, {2{maskSplit_1_2[10]}}};
  wire [7:0]        maskSplit_byteMask_hi_lo_1 = {maskSplit_byteMask_hi_lo_hi_1, maskSplit_byteMask_hi_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_hi_lo_1 = {{2{maskSplit_1_2[13]}}, {2{maskSplit_1_2[12]}}};
  wire [3:0]        maskSplit_byteMask_hi_hi_hi_1 = {{2{maskSplit_1_2[15]}}, {2{maskSplit_1_2[14]}}};
  wire [7:0]        maskSplit_byteMask_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_1, maskSplit_byteMask_hi_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [31:0]       maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_2};
  wire [511:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_2};
  wire [511:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire              maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[2:0]);
  wire [7:0]        maskSplit_lastexecuteGroup_2 = instReg_vl[10:3] - {7'h0, ~maskSplit_vlMisAlign_2};
  wire [7:0]        _GEN_46 = {2'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_2 = _GEN_46 == maskSplit_lastexecuteGroup_2;
  wire              maskSplit_validExecuteGroup_2 = _GEN_46 <= maskSplit_lastexecuteGroup_2;
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_46 = _maskSplit_vlBoundaryCorrection_T_43 | {_maskSplit_vlBoundaryCorrection_T_43[6:0], 1'h0};
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_49 = _maskSplit_vlBoundaryCorrection_T_46 | {_maskSplit_vlBoundaryCorrection_T_46[5:0], 2'h0};
  wire [7:0]        maskSplit_vlBoundaryCorrection_2 =
    ~({8{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_49 | {_maskSplit_vlBoundaryCorrection_T_49[3:0], 4'h0})) & {8{maskSplit_validExecuteGroup_2}};
  wire [63:0][7:0]  _GEN_47 =
    {{maskSplit_maskSelect_lo_2[511:504]},
     {maskSplit_maskSelect_lo_2[503:496]},
     {maskSplit_maskSelect_lo_2[495:488]},
     {maskSplit_maskSelect_lo_2[487:480]},
     {maskSplit_maskSelect_lo_2[479:472]},
     {maskSplit_maskSelect_lo_2[471:464]},
     {maskSplit_maskSelect_lo_2[463:456]},
     {maskSplit_maskSelect_lo_2[455:448]},
     {maskSplit_maskSelect_lo_2[447:440]},
     {maskSplit_maskSelect_lo_2[439:432]},
     {maskSplit_maskSelect_lo_2[431:424]},
     {maskSplit_maskSelect_lo_2[423:416]},
     {maskSplit_maskSelect_lo_2[415:408]},
     {maskSplit_maskSelect_lo_2[407:400]},
     {maskSplit_maskSelect_lo_2[399:392]},
     {maskSplit_maskSelect_lo_2[391:384]},
     {maskSplit_maskSelect_lo_2[383:376]},
     {maskSplit_maskSelect_lo_2[375:368]},
     {maskSplit_maskSelect_lo_2[367:360]},
     {maskSplit_maskSelect_lo_2[359:352]},
     {maskSplit_maskSelect_lo_2[351:344]},
     {maskSplit_maskSelect_lo_2[343:336]},
     {maskSplit_maskSelect_lo_2[335:328]},
     {maskSplit_maskSelect_lo_2[327:320]},
     {maskSplit_maskSelect_lo_2[319:312]},
     {maskSplit_maskSelect_lo_2[311:304]},
     {maskSplit_maskSelect_lo_2[303:296]},
     {maskSplit_maskSelect_lo_2[295:288]},
     {maskSplit_maskSelect_lo_2[287:280]},
     {maskSplit_maskSelect_lo_2[279:272]},
     {maskSplit_maskSelect_lo_2[271:264]},
     {maskSplit_maskSelect_lo_2[263:256]},
     {maskSplit_maskSelect_lo_2[255:248]},
     {maskSplit_maskSelect_lo_2[247:240]},
     {maskSplit_maskSelect_lo_2[239:232]},
     {maskSplit_maskSelect_lo_2[231:224]},
     {maskSplit_maskSelect_lo_2[223:216]},
     {maskSplit_maskSelect_lo_2[215:208]},
     {maskSplit_maskSelect_lo_2[207:200]},
     {maskSplit_maskSelect_lo_2[199:192]},
     {maskSplit_maskSelect_lo_2[191:184]},
     {maskSplit_maskSelect_lo_2[183:176]},
     {maskSplit_maskSelect_lo_2[175:168]},
     {maskSplit_maskSelect_lo_2[167:160]},
     {maskSplit_maskSelect_lo_2[159:152]},
     {maskSplit_maskSelect_lo_2[151:144]},
     {maskSplit_maskSelect_lo_2[143:136]},
     {maskSplit_maskSelect_lo_2[135:128]},
     {maskSplit_maskSelect_lo_2[127:120]},
     {maskSplit_maskSelect_lo_2[119:112]},
     {maskSplit_maskSelect_lo_2[111:104]},
     {maskSplit_maskSelect_lo_2[103:96]},
     {maskSplit_maskSelect_lo_2[95:88]},
     {maskSplit_maskSelect_lo_2[87:80]},
     {maskSplit_maskSelect_lo_2[79:72]},
     {maskSplit_maskSelect_lo_2[71:64]},
     {maskSplit_maskSelect_lo_2[63:56]},
     {maskSplit_maskSelect_lo_2[55:48]},
     {maskSplit_maskSelect_lo_2[47:40]},
     {maskSplit_maskSelect_lo_2[39:32]},
     {maskSplit_maskSelect_lo_2[31:24]},
     {maskSplit_maskSelect_lo_2[23:16]},
     {maskSplit_maskSelect_lo_2[15:8]},
     {maskSplit_maskSelect_lo_2[7:0]}};
  wire [7:0]        maskSplit_2_2 = (instReg_maskType ? _GEN_47[executeGroupCounter] : 8'hFF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]        maskSplit_byteMask_lo_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]        maskSplit_byteMask_lo_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]       maskSplit_byteMask_lo_2 = {maskSplit_byteMask_lo_hi_2, maskSplit_byteMask_lo_lo_2};
  wire [7:0]        maskSplit_byteMask_hi_lo_2 = {{4{maskSplit_2_2[5]}}, {4{maskSplit_2_2[4]}}};
  wire [7:0]        maskSplit_byteMask_hi_hi_2 = {{4{maskSplit_2_2[7]}}, {4{maskSplit_2_2[6]}}};
  wire [15:0]       maskSplit_byteMask_hi_2 = {maskSplit_byteMask_hi_hi_2, maskSplit_byteMask_hi_lo_2};
  wire [31:0]       maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [31:0]       executeByteMask = (sew1H[0] ? maskSplit_0_1 : 32'h0) | (sew1H[1] ? maskSplit_1_1 : 32'h0) | (sew1H[2] ? maskSplit_2_1 : 32'h0);
  wire [31:0]       _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 32'h0;
  wire [15:0]       _GEN_48 = _executeElementMask_T_3[15:0] | (sew1H[1] ? maskSplit_1_2 : 16'h0);
  wire [31:0]       executeElementMask = {_executeElementMask_T_3[31:16], _GEN_48[15:8], _GEN_48[7:0] | (sew1H[2] ? maskSplit_2_2 : 8'h0)};
  wire [127:0]      maskForDestination_lo_lo_lo = {maskForDestination_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo};
  wire [127:0]      maskForDestination_lo_lo_hi = {maskForDestination_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo};
  wire [255:0]      maskForDestination_lo_lo = {maskForDestination_lo_lo_hi, maskForDestination_lo_lo_lo};
  wire [127:0]      maskForDestination_lo_hi_lo = {maskForDestination_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo};
  wire [127:0]      maskForDestination_lo_hi_hi = {maskForDestination_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo};
  wire [255:0]      maskForDestination_lo_hi = {maskForDestination_lo_hi_hi, maskForDestination_lo_hi_lo};
  wire [511:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]      maskForDestination_hi_lo_lo = {maskForDestination_hi_lo_lo_hi, maskForDestination_hi_lo_lo_lo};
  wire [127:0]      maskForDestination_hi_lo_hi = {maskForDestination_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo};
  wire [255:0]      maskForDestination_hi_lo = {maskForDestination_hi_lo_hi, maskForDestination_hi_lo_lo};
  wire [127:0]      maskForDestination_hi_hi_lo = {maskForDestination_hi_hi_lo_hi, maskForDestination_hi_hi_lo_lo};
  wire [127:0]      maskForDestination_hi_hi_hi = {maskForDestination_hi_hi_hi_hi, maskForDestination_hi_hi_hi_lo};
  wire [255:0]      maskForDestination_hi_hi = {maskForDestination_hi_hi_hi, maskForDestination_hi_hi_lo};
  wire [511:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire [1:0]        vs1Split_vs1SetIndex_1 = requestCounter[1:0];
  wire [255:0]      _lastGroupMask_T = 256'h1 << elementTailForMaskDestination;
  wire [254:0]      _GEN_49 = _lastGroupMask_T[254:0] | _lastGroupMask_T[255:1];
  wire [253:0]      _GEN_50 = _GEN_49[253:0] | {_lastGroupMask_T[255], _GEN_49[254:2]};
  wire [251:0]      _GEN_51 = _GEN_50[251:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:4]};
  wire [247:0]      _GEN_52 = _GEN_51[247:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:252], _GEN_51[251:8]};
  wire [239:0]      _GEN_53 = _GEN_52[239:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:252], _GEN_51[251:248], _GEN_52[247:16]};
  wire [223:0]      _GEN_54 = _GEN_53[223:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:252], _GEN_51[251:248], _GEN_52[247:240], _GEN_53[239:32]};
  wire [191:0]      _GEN_55 = _GEN_54[191:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:252], _GEN_51[251:248], _GEN_52[247:240], _GEN_53[239:224], _GEN_54[223:64]};
  wire [255:0]      lastGroupMask =
    {_lastGroupMask_T[255],
     _GEN_49[254],
     _GEN_50[253:252],
     _GEN_51[251:248],
     _GEN_52[247:240],
     _GEN_53[239:224],
     _GEN_54[223:192],
     _GEN_55[191:128],
     _GEN_55[127:0] | {_lastGroupMask_T[255], _GEN_49[254], _GEN_50[253:252], _GEN_51[251:248], _GEN_52[247:240], _GEN_53[239:224], _GEN_54[223:192], _GEN_55[191:128]}};
  wire [3:0][255:0] _GEN_56 = {{maskForDestination_hi[511:256]}, {maskForDestination_hi[255:0]}, {maskForDestination_lo[511:256]}, {maskForDestination_lo[255:0]}};
  wire [255:0]      currentMaskGroupForDestination =
    (lastGroup ? lastGroupMask : 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
    & (instReg_maskType & ~instReg_decodeResult_maskSource ? _GEN_56[vs1Split_vs1SetIndex_1] : 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]       _GEN_57 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]       groupSourceData_lo_lo;
  assign groupSourceData_lo_lo = _GEN_57;
  wire [63:0]       source1_lo_lo;
  assign source1_lo_lo = _GEN_57;
  wire [63:0]       _GEN_58 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]       groupSourceData_lo_hi;
  assign groupSourceData_lo_hi = _GEN_58;
  wire [63:0]       source1_lo_hi;
  assign source1_lo_hi = _GEN_58;
  wire [127:0]      groupSourceData_lo = {groupSourceData_lo_hi, groupSourceData_lo_lo};
  wire [63:0]       _GEN_59 = {exeReqReg_5_bits_source1, exeReqReg_4_bits_source1};
  wire [63:0]       groupSourceData_hi_lo;
  assign groupSourceData_hi_lo = _GEN_59;
  wire [63:0]       source1_hi_lo;
  assign source1_hi_lo = _GEN_59;
  wire [63:0]       _GEN_60 = {exeReqReg_7_bits_source1, exeReqReg_6_bits_source1};
  wire [63:0]       groupSourceData_hi_hi;
  assign groupSourceData_hi_hi = _GEN_60;
  wire [63:0]       source1_hi_hi;
  assign source1_hi_hi = _GEN_60;
  wire [127:0]      groupSourceData_hi = {groupSourceData_hi_hi, groupSourceData_hi_lo};
  wire [255:0]      groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]        _GEN_61 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]        groupSourceValid_lo_lo;
  assign groupSourceValid_lo_lo = _GEN_61;
  wire [1:0]        view__in_bits_validInput_lo_lo;
  assign view__in_bits_validInput_lo_lo = _GEN_61;
  wire [1:0]        view__in_bits_sourceValid_lo_lo;
  assign view__in_bits_sourceValid_lo_lo = _GEN_61;
  wire [1:0]        _GEN_62 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]        groupSourceValid_lo_hi;
  assign groupSourceValid_lo_hi = _GEN_62;
  wire [1:0]        view__in_bits_validInput_lo_hi;
  assign view__in_bits_validInput_lo_hi = _GEN_62;
  wire [1:0]        view__in_bits_sourceValid_lo_hi;
  assign view__in_bits_sourceValid_lo_hi = _GEN_62;
  wire [3:0]        groupSourceValid_lo = {groupSourceValid_lo_hi, groupSourceValid_lo_lo};
  wire [1:0]        _GEN_63 = {exeReqReg_5_valid, exeReqReg_4_valid};
  wire [1:0]        groupSourceValid_hi_lo;
  assign groupSourceValid_hi_lo = _GEN_63;
  wire [1:0]        view__in_bits_validInput_hi_lo;
  assign view__in_bits_validInput_hi_lo = _GEN_63;
  wire [1:0]        view__in_bits_sourceValid_hi_lo;
  assign view__in_bits_sourceValid_hi_lo = _GEN_63;
  wire [1:0]        _GEN_64 = {exeReqReg_7_valid, exeReqReg_6_valid};
  wire [1:0]        groupSourceValid_hi_hi;
  assign groupSourceValid_hi_hi = _GEN_64;
  wire [1:0]        view__in_bits_validInput_hi_hi;
  assign view__in_bits_validInput_hi_hi = _GEN_64;
  wire [1:0]        view__in_bits_sourceValid_hi_hi;
  assign view__in_bits_sourceValid_hi_hi = _GEN_64;
  wire [3:0]        groupSourceValid_hi = {groupSourceValid_hi_hi, groupSourceValid_hi_lo};
  wire [7:0]        groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]        shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]        _shifterSource_T = 4'h1 << shifterSize;
  wire [255:0]      _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 256'h0;
  wire [191:0]      _GEN_65 = _shifterSource_T_8[191:0] | (_shifterSource_T[1] ? groupSourceData[255:64] : 192'h0);
  wire [127:0]      _GEN_66 = _GEN_65[127:0] | (_shifterSource_T[2] ? groupSourceData[255:128] : 128'h0);
  wire [255:0]      shifterSource = {_shifterSource_T_8[255:192], _GEN_65[191:128], _GEN_66[127:64], _GEN_66[63:0] | (_shifterSource_T[3] ? groupSourceData[255:192] : 64'h0)};
  wire [7:0]        selectValid_lo_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]        selectValid_lo_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [15:0]       selectValid_lo = {selectValid_lo_hi, selectValid_lo_lo};
  wire [7:0]        selectValid_hi_lo = {{4{groupSourceValid[5]}}, {4{groupSourceValid[4]}}};
  wire [7:0]        selectValid_hi_hi = {{4{groupSourceValid[7]}}, {4{groupSourceValid[6]}}};
  wire [15:0]       selectValid_hi = {selectValid_hi_hi, selectValid_hi_lo};
  wire [3:0]        selectValid_lo_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]        selectValid_lo_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [7:0]        selectValid_lo_1 = {selectValid_lo_hi_1, selectValid_lo_lo_1};
  wire [3:0]        selectValid_hi_lo_1 = {{2{groupSourceValid[5]}}, {2{groupSourceValid[4]}}};
  wire [3:0]        selectValid_hi_hi_1 = {{2{groupSourceValid[7]}}, {2{groupSourceValid[6]}}};
  wire [7:0]        selectValid_hi_1 = {selectValid_hi_hi_1, selectValid_hi_lo_1};
  wire [3:0][7:0]   _GEN_67 = {{selectValid_hi[15:8]}, {selectValid_hi[7:0]}, {selectValid_lo[15:8]}, {selectValid_lo[7:0]}};
  wire [7:0]        selectValid = (sourceDataEEW1H[0] ? _GEN_67[executeIndex] : 8'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 8'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 8'h0);
  wire [31:0]       source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]       source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]       source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]       source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [31:0]       source_4 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[39:32] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[79:64] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[159:128] : 32'h0);
  wire [31:0]       source_5 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[47:40] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[95:80] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[191:160] : 32'h0);
  wire [31:0]       source_6 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[55:48] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[111:96] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[223:192] : 32'h0);
  wire [31:0]       source_7 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[63:56] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[127:112] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[255:224] : 32'h0);
  wire [7:0]        _GEN_68 = selectValid & readMaskCorrection;
  wire [7:0]        checkVec_validVec;
  assign checkVec_validVec = _GEN_68;
  wire [7:0]        checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_68;
  wire [7:0]        checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_68;
  wire              checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]        _GEN_69 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]        checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_12;
  assign checkVec_checkResultVec_intLMULInput_12 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_13;
  assign checkVec_checkResultVec_intLMULInput_13 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_14;
  assign checkVec_checkResultVec_intLMULInput_14 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_15;
  assign checkVec_checkResultVec_intLMULInput_15 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_16;
  assign checkVec_checkResultVec_intLMULInput_16 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_17;
  assign checkVec_checkResultVec_intLMULInput_17 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_18;
  assign checkVec_checkResultVec_intLMULInput_18 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_19;
  assign checkVec_checkResultVec_intLMULInput_19 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_20;
  assign checkVec_checkResultVec_intLMULInput_20 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_21;
  assign checkVec_checkResultVec_intLMULInput_21 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_22;
  assign checkVec_checkResultVec_intLMULInput_22 = _GEN_69;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_23;
  assign checkVec_checkResultVec_intLMULInput_23 = _GEN_69;
  wire [9:0]        checkVec_checkResultVec_dataPosition = source_0[9:0];
  wire [3:0]        checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]        checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [2:0]        checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[9:5];
  wire [1:0]        checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[4:2];
  wire [2:0]        checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [4:0]        checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]        checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion[4:2];
  wire              checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:10]};
  wire              checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire              checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_1 = source_1[9:0];
  wire [3:0]        checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]        checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [2:0]        checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[9:5];
  wire [1:0]        checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[4:2];
  wire [2:0]        checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]        checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1[4:2];
  wire              checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:10]};
  wire              checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire              checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_2 = source_2[9:0];
  wire [3:0]        checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]        checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [2:0]        checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[9:5];
  wire [1:0]        checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[4:2];
  wire [2:0]        checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2[4:2];
  wire              checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:10]};
  wire              checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire              checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_3 = source_3[9:0];
  wire [3:0]        checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]        checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [2:0]        checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[9:5];
  wire [1:0]        checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[4:2];
  wire [2:0]        checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]        checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3[4:2];
  wire              checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:10]};
  wire              checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire              checkVec_checkResultVec_4_6 = checkVec_validVec[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_4 = source_4[9:0];
  wire [3:0]        checkVec_checkResultVec_4_0 = 4'h1 << checkVec_checkResultVec_dataPosition_4[1:0];
  wire [1:0]        checkVec_checkResultVec_4_1 = checkVec_checkResultVec_dataPosition_4[1:0];
  wire [2:0]        checkVec_checkResultVec_4_2 = checkVec_checkResultVec_dataPosition_4[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[9:5];
  wire [1:0]        checkVec_checkResultVec_4_3 = checkVec_checkResultVec_dataGroup_4[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[4:2];
  wire [2:0]        checkVec_checkResultVec_4_4 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_4_3, checkVec_checkResultVec_4_2};
  wire [2:0]        checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4[4:2];
  wire              checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_4[31:10]};
  wire              checkVec_checkResultVec_4_5 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_4_6;
  wire              checkVec_checkResultVec_5_6 = checkVec_validVec[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_5 = source_5[9:0];
  wire [3:0]        checkVec_checkResultVec_5_0 = 4'h1 << checkVec_checkResultVec_dataPosition_5[1:0];
  wire [1:0]        checkVec_checkResultVec_5_1 = checkVec_checkResultVec_dataPosition_5[1:0];
  wire [2:0]        checkVec_checkResultVec_5_2 = checkVec_checkResultVec_dataPosition_5[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[9:5];
  wire [1:0]        checkVec_checkResultVec_5_3 = checkVec_checkResultVec_dataGroup_5[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[4:2];
  wire [2:0]        checkVec_checkResultVec_5_4 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_5_2};
  wire [2:0]        checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5[4:2];
  wire              checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_5[31:10]};
  wire              checkVec_checkResultVec_5_5 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_5_6;
  wire              checkVec_checkResultVec_6_6 = checkVec_validVec[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_6 = source_6[9:0];
  wire [3:0]        checkVec_checkResultVec_6_0 = 4'h1 << checkVec_checkResultVec_dataPosition_6[1:0];
  wire [1:0]        checkVec_checkResultVec_6_1 = checkVec_checkResultVec_dataPosition_6[1:0];
  wire [2:0]        checkVec_checkResultVec_6_2 = checkVec_checkResultVec_dataPosition_6[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[9:5];
  wire [1:0]        checkVec_checkResultVec_6_3 = checkVec_checkResultVec_dataGroup_6[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[4:2];
  wire [2:0]        checkVec_checkResultVec_6_4 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_6_3, checkVec_checkResultVec_6_2};
  wire [2:0]        checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6[4:2];
  wire              checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_6[31:10]};
  wire              checkVec_checkResultVec_6_5 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_6_6;
  wire              checkVec_checkResultVec_7_6 = checkVec_validVec[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_7 = source_7[9:0];
  wire [3:0]        checkVec_checkResultVec_7_0 = 4'h1 << checkVec_checkResultVec_dataPosition_7[1:0];
  wire [1:0]        checkVec_checkResultVec_7_1 = checkVec_checkResultVec_dataPosition_7[1:0];
  wire [2:0]        checkVec_checkResultVec_7_2 = checkVec_checkResultVec_dataPosition_7[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[9:5];
  wire [1:0]        checkVec_checkResultVec_7_3 = checkVec_checkResultVec_dataGroup_7[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[4:2];
  wire [2:0]        checkVec_checkResultVec_7_4 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_7_2};
  wire [2:0]        checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7[4:2];
  wire              checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_7[31:10]};
  wire              checkVec_checkResultVec_7_5 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_7_6;
  wire [7:0]        checkVec_checkResult_lo_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]        checkVec_checkResult_lo_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]       checkVec_checkResult_lo = {checkVec_checkResult_lo_hi, checkVec_checkResult_lo_lo};
  wire [7:0]        checkVec_checkResult_hi_lo = {checkVec_checkResultVec_5_0, checkVec_checkResultVec_4_0};
  wire [7:0]        checkVec_checkResult_hi_hi = {checkVec_checkResultVec_7_0, checkVec_checkResultVec_6_0};
  wire [15:0]       checkVec_checkResult_hi = {checkVec_checkResult_hi_hi, checkVec_checkResult_hi_lo};
  wire [31:0]       checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]        checkVec_checkResult_lo_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]        checkVec_checkResult_lo_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]        checkVec_checkResult_lo_1 = {checkVec_checkResult_lo_hi_1, checkVec_checkResult_lo_lo_1};
  wire [3:0]        checkVec_checkResult_hi_lo_1 = {checkVec_checkResultVec_5_1, checkVec_checkResultVec_4_1};
  wire [3:0]        checkVec_checkResult_hi_hi_1 = {checkVec_checkResultVec_7_1, checkVec_checkResultVec_6_1};
  wire [7:0]        checkVec_checkResult_hi_1 = {checkVec_checkResult_hi_hi_1, checkVec_checkResult_hi_lo_1};
  wire [15:0]       checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [5:0]        checkVec_checkResult_lo_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [5:0]        checkVec_checkResult_lo_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [11:0]       checkVec_checkResult_lo_2 = {checkVec_checkResult_lo_hi_2, checkVec_checkResult_lo_lo_2};
  wire [5:0]        checkVec_checkResult_hi_lo_2 = {checkVec_checkResultVec_5_2, checkVec_checkResultVec_4_2};
  wire [5:0]        checkVec_checkResult_hi_hi_2 = {checkVec_checkResultVec_7_2, checkVec_checkResultVec_6_2};
  wire [11:0]       checkVec_checkResult_hi_2 = {checkVec_checkResult_hi_hi_2, checkVec_checkResult_hi_lo_2};
  wire [23:0]       checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [3:0]        checkVec_checkResult_lo_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [3:0]        checkVec_checkResult_lo_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [7:0]        checkVec_checkResult_lo_3 = {checkVec_checkResult_lo_hi_3, checkVec_checkResult_lo_lo_3};
  wire [3:0]        checkVec_checkResult_hi_lo_3 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_4_3};
  wire [3:0]        checkVec_checkResult_hi_hi_3 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_6_3};
  wire [7:0]        checkVec_checkResult_hi_3 = {checkVec_checkResult_hi_hi_3, checkVec_checkResult_hi_lo_3};
  wire [15:0]       checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]        checkVec_checkResult_lo_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]        checkVec_checkResult_lo_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]       checkVec_checkResult_lo_4 = {checkVec_checkResult_lo_hi_4, checkVec_checkResult_lo_lo_4};
  wire [5:0]        checkVec_checkResult_hi_lo_4 = {checkVec_checkResultVec_5_4, checkVec_checkResultVec_4_4};
  wire [5:0]        checkVec_checkResult_hi_hi_4 = {checkVec_checkResultVec_7_4, checkVec_checkResultVec_6_4};
  wire [11:0]       checkVec_checkResult_hi_4 = {checkVec_checkResult_hi_hi_4, checkVec_checkResult_hi_lo_4};
  wire [23:0]       checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]        checkVec_checkResult_lo_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]        checkVec_checkResult_lo_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]        checkVec_checkResult_lo_5 = {checkVec_checkResult_lo_hi_5, checkVec_checkResult_lo_lo_5};
  wire [1:0]        checkVec_checkResult_hi_lo_5 = {checkVec_checkResultVec_5_5, checkVec_checkResultVec_4_5};
  wire [1:0]        checkVec_checkResult_hi_hi_5 = {checkVec_checkResultVec_7_5, checkVec_checkResultVec_6_5};
  wire [3:0]        checkVec_checkResult_hi_5 = {checkVec_checkResult_hi_hi_5, checkVec_checkResult_hi_lo_5};
  wire [7:0]        checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]        checkVec_checkResult_lo_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]        checkVec_checkResult_lo_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]        checkVec_checkResult_lo_6 = {checkVec_checkResult_lo_hi_6, checkVec_checkResult_lo_lo_6};
  wire [1:0]        checkVec_checkResult_hi_lo_6 = {checkVec_checkResultVec_5_6, checkVec_checkResultVec_4_6};
  wire [1:0]        checkVec_checkResult_hi_hi_6 = {checkVec_checkResultVec_7_6, checkVec_checkResultVec_6_6};
  wire [3:0]        checkVec_checkResult_hi_6 = {checkVec_checkResult_hi_hi_6, checkVec_checkResult_hi_lo_6};
  wire [7:0]        checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire              checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [9:0]        checkVec_checkResultVec_dataPosition_8 = {source_0[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_67 = 2'h1 << checkVec_checkResultVec_dataPosition_8[1];
  wire [3:0]        checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_67[1]}}, {2{_checkVec_checkResultVec_accessMask_T_67[0]}}};
  wire [1:0]        checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_8[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_8[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[9:5];
  wire [1:0]        checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_8[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[4:2];
  wire [2:0]        checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8[4:2];
  wire              checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_0[31:10]};
  wire              checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_0_6_1;
  wire              checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_9 = {source_1[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_75 = 2'h1 << checkVec_checkResultVec_dataPosition_9[1];
  wire [3:0]        checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_75[1]}}, {2{_checkVec_checkResultVec_accessMask_T_75[0]}}};
  wire [1:0]        checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_9[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_9[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[9:5];
  wire [1:0]        checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_9[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[4:2];
  wire [2:0]        checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9[4:2];
  wire              checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_1[31:10]};
  wire              checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_1_6_1;
  wire              checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_10 = {source_2[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_83 = 2'h1 << checkVec_checkResultVec_dataPosition_10[1];
  wire [3:0]        checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_83[1]}}, {2{_checkVec_checkResultVec_accessMask_T_83[0]}}};
  wire [1:0]        checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_10[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_10[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[9:5];
  wire [1:0]        checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_10[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[4:2];
  wire [2:0]        checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10[4:2];
  wire              checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_2[31:10]};
  wire              checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_2_6_1;
  wire              checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_11 = {source_3[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_91 = 2'h1 << checkVec_checkResultVec_dataPosition_11[1];
  wire [3:0]        checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_91[1]}}, {2{_checkVec_checkResultVec_accessMask_T_91[0]}}};
  wire [1:0]        checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_11[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_11[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[9:5];
  wire [1:0]        checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_11[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[4:2];
  wire [2:0]        checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11[4:2];
  wire              checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_3[31:10]};
  wire              checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_3_6_1;
  wire              checkVec_checkResultVec_4_6_1 = checkVec_validVec_1[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_12 = {source_4[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_99 = 2'h1 << checkVec_checkResultVec_dataPosition_12[1];
  wire [3:0]        checkVec_checkResultVec_4_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_99[1]}}, {2{_checkVec_checkResultVec_accessMask_T_99[0]}}};
  wire [1:0]        checkVec_checkResultVec_4_1_1 = {checkVec_checkResultVec_dataPosition_12[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_4_2_1 = checkVec_checkResultVec_dataPosition_12[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_12 = checkVec_checkResultVec_dataPosition_12[9:5];
  wire [1:0]        checkVec_checkResultVec_4_3_1 = checkVec_checkResultVec_dataGroup_12[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_12 = checkVec_checkResultVec_dataGroup_12[4:2];
  wire [2:0]        checkVec_checkResultVec_4_4_1 = checkVec_checkResultVec_accessRegGrowth_12;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_12 = {checkVec_checkResultVec_4_3_1, checkVec_checkResultVec_4_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_12 = checkVec_checkResultVec_decimalProportion_12[4:2];
  wire              checkVec_checkResultVec_overlap_12 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_12 >= checkVec_checkResultVec_intLMULInput_12[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_12} >= checkVec_checkResultVec_intLMULInput_12,
      source_4[31:10]};
  wire              checkVec_checkResultVec_4_5_1 = checkVec_checkResultVec_overlap_12 | ~checkVec_checkResultVec_4_6_1;
  wire              checkVec_checkResultVec_5_6_1 = checkVec_validVec_1[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_13 = {source_5[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_107 = 2'h1 << checkVec_checkResultVec_dataPosition_13[1];
  wire [3:0]        checkVec_checkResultVec_5_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_107[1]}}, {2{_checkVec_checkResultVec_accessMask_T_107[0]}}};
  wire [1:0]        checkVec_checkResultVec_5_1_1 = {checkVec_checkResultVec_dataPosition_13[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_5_2_1 = checkVec_checkResultVec_dataPosition_13[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_13 = checkVec_checkResultVec_dataPosition_13[9:5];
  wire [1:0]        checkVec_checkResultVec_5_3_1 = checkVec_checkResultVec_dataGroup_13[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_13 = checkVec_checkResultVec_dataGroup_13[4:2];
  wire [2:0]        checkVec_checkResultVec_5_4_1 = checkVec_checkResultVec_accessRegGrowth_13;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_13 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_5_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_13 = checkVec_checkResultVec_decimalProportion_13[4:2];
  wire              checkVec_checkResultVec_overlap_13 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_13 >= checkVec_checkResultVec_intLMULInput_13[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_13} >= checkVec_checkResultVec_intLMULInput_13,
      source_5[31:10]};
  wire              checkVec_checkResultVec_5_5_1 = checkVec_checkResultVec_overlap_13 | ~checkVec_checkResultVec_5_6_1;
  wire              checkVec_checkResultVec_6_6_1 = checkVec_validVec_1[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_14 = {source_6[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_115 = 2'h1 << checkVec_checkResultVec_dataPosition_14[1];
  wire [3:0]        checkVec_checkResultVec_6_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_115[1]}}, {2{_checkVec_checkResultVec_accessMask_T_115[0]}}};
  wire [1:0]        checkVec_checkResultVec_6_1_1 = {checkVec_checkResultVec_dataPosition_14[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_6_2_1 = checkVec_checkResultVec_dataPosition_14[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_14 = checkVec_checkResultVec_dataPosition_14[9:5];
  wire [1:0]        checkVec_checkResultVec_6_3_1 = checkVec_checkResultVec_dataGroup_14[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_14 = checkVec_checkResultVec_dataGroup_14[4:2];
  wire [2:0]        checkVec_checkResultVec_6_4_1 = checkVec_checkResultVec_accessRegGrowth_14;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_14 = {checkVec_checkResultVec_6_3_1, checkVec_checkResultVec_6_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_14 = checkVec_checkResultVec_decimalProportion_14[4:2];
  wire              checkVec_checkResultVec_overlap_14 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_14 >= checkVec_checkResultVec_intLMULInput_14[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_14} >= checkVec_checkResultVec_intLMULInput_14,
      source_6[31:10]};
  wire              checkVec_checkResultVec_6_5_1 = checkVec_checkResultVec_overlap_14 | ~checkVec_checkResultVec_6_6_1;
  wire              checkVec_checkResultVec_7_6_1 = checkVec_validVec_1[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_15 = {source_7[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_123 = 2'h1 << checkVec_checkResultVec_dataPosition_15[1];
  wire [3:0]        checkVec_checkResultVec_7_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_123[1]}}, {2{_checkVec_checkResultVec_accessMask_T_123[0]}}};
  wire [1:0]        checkVec_checkResultVec_7_1_1 = {checkVec_checkResultVec_dataPosition_15[1], 1'h0};
  wire [2:0]        checkVec_checkResultVec_7_2_1 = checkVec_checkResultVec_dataPosition_15[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_15 = checkVec_checkResultVec_dataPosition_15[9:5];
  wire [1:0]        checkVec_checkResultVec_7_3_1 = checkVec_checkResultVec_dataGroup_15[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_15 = checkVec_checkResultVec_dataGroup_15[4:2];
  wire [2:0]        checkVec_checkResultVec_7_4_1 = checkVec_checkResultVec_accessRegGrowth_15;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_15 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_7_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_15 = checkVec_checkResultVec_decimalProportion_15[4:2];
  wire              checkVec_checkResultVec_overlap_15 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_15 >= checkVec_checkResultVec_intLMULInput_15[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_15} >= checkVec_checkResultVec_intLMULInput_15,
      source_7[31:10]};
  wire              checkVec_checkResultVec_7_5_1 = checkVec_checkResultVec_overlap_15 | ~checkVec_checkResultVec_7_6_1;
  wire [7:0]        checkVec_checkResult_lo_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]        checkVec_checkResult_lo_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]       checkVec_checkResult_lo_7 = {checkVec_checkResult_lo_hi_7, checkVec_checkResult_lo_lo_7};
  wire [7:0]        checkVec_checkResult_hi_lo_7 = {checkVec_checkResultVec_5_0_1, checkVec_checkResultVec_4_0_1};
  wire [7:0]        checkVec_checkResult_hi_hi_7 = {checkVec_checkResultVec_7_0_1, checkVec_checkResultVec_6_0_1};
  wire [15:0]       checkVec_checkResult_hi_7 = {checkVec_checkResult_hi_hi_7, checkVec_checkResult_hi_lo_7};
  wire [31:0]       checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]        checkVec_checkResult_lo_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]        checkVec_checkResult_lo_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]        checkVec_checkResult_lo_8 = {checkVec_checkResult_lo_hi_8, checkVec_checkResult_lo_lo_8};
  wire [3:0]        checkVec_checkResult_hi_lo_8 = {checkVec_checkResultVec_5_1_1, checkVec_checkResultVec_4_1_1};
  wire [3:0]        checkVec_checkResult_hi_hi_8 = {checkVec_checkResultVec_7_1_1, checkVec_checkResultVec_6_1_1};
  wire [7:0]        checkVec_checkResult_hi_8 = {checkVec_checkResult_hi_hi_8, checkVec_checkResult_hi_lo_8};
  wire [15:0]       checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [5:0]        checkVec_checkResult_lo_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [5:0]        checkVec_checkResult_lo_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [11:0]       checkVec_checkResult_lo_9 = {checkVec_checkResult_lo_hi_9, checkVec_checkResult_lo_lo_9};
  wire [5:0]        checkVec_checkResult_hi_lo_9 = {checkVec_checkResultVec_5_2_1, checkVec_checkResultVec_4_2_1};
  wire [5:0]        checkVec_checkResult_hi_hi_9 = {checkVec_checkResultVec_7_2_1, checkVec_checkResultVec_6_2_1};
  wire [11:0]       checkVec_checkResult_hi_9 = {checkVec_checkResult_hi_hi_9, checkVec_checkResult_hi_lo_9};
  wire [23:0]       checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [3:0]        checkVec_checkResult_lo_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [3:0]        checkVec_checkResult_lo_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [7:0]        checkVec_checkResult_lo_10 = {checkVec_checkResult_lo_hi_10, checkVec_checkResult_lo_lo_10};
  wire [3:0]        checkVec_checkResult_hi_lo_10 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_4_3_1};
  wire [3:0]        checkVec_checkResult_hi_hi_10 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_6_3_1};
  wire [7:0]        checkVec_checkResult_hi_10 = {checkVec_checkResult_hi_hi_10, checkVec_checkResult_hi_lo_10};
  wire [15:0]       checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]        checkVec_checkResult_lo_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]        checkVec_checkResult_lo_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]       checkVec_checkResult_lo_11 = {checkVec_checkResult_lo_hi_11, checkVec_checkResult_lo_lo_11};
  wire [5:0]        checkVec_checkResult_hi_lo_11 = {checkVec_checkResultVec_5_4_1, checkVec_checkResultVec_4_4_1};
  wire [5:0]        checkVec_checkResult_hi_hi_11 = {checkVec_checkResultVec_7_4_1, checkVec_checkResultVec_6_4_1};
  wire [11:0]       checkVec_checkResult_hi_11 = {checkVec_checkResult_hi_hi_11, checkVec_checkResult_hi_lo_11};
  wire [23:0]       checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]        checkVec_checkResult_lo_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]        checkVec_checkResult_lo_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]        checkVec_checkResult_lo_12 = {checkVec_checkResult_lo_hi_12, checkVec_checkResult_lo_lo_12};
  wire [1:0]        checkVec_checkResult_hi_lo_12 = {checkVec_checkResultVec_5_5_1, checkVec_checkResultVec_4_5_1};
  wire [1:0]        checkVec_checkResult_hi_hi_12 = {checkVec_checkResultVec_7_5_1, checkVec_checkResultVec_6_5_1};
  wire [3:0]        checkVec_checkResult_hi_12 = {checkVec_checkResult_hi_hi_12, checkVec_checkResult_hi_lo_12};
  wire [7:0]        checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]        checkVec_checkResult_lo_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]        checkVec_checkResult_lo_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]        checkVec_checkResult_lo_13 = {checkVec_checkResult_lo_hi_13, checkVec_checkResult_lo_lo_13};
  wire [1:0]        checkVec_checkResult_hi_lo_13 = {checkVec_checkResultVec_5_6_1, checkVec_checkResultVec_4_6_1};
  wire [1:0]        checkVec_checkResult_hi_hi_13 = {checkVec_checkResultVec_7_6_1, checkVec_checkResultVec_6_6_1};
  wire [3:0]        checkVec_checkResult_hi_13 = {checkVec_checkResult_hi_hi_13, checkVec_checkResult_hi_lo_13};
  wire [7:0]        checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire              checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [9:0]        checkVec_checkResultVec_dataPosition_16 = {source_0[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_16[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_16 = checkVec_checkResultVec_dataPosition_16[9:5];
  wire [1:0]        checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_16[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_16 = checkVec_checkResultVec_dataGroup_16[4:2];
  wire [2:0]        checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_16;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_16 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_16 = checkVec_checkResultVec_decimalProportion_16[4:2];
  wire              checkVec_checkResultVec_overlap_16 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_16 >= checkVec_checkResultVec_intLMULInput_16[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_16} >= checkVec_checkResultVec_intLMULInput_16,
      source_0[31:10]};
  wire              checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_16 | ~checkVec_checkResultVec_0_6_2;
  wire              checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_17 = {source_1[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_17[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_17 = checkVec_checkResultVec_dataPosition_17[9:5];
  wire [1:0]        checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_17[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_17 = checkVec_checkResultVec_dataGroup_17[4:2];
  wire [2:0]        checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_17;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_17 = checkVec_checkResultVec_decimalProportion_17[4:2];
  wire              checkVec_checkResultVec_overlap_17 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_17 >= checkVec_checkResultVec_intLMULInput_17[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_17} >= checkVec_checkResultVec_intLMULInput_17,
      source_1[31:10]};
  wire              checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_17 | ~checkVec_checkResultVec_1_6_2;
  wire              checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_18 = {source_2[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_18[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_18 = checkVec_checkResultVec_dataPosition_18[9:5];
  wire [1:0]        checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_18[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_18 = checkVec_checkResultVec_dataGroup_18[4:2];
  wire [2:0]        checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_18;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_18 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_18 = checkVec_checkResultVec_decimalProportion_18[4:2];
  wire              checkVec_checkResultVec_overlap_18 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_18 >= checkVec_checkResultVec_intLMULInput_18[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_18} >= checkVec_checkResultVec_intLMULInput_18,
      source_2[31:10]};
  wire              checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_18 | ~checkVec_checkResultVec_2_6_2;
  wire              checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_19 = {source_3[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_19[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_19 = checkVec_checkResultVec_dataPosition_19[9:5];
  wire [1:0]        checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_19[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_19 = checkVec_checkResultVec_dataGroup_19[4:2];
  wire [2:0]        checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_19;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_19 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_19 = checkVec_checkResultVec_decimalProportion_19[4:2];
  wire              checkVec_checkResultVec_overlap_19 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_19 >= checkVec_checkResultVec_intLMULInput_19[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_19} >= checkVec_checkResultVec_intLMULInput_19,
      source_3[31:10]};
  wire              checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_19 | ~checkVec_checkResultVec_3_6_2;
  wire              checkVec_checkResultVec_4_6_2 = checkVec_validVec_2[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_20 = {source_4[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_4_2_2 = checkVec_checkResultVec_dataPosition_20[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_20 = checkVec_checkResultVec_dataPosition_20[9:5];
  wire [1:0]        checkVec_checkResultVec_4_3_2 = checkVec_checkResultVec_dataGroup_20[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_20 = checkVec_checkResultVec_dataGroup_20[4:2];
  wire [2:0]        checkVec_checkResultVec_4_4_2 = checkVec_checkResultVec_accessRegGrowth_20;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_20 = {checkVec_checkResultVec_4_3_2, checkVec_checkResultVec_4_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_20 = checkVec_checkResultVec_decimalProportion_20[4:2];
  wire              checkVec_checkResultVec_overlap_20 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_20 >= checkVec_checkResultVec_intLMULInput_20[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_20} >= checkVec_checkResultVec_intLMULInput_20,
      source_4[31:10]};
  wire              checkVec_checkResultVec_4_5_2 = checkVec_checkResultVec_overlap_20 | ~checkVec_checkResultVec_4_6_2;
  wire              checkVec_checkResultVec_5_6_2 = checkVec_validVec_2[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_21 = {source_5[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_5_2_2 = checkVec_checkResultVec_dataPosition_21[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_21 = checkVec_checkResultVec_dataPosition_21[9:5];
  wire [1:0]        checkVec_checkResultVec_5_3_2 = checkVec_checkResultVec_dataGroup_21[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_21 = checkVec_checkResultVec_dataGroup_21[4:2];
  wire [2:0]        checkVec_checkResultVec_5_4_2 = checkVec_checkResultVec_accessRegGrowth_21;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_21 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_5_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_21 = checkVec_checkResultVec_decimalProportion_21[4:2];
  wire              checkVec_checkResultVec_overlap_21 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_21 >= checkVec_checkResultVec_intLMULInput_21[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_21} >= checkVec_checkResultVec_intLMULInput_21,
      source_5[31:10]};
  wire              checkVec_checkResultVec_5_5_2 = checkVec_checkResultVec_overlap_21 | ~checkVec_checkResultVec_5_6_2;
  wire              checkVec_checkResultVec_6_6_2 = checkVec_validVec_2[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_22 = {source_6[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_6_2_2 = checkVec_checkResultVec_dataPosition_22[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_22 = checkVec_checkResultVec_dataPosition_22[9:5];
  wire [1:0]        checkVec_checkResultVec_6_3_2 = checkVec_checkResultVec_dataGroup_22[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_22 = checkVec_checkResultVec_dataGroup_22[4:2];
  wire [2:0]        checkVec_checkResultVec_6_4_2 = checkVec_checkResultVec_accessRegGrowth_22;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_22 = {checkVec_checkResultVec_6_3_2, checkVec_checkResultVec_6_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_22 = checkVec_checkResultVec_decimalProportion_22[4:2];
  wire              checkVec_checkResultVec_overlap_22 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_22 >= checkVec_checkResultVec_intLMULInput_22[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_22} >= checkVec_checkResultVec_intLMULInput_22,
      source_6[31:10]};
  wire              checkVec_checkResultVec_6_5_2 = checkVec_checkResultVec_overlap_22 | ~checkVec_checkResultVec_6_6_2;
  wire              checkVec_checkResultVec_7_6_2 = checkVec_validVec_2[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_23 = {source_7[7:0], 2'h0};
  wire [2:0]        checkVec_checkResultVec_7_2_2 = checkVec_checkResultVec_dataPosition_23[4:2];
  wire [4:0]        checkVec_checkResultVec_dataGroup_23 = checkVec_checkResultVec_dataPosition_23[9:5];
  wire [1:0]        checkVec_checkResultVec_7_3_2 = checkVec_checkResultVec_dataGroup_23[1:0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_23 = checkVec_checkResultVec_dataGroup_23[4:2];
  wire [2:0]        checkVec_checkResultVec_7_4_2 = checkVec_checkResultVec_accessRegGrowth_23;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_23 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_7_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_23 = checkVec_checkResultVec_decimalProportion_23[4:2];
  wire              checkVec_checkResultVec_overlap_23 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_23 >= checkVec_checkResultVec_intLMULInput_23[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_23} >= checkVec_checkResultVec_intLMULInput_23,
      source_7[31:10]};
  wire              checkVec_checkResultVec_7_5_2 = checkVec_checkResultVec_overlap_23 | ~checkVec_checkResultVec_7_6_2;
  wire [5:0]        checkVec_checkResult_lo_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [5:0]        checkVec_checkResult_lo_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [11:0]       checkVec_checkResult_lo_16 = {checkVec_checkResult_lo_hi_16, checkVec_checkResult_lo_lo_16};
  wire [5:0]        checkVec_checkResult_hi_lo_16 = {checkVec_checkResultVec_5_2_2, checkVec_checkResultVec_4_2_2};
  wire [5:0]        checkVec_checkResult_hi_hi_16 = {checkVec_checkResultVec_7_2_2, checkVec_checkResultVec_6_2_2};
  wire [11:0]       checkVec_checkResult_hi_16 = {checkVec_checkResult_hi_hi_16, checkVec_checkResult_hi_lo_16};
  wire [23:0]       checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [3:0]        checkVec_checkResult_lo_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [3:0]        checkVec_checkResult_lo_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [7:0]        checkVec_checkResult_lo_17 = {checkVec_checkResult_lo_hi_17, checkVec_checkResult_lo_lo_17};
  wire [3:0]        checkVec_checkResult_hi_lo_17 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_4_3_2};
  wire [3:0]        checkVec_checkResult_hi_hi_17 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_6_3_2};
  wire [7:0]        checkVec_checkResult_hi_17 = {checkVec_checkResult_hi_hi_17, checkVec_checkResult_hi_lo_17};
  wire [15:0]       checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]        checkVec_checkResult_lo_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]        checkVec_checkResult_lo_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]       checkVec_checkResult_lo_18 = {checkVec_checkResult_lo_hi_18, checkVec_checkResult_lo_lo_18};
  wire [5:0]        checkVec_checkResult_hi_lo_18 = {checkVec_checkResultVec_5_4_2, checkVec_checkResultVec_4_4_2};
  wire [5:0]        checkVec_checkResult_hi_hi_18 = {checkVec_checkResultVec_7_4_2, checkVec_checkResultVec_6_4_2};
  wire [11:0]       checkVec_checkResult_hi_18 = {checkVec_checkResult_hi_hi_18, checkVec_checkResult_hi_lo_18};
  wire [23:0]       checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]        checkVec_checkResult_lo_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]        checkVec_checkResult_lo_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]        checkVec_checkResult_lo_19 = {checkVec_checkResult_lo_hi_19, checkVec_checkResult_lo_lo_19};
  wire [1:0]        checkVec_checkResult_hi_lo_19 = {checkVec_checkResultVec_5_5_2, checkVec_checkResultVec_4_5_2};
  wire [1:0]        checkVec_checkResult_hi_hi_19 = {checkVec_checkResultVec_7_5_2, checkVec_checkResultVec_6_5_2};
  wire [3:0]        checkVec_checkResult_hi_19 = {checkVec_checkResult_hi_hi_19, checkVec_checkResult_hi_lo_19};
  wire [7:0]        checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]        checkVec_checkResult_lo_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]        checkVec_checkResult_lo_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]        checkVec_checkResult_lo_20 = {checkVec_checkResult_lo_hi_20, checkVec_checkResult_lo_lo_20};
  wire [1:0]        checkVec_checkResult_hi_lo_20 = {checkVec_checkResultVec_5_6_2, checkVec_checkResultVec_4_6_2};
  wire [1:0]        checkVec_checkResult_hi_hi_20 = {checkVec_checkResultVec_7_6_2, checkVec_checkResultVec_6_6_2};
  wire [3:0]        checkVec_checkResult_hi_20 = {checkVec_checkResult_hi_hi_20, checkVec_checkResult_hi_lo_20};
  wire [7:0]        checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [15:0]       dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 16'h0) | (sew1H[1] ? checkVec_1_1 : 16'h0);
  wire [23:0]       accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 24'h0) | (sew1H[1] ? checkVec_1_2 : 24'h0) | (sew1H[2] ? checkVec_2_2 : 24'h0);
  wire [15:0]       offsetSelect = (sew1H[0] ? checkVec_0_3 : 16'h0) | (sew1H[1] ? checkVec_1_3 : 16'h0) | (sew1H[2] ? checkVec_2_3 : 16'h0);
  wire [23:0]       growthSelect = (sew1H[0] ? checkVec_0_4 : 24'h0) | (sew1H[1] ? checkVec_1_4 : 24'h0) | (sew1H[2] ? checkVec_2_4 : 24'h0);
  wire [7:0]        notReadSelect = (sew1H[0] ? checkVec_0_5 : 8'h0) | (sew1H[1] ? checkVec_1_5 : 8'h0) | (sew1H[2] ? checkVec_2_5 : 8'h0);
  wire [7:0]        elementValidSelect = (sew1H[0] ? checkVec_0_6 : 8'h0) | (sew1H[1] ? checkVec_1_6 : 8'h0) | (sew1H[2] ? checkVec_2_6 : 8'h0);
  wire              readTypeRequestDeq;
  wire              waiteStageEnqReady;
  wire              readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [7:0]        readWaitQueue_dataOut_executeGroup;
  wire [7:0]        readWaitQueue_dataOut_sourceValid;
  wire [7:0]        readWaitQueue_dataOut_replaceVs1;
  wire [7:0]        readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_dataOut_last;
  wire [8:0]        readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [15:0]       readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [23:0]       readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [32:0]       readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[8:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[16:9];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[24:17];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[32:25];
  wire [7:0]        readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [7:0]        readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [7:0]        readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [7:0]        readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire              readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire              readWaitQueue_enq_valid;
  wire              readWaitQueue_deq_ready;
  wire              _GEN_70 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_70;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_70;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_70;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_70;
  assign exeRequestQueue_4_deq_ready = ~exeReqReg_4_valid | _GEN_70;
  assign exeRequestQueue_5_deq_ready = ~exeReqReg_5_valid | _GEN_70;
  assign exeRequestQueue_6_deq_ready = ~exeReqReg_6_valid | _GEN_70;
  assign exeRequestQueue_7_deq_ready = ~exeReqReg_7_valid | _GEN_70;
  wire              isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire              allDataValid =
    (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3])) & (exeReqReg_4_valid | ~(groupDataNeed[4]))
    & (exeReqReg_5_valid | ~(groupDataNeed[5])) & (exeReqReg_6_valid | ~(groupDataNeed[6])) & (exeReqReg_7_valid | ~(groupDataNeed[7]));
  wire              anyDataValid = exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid | exeReqReg_4_valid | exeReqReg_5_valid | exeReqReg_6_valid | exeReqReg_7_valid;
  wire              _GEN_71 = compress | mvRd;
  wire              readVs1Valid = (unitType[2] | _GEN_71) & ~readVS1Reg_requestSend | gatherSRead;
  wire              _GEN_72 = compress | ~gatherSRead;
  wire [4:0]        readVS1Req_vs = _GEN_72 ? instReg_vs1 : instReg_vs1 + {2'h0, gatherGrowth};
  wire [1:0]        readVS1Req_offset = compress ? readVS1Reg_readIndex[4:3] : gatherSRead ? gatherOffset : 2'h0;
  wire [2:0]        readVS1Req_readLane = compress ? readVS1Reg_readIndex[2:0] : gatherSRead ? gatherLane : 3'h0;
  wire [1:0]        readVS1Req_dataOffset = _GEN_72 ? 2'h0 : gatherDatOffset;
  wire [1:0]        selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[3:2];
  wire [1:0]        selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[5:4];
  wire [1:0]        selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[7:6];
  wire [1:0]        selectExecuteReq_4_bits_offset = readIssueStageState_readOffset[9:8];
  wire [1:0]        selectExecuteReq_5_bits_offset = readIssueStageState_readOffset[11:10];
  wire [1:0]        selectExecuteReq_6_bits_offset = readIssueStageState_readOffset[13:12];
  wire [1:0]        selectExecuteReq_7_bits_offset = readIssueStageState_readOffset[15:14];
  wire [1:0]        selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]        selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]        selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire [1:0]        selectExecuteReq_4_bits_dataOffset = readIssueStageState_readDataOffset[9:8];
  wire [1:0]        selectExecuteReq_5_bits_dataOffset = readIssueStageState_readDataOffset[11:10];
  wire [1:0]        selectExecuteReq_6_bits_dataOffset = readIssueStageState_readDataOffset[13:12];
  wire [1:0]        selectExecuteReq_7_bits_dataOffset = readIssueStageState_readDataOffset[15:14];
  wire              selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]        selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire [1:0]        selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[1:0];
  wire [2:0]        selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]        selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire              _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire              pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]        selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire              selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire              pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]        selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire              selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire              pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]        selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire              selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire              pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  wire [4:0]        selectExecuteReq_4_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_4};
  wire              selectExecuteReq_4_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[4]) & readIssueStageState_needRead[4] & readType;
  wire              pipeReadFire_4 = _readCrossBar_input_4_ready & readCrossBar_input_4_valid;
  wire [4:0]        selectExecuteReq_5_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_5};
  wire              selectExecuteReq_5_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[5]) & readIssueStageState_needRead[5] & readType;
  wire              pipeReadFire_5 = _readCrossBar_input_5_ready & readCrossBar_input_5_valid;
  wire [4:0]        selectExecuteReq_6_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_6};
  wire              selectExecuteReq_6_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[6]) & readIssueStageState_needRead[6] & readType;
  wire              pipeReadFire_6 = _readCrossBar_input_6_ready & readCrossBar_input_6_valid;
  wire [4:0]        selectExecuteReq_7_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_7};
  wire              selectExecuteReq_7_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[7]) & readIssueStageState_needRead[7] & readType;
  wire              pipeReadFire_7 = _readCrossBar_input_7_ready & readCrossBar_input_7_valid;
  reg  [3:0]        tokenCheck_counter;
  wire [3:0]        tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire              tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]        tokenCheck_counter_1;
  wire [3:0]        tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire              tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]        tokenCheck_counter_2;
  wire [3:0]        tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire              tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]        tokenCheck_counter_3;
  wire [3:0]        tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire              tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  reg  [3:0]        tokenCheck_counter_4;
  wire [3:0]        tokenCheck_counterChange_4 = pipeReadFire_4 ? 4'h1 : 4'hF;
  wire              tokenCheck_4 = ~(tokenCheck_counter_4[3]);
  assign readCrossBar_input_4_valid = selectExecuteReq_4_valid & tokenCheck_4;
  reg  [3:0]        tokenCheck_counter_5;
  wire [3:0]        tokenCheck_counterChange_5 = pipeReadFire_5 ? 4'h1 : 4'hF;
  wire              tokenCheck_5 = ~(tokenCheck_counter_5[3]);
  assign readCrossBar_input_5_valid = selectExecuteReq_5_valid & tokenCheck_5;
  reg  [3:0]        tokenCheck_counter_6;
  wire [3:0]        tokenCheck_counterChange_6 = pipeReadFire_6 ? 4'h1 : 4'hF;
  wire              tokenCheck_6 = ~(tokenCheck_counter_6[3]);
  assign readCrossBar_input_6_valid = selectExecuteReq_6_valid & tokenCheck_6;
  reg  [3:0]        tokenCheck_counter_7;
  wire [3:0]        tokenCheck_counterChange_7 = pipeReadFire_7 ? 4'h1 : 4'hF;
  wire              tokenCheck_7 = ~(tokenCheck_counter_7[3]);
  assign readCrossBar_input_7_valid = selectExecuteReq_7_valid & tokenCheck_7;
  wire [1:0]        readFire_lo_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]        readFire_lo_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]        readFire_lo = {readFire_lo_hi, readFire_lo_lo};
  wire [1:0]        readFire_hi_lo = {pipeReadFire_5, pipeReadFire_4};
  wire [1:0]        readFire_hi_hi = {pipeReadFire_7, pipeReadFire_6};
  wire [3:0]        readFire_hi = {readFire_hi_hi, readFire_hi_lo};
  wire [7:0]        readFire = {readFire_hi, readFire_lo};
  wire              anyReadFire = |readFire;
  wire [7:0]        readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire              groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 8'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [7:0]        compressUnitResultQueue_enq_bits_ffoOutput;
  wire              compressUnitResultQueue_enq_bits_compressValid;
  wire [8:0]        compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [255:0]      compressUnitResultQueue_enq_bits_data;
  wire [31:0]       compressUnitResultQueue_enq_bits_mask;
  wire [287:0]      compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [5:0]        compressUnitResultQueue_enq_bits_groupCounter;
  wire [293:0]      compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [302:0]      compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire              compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [7:0]        compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[8:1];
  wire [5:0]        compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[14:9];
  wire [31:0]       compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[46:15];
  wire [255:0]      compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[302:47];
  wire              compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire              compressUnitResultQueue_deq_ready;
  wire              compressUnitResultQueue_enq_valid;
  wire              compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [255:0]      compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [31:0]       compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [5:0]        compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [7:0]        compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire              compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire              noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire              vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_71);
  wire [1:0]        _GEN_73 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]        executeDeqReady_lo_lo;
  assign executeDeqReady_lo_lo = _GEN_73;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_lo;
  assign compressUnitResultQueue_deq_ready_lo_lo = _GEN_73;
  wire [1:0]        _GEN_74 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]        executeDeqReady_lo_hi;
  assign executeDeqReady_lo_hi = _GEN_74;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_hi;
  assign compressUnitResultQueue_deq_ready_lo_hi = _GEN_74;
  wire [3:0]        executeDeqReady_lo = {executeDeqReady_lo_hi, executeDeqReady_lo_lo};
  wire [1:0]        _GEN_75 = {_maskedWrite_in_5_ready, _maskedWrite_in_4_ready};
  wire [1:0]        executeDeqReady_hi_lo;
  assign executeDeqReady_hi_lo = _GEN_75;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_lo;
  assign compressUnitResultQueue_deq_ready_hi_lo = _GEN_75;
  wire [1:0]        _GEN_76 = {_maskedWrite_in_7_ready, _maskedWrite_in_6_ready};
  wire [1:0]        executeDeqReady_hi_hi;
  assign executeDeqReady_hi_hi = _GEN_76;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_hi;
  assign compressUnitResultQueue_deq_ready_hi_hi = _GEN_76;
  wire [3:0]        executeDeqReady_hi = {executeDeqReady_hi_hi, executeDeqReady_hi_lo};
  wire              compressUnitResultQueue_empty;
  wire              executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire              otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire              reorderQueueAllocate;
  wire              _GEN_77 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_77;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire              executeReady;
  wire              requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire              slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_77;
  wire              _GEN_78 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire              _GEN_79 = readIssueStageEnq & _GEN_78;
  assign accessCountEnq_0 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h0 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h0 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h0 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h0 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h0 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h0 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h0 & ~(notReadSelect[7])}}};
  assign accessCountEnq_1 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h1 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h1 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h1 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h1 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h1 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h1 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h1 & ~(notReadSelect[7])}}};
  assign accessCountEnq_2 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h2 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h2 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h2 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h2 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h2 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h2 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h2 & ~(notReadSelect[7])}}};
  assign accessCountEnq_3 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h3 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h3 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h3 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h3 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h3 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h3 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h3 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h3 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h3 & ~(notReadSelect[7])}}};
  assign accessCountEnq_4 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h4 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h4 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h4 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h4 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h4 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h4 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h4 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h4 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h4 & ~(notReadSelect[7])}}};
  assign accessCountEnq_5 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h5 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h5 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h5 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h5 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h5 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h5 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h5 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h5 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h5 & ~(notReadSelect[7])}}};
  assign accessCountEnq_6 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 3'h6 & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, accessLaneSelect[2:0] == 3'h6 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[5:3] == 3'h6 & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, accessLaneSelect[8:6] == 3'h6 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[11:9] == 3'h6 & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, accessLaneSelect[14:12] == 3'h6 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[17:15] == 3'h6 & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, accessLaneSelect[20:18] == 3'h6 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[23:21] == 3'h6 & ~(notReadSelect[7])}}};
  assign accessCountEnq_7 =
    _GEN_79
      ? {1'h0,
         {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
           + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}}
        + {1'h0,
           {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_4) & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_5) & _slideAddressGen_indexDeq_bits_needRead[5]}}
             + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_6) & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_7) & _slideAddressGen_indexDeq_bits_needRead[7]}}}
      : {1'h0,
         {1'h0, {1'h0, (&(accessLaneSelect[2:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[5:3])) & ~(notReadSelect[1])}}
           + {1'h0, {1'h0, (&(accessLaneSelect[8:6])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[11:9])) & ~(notReadSelect[3])}}}
        + {1'h0,
           {1'h0, {1'h0, (&(accessLaneSelect[14:12])) & ~(notReadSelect[4])} + {1'h0, (&(accessLaneSelect[17:15])) & ~(notReadSelect[5])}}
             + {1'h0, {1'h0, (&(accessLaneSelect[20:18])) & ~(notReadSelect[6])} + {1'h0, (&(accessLaneSelect[23:21])) & ~(notReadSelect[7])}}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [7:0]        readMessageQueue_deq_bits_readSource;
  wire              deqAllocate;
  wire              reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]       reorderQueueVec_dataOut_data;
  wire [7:0]        reorderQueueVec_dataOut_write1H;
  wire [31:0]       dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_enq_bits_data;
  wire [7:0]        reorderQueueVec_0_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[7:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[39:8];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [7:0]        reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire              reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire              reorderQueueVec_0_deq_ready;
  wire [7:0]        readMessageQueue_1_deq_bits_readSource;
  wire              deqAllocate_1;
  wire              reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]       reorderQueueVec_dataOut_1_data;
  wire [7:0]        reorderQueueVec_dataOut_1_write1H;
  wire [31:0]       dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_enq_bits_data;
  wire [7:0]        reorderQueueVec_1_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[7:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[39:8];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [7:0]        reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire              reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_1_deq_ready;
  wire [7:0]        readMessageQueue_2_deq_bits_readSource;
  wire              deqAllocate_2;
  wire              reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]       reorderQueueVec_dataOut_2_data;
  wire [7:0]        reorderQueueVec_dataOut_2_write1H;
  wire [31:0]       dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_enq_bits_data;
  wire [7:0]        reorderQueueVec_2_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[7:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[39:8];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [7:0]        reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire              reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_2_deq_ready;
  wire [7:0]        readMessageQueue_3_deq_bits_readSource;
  wire              deqAllocate_3;
  wire              reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]       reorderQueueVec_dataOut_3_data;
  wire [7:0]        reorderQueueVec_dataOut_3_write1H;
  wire [31:0]       dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_3_enq_bits_data;
  wire [7:0]        reorderQueueVec_3_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[7:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[39:8];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [7:0]        reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire              reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire              reorderQueueVec_3_deq_ready;
  wire [7:0]        readMessageQueue_4_deq_bits_readSource;
  wire              deqAllocate_4;
  wire              reorderQueueVec_4_deq_valid;
  assign reorderQueueVec_4_deq_valid = ~_reorderQueueVec_fifo_4_empty;
  wire [31:0]       reorderQueueVec_dataOut_4_data;
  wire [7:0]        reorderQueueVec_dataOut_4_write1H;
  wire [31:0]       dataAfterReorderCheck_4 = reorderQueueVec_4_deq_bits_data;
  wire [31:0]       reorderQueueVec_4_enq_bits_data;
  wire [7:0]        reorderQueueVec_4_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_4 = {reorderQueueVec_4_enq_bits_data, reorderQueueVec_4_enq_bits_write1H};
  assign reorderQueueVec_dataOut_4_write1H = _reorderQueueVec_fifo_4_data_out[7:0];
  assign reorderQueueVec_dataOut_4_data = _reorderQueueVec_fifo_4_data_out[39:8];
  assign reorderQueueVec_4_deq_bits_data = reorderQueueVec_dataOut_4_data;
  wire [7:0]        reorderQueueVec_4_deq_bits_write1H = reorderQueueVec_dataOut_4_write1H;
  wire              reorderQueueVec_4_enq_ready = ~_reorderQueueVec_fifo_4_full;
  wire              reorderQueueVec_4_deq_ready;
  wire [7:0]        readMessageQueue_5_deq_bits_readSource;
  wire              deqAllocate_5;
  wire              reorderQueueVec_5_deq_valid;
  assign reorderQueueVec_5_deq_valid = ~_reorderQueueVec_fifo_5_empty;
  wire [31:0]       reorderQueueVec_dataOut_5_data;
  wire [7:0]        reorderQueueVec_dataOut_5_write1H;
  wire [31:0]       dataAfterReorderCheck_5 = reorderQueueVec_5_deq_bits_data;
  wire [31:0]       reorderQueueVec_5_enq_bits_data;
  wire [7:0]        reorderQueueVec_5_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_5 = {reorderQueueVec_5_enq_bits_data, reorderQueueVec_5_enq_bits_write1H};
  assign reorderQueueVec_dataOut_5_write1H = _reorderQueueVec_fifo_5_data_out[7:0];
  assign reorderQueueVec_dataOut_5_data = _reorderQueueVec_fifo_5_data_out[39:8];
  assign reorderQueueVec_5_deq_bits_data = reorderQueueVec_dataOut_5_data;
  wire [7:0]        reorderQueueVec_5_deq_bits_write1H = reorderQueueVec_dataOut_5_write1H;
  wire              reorderQueueVec_5_enq_ready = ~_reorderQueueVec_fifo_5_full;
  wire              reorderQueueVec_5_deq_ready;
  wire [7:0]        readMessageQueue_6_deq_bits_readSource;
  wire              deqAllocate_6;
  wire              reorderQueueVec_6_deq_valid;
  assign reorderQueueVec_6_deq_valid = ~_reorderQueueVec_fifo_6_empty;
  wire [31:0]       reorderQueueVec_dataOut_6_data;
  wire [7:0]        reorderQueueVec_dataOut_6_write1H;
  wire [31:0]       dataAfterReorderCheck_6 = reorderQueueVec_6_deq_bits_data;
  wire [31:0]       reorderQueueVec_6_enq_bits_data;
  wire [7:0]        reorderQueueVec_6_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_6 = {reorderQueueVec_6_enq_bits_data, reorderQueueVec_6_enq_bits_write1H};
  assign reorderQueueVec_dataOut_6_write1H = _reorderQueueVec_fifo_6_data_out[7:0];
  assign reorderQueueVec_dataOut_6_data = _reorderQueueVec_fifo_6_data_out[39:8];
  assign reorderQueueVec_6_deq_bits_data = reorderQueueVec_dataOut_6_data;
  wire [7:0]        reorderQueueVec_6_deq_bits_write1H = reorderQueueVec_dataOut_6_write1H;
  wire              reorderQueueVec_6_enq_ready = ~_reorderQueueVec_fifo_6_full;
  wire              reorderQueueVec_6_deq_ready;
  wire [7:0]        readMessageQueue_7_deq_bits_readSource;
  wire              deqAllocate_7;
  wire              reorderQueueVec_7_deq_valid;
  assign reorderQueueVec_7_deq_valid = ~_reorderQueueVec_fifo_7_empty;
  wire [31:0]       reorderQueueVec_dataOut_7_data;
  wire [7:0]        reorderQueueVec_dataOut_7_write1H;
  wire [31:0]       dataAfterReorderCheck_7 = reorderQueueVec_7_deq_bits_data;
  wire [31:0]       reorderQueueVec_7_enq_bits_data;
  wire [7:0]        reorderQueueVec_7_enq_bits_write1H;
  wire [39:0]       reorderQueueVec_dataIn_7 = {reorderQueueVec_7_enq_bits_data, reorderQueueVec_7_enq_bits_write1H};
  assign reorderQueueVec_dataOut_7_write1H = _reorderQueueVec_fifo_7_data_out[7:0];
  assign reorderQueueVec_dataOut_7_data = _reorderQueueVec_fifo_7_data_out[39:8];
  assign reorderQueueVec_7_deq_bits_data = reorderQueueVec_dataOut_7_data;
  wire [7:0]        reorderQueueVec_7_deq_bits_write1H = reorderQueueVec_dataOut_7_write1H;
  wire              reorderQueueVec_7_enq_ready = ~_reorderQueueVec_fifo_7_full;
  wire              reorderQueueVec_7_deq_ready;
  reg  [4:0]        reorderQueueAllocate_counter;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate;
  wire              _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire              reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {4'h0, reorderQueueAllocate_release};
  reg  [4:0]        reorderQueueAllocate_counter_1;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_1;
  wire              _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire              reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {4'h0, reorderQueueAllocate_release_1};
  reg  [4:0]        reorderQueueAllocate_counter_2;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_2;
  wire              _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire              reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {4'h0, reorderQueueAllocate_release_2};
  reg  [4:0]        reorderQueueAllocate_counter_3;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_3;
  wire              _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire              reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {4'h0, reorderQueueAllocate_release_3};
  reg  [4:0]        reorderQueueAllocate_counter_4;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_4;
  wire              _write1HPipe_4_T = reorderQueueVec_4_deq_ready & reorderQueueVec_4_deq_valid;
  wire              reorderQueueAllocate_release_4 = _write1HPipe_4_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_4 = readIssueStageEnq ? accessCountEnq_4 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_4 = reorderQueueAllocate_counter_4 + {1'h0, reorderQueueAllocate_allocate_4} - {4'h0, reorderQueueAllocate_release_4};
  reg  [4:0]        reorderQueueAllocate_counter_5;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_5;
  wire              _write1HPipe_5_T = reorderQueueVec_5_deq_ready & reorderQueueVec_5_deq_valid;
  wire              reorderQueueAllocate_release_5 = _write1HPipe_5_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_5 = readIssueStageEnq ? accessCountEnq_5 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_5 = reorderQueueAllocate_counter_5 + {1'h0, reorderQueueAllocate_allocate_5} - {4'h0, reorderQueueAllocate_release_5};
  reg  [4:0]        reorderQueueAllocate_counter_6;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_6;
  wire              _write1HPipe_6_T = reorderQueueVec_6_deq_ready & reorderQueueVec_6_deq_valid;
  wire              reorderQueueAllocate_release_6 = _write1HPipe_6_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_6 = readIssueStageEnq ? accessCountEnq_6 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_6 = reorderQueueAllocate_counter_6 + {1'h0, reorderQueueAllocate_allocate_6} - {4'h0, reorderQueueAllocate_release_6};
  reg  [4:0]        reorderQueueAllocate_counter_7;
  reg  [4:0]        reorderQueueAllocate_counterWillUpdate_7;
  wire              _write1HPipe_7_T = reorderQueueVec_7_deq_ready & reorderQueueVec_7_deq_valid;
  wire              reorderQueueAllocate_release_7 = _write1HPipe_7_T & readValid;
  wire [3:0]        reorderQueueAllocate_allocate_7 = readIssueStageEnq ? accessCountEnq_7 : 4'h0;
  wire [4:0]        reorderQueueAllocate_counterUpdate_7 = reorderQueueAllocate_counter_7 + {1'h0, reorderQueueAllocate_allocate_7} - {4'h0, reorderQueueAllocate_release_7};
  assign reorderQueueAllocate =
    ~(reorderQueueAllocate_counterWillUpdate[4]) & ~(reorderQueueAllocate_counterWillUpdate_1[4]) & ~(reorderQueueAllocate_counterWillUpdate_2[4]) & ~(reorderQueueAllocate_counterWillUpdate_3[4])
    & ~(reorderQueueAllocate_counterWillUpdate_4[4]) & ~(reorderQueueAllocate_counterWillUpdate_5[4]) & ~(reorderQueueAllocate_counterWillUpdate_6[4]) & ~(reorderQueueAllocate_counterWillUpdate_7[4]);
  reg               reorderStageValid;
  reg  [3:0]        reorderStageState_0;
  reg  [3:0]        reorderStageState_1;
  reg  [3:0]        reorderStageState_2;
  reg  [3:0]        reorderStageState_3;
  reg  [3:0]        reorderStageState_4;
  reg  [3:0]        reorderStageState_5;
  reg  [3:0]        reorderStageState_6;
  reg  [3:0]        reorderStageState_7;
  reg  [3:0]        reorderStageNeed_0;
  reg  [3:0]        reorderStageNeed_1;
  reg  [3:0]        reorderStageNeed_2;
  reg  [3:0]        reorderStageNeed_3;
  reg  [3:0]        reorderStageNeed_4;
  reg  [3:0]        reorderStageNeed_5;
  reg  [3:0]        reorderStageNeed_6;
  reg  [3:0]        reorderStageNeed_7;
  wire              stateCheck =
    reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3 & reorderStageState_4 == reorderStageNeed_4
    & reorderStageState_5 == reorderStageNeed_5 & reorderStageState_6 == reorderStageNeed_6 & reorderStageState_7 == reorderStageNeed_7;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire              reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire              reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [7:0]        sourceLane;
  wire              readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [7:0]        readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_dataOffset;
  wire [7:0]        readMessageQueue_enq_bits_readSource;
  wire [1:0]        readMessageQueue_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[9:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]        readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire              readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire              readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 8'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire              readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]        readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire [1:0]        readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_1;
  wire              readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [7:0]        readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_1_dataOffset;
  wire [7:0]        readMessageQueue_1_enq_bits_readSource;
  wire [1:0]        readMessageQueue_1_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[9:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]        readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire              readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire              readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 8'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire              readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]        readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire [1:0]        readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_2;
  wire              readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [7:0]        readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_2_dataOffset;
  wire [7:0]        readMessageQueue_2_enq_bits_readSource;
  wire [1:0]        readMessageQueue_2_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[9:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]        readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire              readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire              readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 8'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire              readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]        readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire [1:0]        readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_3;
  wire              readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [7:0]        readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_3_dataOffset;
  wire [7:0]        readMessageQueue_3_enq_bits_readSource;
  wire [1:0]        readMessageQueue_3_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[9:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]        readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire              readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire              readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 8'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire              readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]        readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire [1:0]        readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_4;
  wire              readMessageQueue_4_deq_valid;
  assign readMessageQueue_4_deq_valid = ~_readMessageQueue_fifo_4_empty;
  wire [7:0]        readMessageQueue_dataOut_4_readSource;
  assign reorderQueueVec_4_enq_bits_write1H = readMessageQueue_4_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_4_dataOffset;
  wire [7:0]        readMessageQueue_4_enq_bits_readSource;
  wire [1:0]        readMessageQueue_4_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_4 = {readMessageQueue_4_enq_bits_readSource, readMessageQueue_4_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_4_dataOffset = _readMessageQueue_fifo_4_data_out[1:0];
  assign readMessageQueue_dataOut_4_readSource = _readMessageQueue_fifo_4_data_out[9:2];
  assign readMessageQueue_4_deq_bits_readSource = readMessageQueue_dataOut_4_readSource;
  wire [1:0]        readMessageQueue_4_deq_bits_dataOffset = readMessageQueue_dataOut_4_dataOffset;
  wire              readMessageQueue_4_enq_ready = ~_readMessageQueue_fifo_4_full;
  wire              readMessageQueue_4_enq_valid;
  assign deqAllocate_4 = ~readValid | reorderStageValid & reorderStageState_4 != reorderStageNeed_4;
  assign reorderQueueVec_4_deq_ready = deqAllocate_4;
  assign sourceLane_4 = 8'h1 << _readCrossBar_output_4_bits_writeIndex;
  assign readMessageQueue_4_enq_bits_readSource = sourceLane_4;
  wire              readChannel_4_valid_0 = maskDestinationType ? _maskedWrite_readChannel_4_valid : _readCrossBar_output_4_valid & readMessageQueue_4_enq_ready;
  wire [4:0]        readChannel_4_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_vs : _readCrossBar_output_4_bits_vs;
  wire [1:0]        readChannel_4_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_offset : _readCrossBar_output_4_bits_offset;
  assign readMessageQueue_4_enq_valid = readChannel_4_ready_0 & readChannel_4_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_4_enq_bits_data = readResult_4_bits >> {27'h0, readMessageQueue_4_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_4 = _write1HPipe_4_T & ~maskDestinationType ? reorderQueueVec_4_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_5;
  wire              readMessageQueue_5_deq_valid;
  assign readMessageQueue_5_deq_valid = ~_readMessageQueue_fifo_5_empty;
  wire [7:0]        readMessageQueue_dataOut_5_readSource;
  assign reorderQueueVec_5_enq_bits_write1H = readMessageQueue_5_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_5_dataOffset;
  wire [7:0]        readMessageQueue_5_enq_bits_readSource;
  wire [1:0]        readMessageQueue_5_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_5 = {readMessageQueue_5_enq_bits_readSource, readMessageQueue_5_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_5_dataOffset = _readMessageQueue_fifo_5_data_out[1:0];
  assign readMessageQueue_dataOut_5_readSource = _readMessageQueue_fifo_5_data_out[9:2];
  assign readMessageQueue_5_deq_bits_readSource = readMessageQueue_dataOut_5_readSource;
  wire [1:0]        readMessageQueue_5_deq_bits_dataOffset = readMessageQueue_dataOut_5_dataOffset;
  wire              readMessageQueue_5_enq_ready = ~_readMessageQueue_fifo_5_full;
  wire              readMessageQueue_5_enq_valid;
  assign deqAllocate_5 = ~readValid | reorderStageValid & reorderStageState_5 != reorderStageNeed_5;
  assign reorderQueueVec_5_deq_ready = deqAllocate_5;
  assign sourceLane_5 = 8'h1 << _readCrossBar_output_5_bits_writeIndex;
  assign readMessageQueue_5_enq_bits_readSource = sourceLane_5;
  wire              readChannel_5_valid_0 = maskDestinationType ? _maskedWrite_readChannel_5_valid : _readCrossBar_output_5_valid & readMessageQueue_5_enq_ready;
  wire [4:0]        readChannel_5_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_vs : _readCrossBar_output_5_bits_vs;
  wire [1:0]        readChannel_5_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_offset : _readCrossBar_output_5_bits_offset;
  assign readMessageQueue_5_enq_valid = readChannel_5_ready_0 & readChannel_5_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_5_enq_bits_data = readResult_5_bits >> {27'h0, readMessageQueue_5_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_5 = _write1HPipe_5_T & ~maskDestinationType ? reorderQueueVec_5_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_6;
  wire              readMessageQueue_6_deq_valid;
  assign readMessageQueue_6_deq_valid = ~_readMessageQueue_fifo_6_empty;
  wire [7:0]        readMessageQueue_dataOut_6_readSource;
  assign reorderQueueVec_6_enq_bits_write1H = readMessageQueue_6_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_6_dataOffset;
  wire [7:0]        readMessageQueue_6_enq_bits_readSource;
  wire [1:0]        readMessageQueue_6_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_6 = {readMessageQueue_6_enq_bits_readSource, readMessageQueue_6_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_6_dataOffset = _readMessageQueue_fifo_6_data_out[1:0];
  assign readMessageQueue_dataOut_6_readSource = _readMessageQueue_fifo_6_data_out[9:2];
  assign readMessageQueue_6_deq_bits_readSource = readMessageQueue_dataOut_6_readSource;
  wire [1:0]        readMessageQueue_6_deq_bits_dataOffset = readMessageQueue_dataOut_6_dataOffset;
  wire              readMessageQueue_6_enq_ready = ~_readMessageQueue_fifo_6_full;
  wire              readMessageQueue_6_enq_valid;
  assign deqAllocate_6 = ~readValid | reorderStageValid & reorderStageState_6 != reorderStageNeed_6;
  assign reorderQueueVec_6_deq_ready = deqAllocate_6;
  assign sourceLane_6 = 8'h1 << _readCrossBar_output_6_bits_writeIndex;
  assign readMessageQueue_6_enq_bits_readSource = sourceLane_6;
  wire              readChannel_6_valid_0 = maskDestinationType ? _maskedWrite_readChannel_6_valid : _readCrossBar_output_6_valid & readMessageQueue_6_enq_ready;
  wire [4:0]        readChannel_6_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_vs : _readCrossBar_output_6_bits_vs;
  wire [1:0]        readChannel_6_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_offset : _readCrossBar_output_6_bits_offset;
  assign readMessageQueue_6_enq_valid = readChannel_6_ready_0 & readChannel_6_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_6_enq_bits_data = readResult_6_bits >> {27'h0, readMessageQueue_6_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_6 = _write1HPipe_6_T & ~maskDestinationType ? reorderQueueVec_6_deq_bits_write1H : 8'h0;
  wire [7:0]        sourceLane_7;
  wire              readMessageQueue_7_deq_valid;
  assign readMessageQueue_7_deq_valid = ~_readMessageQueue_fifo_7_empty;
  wire [7:0]        readMessageQueue_dataOut_7_readSource;
  assign reorderQueueVec_7_enq_bits_write1H = readMessageQueue_7_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_7_dataOffset;
  wire [7:0]        readMessageQueue_7_enq_bits_readSource;
  wire [1:0]        readMessageQueue_7_enq_bits_dataOffset;
  wire [9:0]        readMessageQueue_dataIn_7 = {readMessageQueue_7_enq_bits_readSource, readMessageQueue_7_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_7_dataOffset = _readMessageQueue_fifo_7_data_out[1:0];
  assign readMessageQueue_dataOut_7_readSource = _readMessageQueue_fifo_7_data_out[9:2];
  assign readMessageQueue_7_deq_bits_readSource = readMessageQueue_dataOut_7_readSource;
  wire [1:0]        readMessageQueue_7_deq_bits_dataOffset = readMessageQueue_dataOut_7_dataOffset;
  wire              readMessageQueue_7_enq_ready = ~_readMessageQueue_fifo_7_full;
  wire              readMessageQueue_7_enq_valid;
  assign deqAllocate_7 = ~readValid | reorderStageValid & reorderStageState_7 != reorderStageNeed_7;
  assign reorderQueueVec_7_deq_ready = deqAllocate_7;
  assign sourceLane_7 = 8'h1 << _readCrossBar_output_7_bits_writeIndex;
  assign readMessageQueue_7_enq_bits_readSource = sourceLane_7;
  wire              readChannel_7_valid_0 = maskDestinationType ? _maskedWrite_readChannel_7_valid : _readCrossBar_output_7_valid & readMessageQueue_7_enq_ready;
  wire [4:0]        readChannel_7_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_vs : _readCrossBar_output_7_bits_vs;
  wire [1:0]        readChannel_7_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_offset : _readCrossBar_output_7_bits_offset;
  assign readMessageQueue_7_enq_valid = readChannel_7_ready_0 & readChannel_7_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_7_enq_bits_data = readResult_7_bits >> {27'h0, readMessageQueue_7_deq_bits_dataOffset, 3'h0};
  wire [7:0]        write1HPipe_7 = _write1HPipe_7_T & ~maskDestinationType ? reorderQueueVec_7_deq_bits_write1H : 8'h0;
  wire [31:0]       readData_data;
  wire              readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_deq_ready;
  wire              readData_readDataQueue_enq_valid;
  wire              readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]       readData_readDataQueue_enq_bits;
  wire [31:0]       readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]        readData_readResultSelect_lo_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]        readData_readResultSelect_lo = {readData_readResultSelect_lo_hi, readData_readResultSelect_lo_lo};
  wire [1:0]        readData_readResultSelect_hi_lo = {write1HPipe_5[0], write1HPipe_4[0]};
  wire [1:0]        readData_readResultSelect_hi_hi = {write1HPipe_7[0], write1HPipe_6[0]};
  wire [3:0]        readData_readResultSelect_hi = {readData_readResultSelect_hi_hi, readData_readResultSelect_hi_lo};
  wire [7:0]        readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire              readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]       readData_data_1;
  wire              isWaiteForThisData_1;
  wire              readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_1_deq_ready;
  wire              readData_readDataQueue_1_enq_valid;
  wire              readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]       readData_readDataQueue_1_enq_bits;
  wire [31:0]       readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]        readData_readResultSelect_lo_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]        readData_readResultSelect_lo_1 = {readData_readResultSelect_lo_hi_1, readData_readResultSelect_lo_lo_1};
  wire [1:0]        readData_readResultSelect_hi_lo_1 = {write1HPipe_5[1], write1HPipe_4[1]};
  wire [1:0]        readData_readResultSelect_hi_hi_1 = {write1HPipe_7[1], write1HPipe_6[1]};
  wire [3:0]        readData_readResultSelect_hi_1 = {readData_readResultSelect_hi_hi_1, readData_readResultSelect_hi_lo_1};
  wire [7:0]        readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_1[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_1[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_1[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_1[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire              readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]       readData_data_2;
  wire              isWaiteForThisData_2;
  wire              readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_2_deq_ready;
  wire              readData_readDataQueue_2_enq_valid;
  wire              readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]       readData_readDataQueue_2_enq_bits;
  wire [31:0]       readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]        readData_readResultSelect_lo_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]        readData_readResultSelect_lo_2 = {readData_readResultSelect_lo_hi_2, readData_readResultSelect_lo_lo_2};
  wire [1:0]        readData_readResultSelect_hi_lo_2 = {write1HPipe_5[2], write1HPipe_4[2]};
  wire [1:0]        readData_readResultSelect_hi_hi_2 = {write1HPipe_7[2], write1HPipe_6[2]};
  wire [3:0]        readData_readResultSelect_hi_2 = {readData_readResultSelect_hi_hi_2, readData_readResultSelect_hi_lo_2};
  wire [7:0]        readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_2[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_2[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_2[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_2[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire              readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]       readData_data_3;
  wire              isWaiteForThisData_3;
  wire              readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire              readData_readDataQueue_3_deq_ready;
  wire              readData_readDataQueue_3_enq_valid;
  wire              readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]       readData_readDataQueue_3_enq_bits;
  wire [31:0]       readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]        readData_readResultSelect_lo_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]        readData_readResultSelect_lo_3 = {readData_readResultSelect_lo_hi_3, readData_readResultSelect_lo_lo_3};
  wire [1:0]        readData_readResultSelect_hi_lo_3 = {write1HPipe_5[3], write1HPipe_4[3]};
  wire [1:0]        readData_readResultSelect_hi_hi_3 = {write1HPipe_7[3], write1HPipe_6[3]};
  wire [3:0]        readData_readResultSelect_hi_3 = {readData_readResultSelect_hi_hi_3, readData_readResultSelect_hi_lo_3};
  wire [7:0]        readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_3[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_3[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_3[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_3[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire              readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  wire [31:0]       readData_data_4;
  wire              isWaiteForThisData_4;
  wire              readData_readDataQueue_4_enq_ready = ~_readData_readDataQueue_fifo_4_full;
  wire              readData_readDataQueue_4_deq_ready;
  wire              readData_readDataQueue_4_enq_valid;
  wire              readData_readDataQueue_4_deq_valid = ~_readData_readDataQueue_fifo_4_empty | readData_readDataQueue_4_enq_valid;
  wire [31:0]       readData_readDataQueue_4_enq_bits;
  wire [31:0]       readData_readDataQueue_4_deq_bits = _readData_readDataQueue_fifo_4_empty ? readData_readDataQueue_4_enq_bits : _readData_readDataQueue_fifo_4_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_4 = {write1HPipe_1[4], write1HPipe_0[4]};
  wire [1:0]        readData_readResultSelect_lo_hi_4 = {write1HPipe_3[4], write1HPipe_2[4]};
  wire [3:0]        readData_readResultSelect_lo_4 = {readData_readResultSelect_lo_hi_4, readData_readResultSelect_lo_lo_4};
  wire [1:0]        readData_readResultSelect_hi_lo_4 = {write1HPipe_5[4], write1HPipe_4[4]};
  wire [1:0]        readData_readResultSelect_hi_hi_4 = {write1HPipe_7[4], write1HPipe_6[4]};
  wire [3:0]        readData_readResultSelect_hi_4 = {readData_readResultSelect_hi_hi_4, readData_readResultSelect_hi_lo_4};
  wire [7:0]        readData_readResultSelect_4 = {readData_readResultSelect_hi_4, readData_readResultSelect_lo_4};
  assign readData_data_4 =
    (readData_readResultSelect_4[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_4[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_4[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_4[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_4[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_4[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_4[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_4[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_4_enq_bits = readData_data_4;
  wire              readTokenRelease_4 = readData_readDataQueue_4_deq_ready & readData_readDataQueue_4_deq_valid;
  assign readData_readDataQueue_4_enq_valid = |readData_readResultSelect_4;
  wire [31:0]       readData_data_5;
  wire              isWaiteForThisData_5;
  wire              readData_readDataQueue_5_enq_ready = ~_readData_readDataQueue_fifo_5_full;
  wire              readData_readDataQueue_5_deq_ready;
  wire              readData_readDataQueue_5_enq_valid;
  wire              readData_readDataQueue_5_deq_valid = ~_readData_readDataQueue_fifo_5_empty | readData_readDataQueue_5_enq_valid;
  wire [31:0]       readData_readDataQueue_5_enq_bits;
  wire [31:0]       readData_readDataQueue_5_deq_bits = _readData_readDataQueue_fifo_5_empty ? readData_readDataQueue_5_enq_bits : _readData_readDataQueue_fifo_5_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_5 = {write1HPipe_1[5], write1HPipe_0[5]};
  wire [1:0]        readData_readResultSelect_lo_hi_5 = {write1HPipe_3[5], write1HPipe_2[5]};
  wire [3:0]        readData_readResultSelect_lo_5 = {readData_readResultSelect_lo_hi_5, readData_readResultSelect_lo_lo_5};
  wire [1:0]        readData_readResultSelect_hi_lo_5 = {write1HPipe_5[5], write1HPipe_4[5]};
  wire [1:0]        readData_readResultSelect_hi_hi_5 = {write1HPipe_7[5], write1HPipe_6[5]};
  wire [3:0]        readData_readResultSelect_hi_5 = {readData_readResultSelect_hi_hi_5, readData_readResultSelect_hi_lo_5};
  wire [7:0]        readData_readResultSelect_5 = {readData_readResultSelect_hi_5, readData_readResultSelect_lo_5};
  assign readData_data_5 =
    (readData_readResultSelect_5[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_5[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_5[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_5[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_5[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_5[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_5[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_5[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_5_enq_bits = readData_data_5;
  wire              readTokenRelease_5 = readData_readDataQueue_5_deq_ready & readData_readDataQueue_5_deq_valid;
  assign readData_readDataQueue_5_enq_valid = |readData_readResultSelect_5;
  wire [31:0]       readData_data_6;
  wire              isWaiteForThisData_6;
  wire              readData_readDataQueue_6_enq_ready = ~_readData_readDataQueue_fifo_6_full;
  wire              readData_readDataQueue_6_deq_ready;
  wire              readData_readDataQueue_6_enq_valid;
  wire              readData_readDataQueue_6_deq_valid = ~_readData_readDataQueue_fifo_6_empty | readData_readDataQueue_6_enq_valid;
  wire [31:0]       readData_readDataQueue_6_enq_bits;
  wire [31:0]       readData_readDataQueue_6_deq_bits = _readData_readDataQueue_fifo_6_empty ? readData_readDataQueue_6_enq_bits : _readData_readDataQueue_fifo_6_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_6 = {write1HPipe_1[6], write1HPipe_0[6]};
  wire [1:0]        readData_readResultSelect_lo_hi_6 = {write1HPipe_3[6], write1HPipe_2[6]};
  wire [3:0]        readData_readResultSelect_lo_6 = {readData_readResultSelect_lo_hi_6, readData_readResultSelect_lo_lo_6};
  wire [1:0]        readData_readResultSelect_hi_lo_6 = {write1HPipe_5[6], write1HPipe_4[6]};
  wire [1:0]        readData_readResultSelect_hi_hi_6 = {write1HPipe_7[6], write1HPipe_6[6]};
  wire [3:0]        readData_readResultSelect_hi_6 = {readData_readResultSelect_hi_hi_6, readData_readResultSelect_hi_lo_6};
  wire [7:0]        readData_readResultSelect_6 = {readData_readResultSelect_hi_6, readData_readResultSelect_lo_6};
  assign readData_data_6 =
    (readData_readResultSelect_6[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_6[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_6[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_6[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_6[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_6[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_6[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_6[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_6_enq_bits = readData_data_6;
  wire              readTokenRelease_6 = readData_readDataQueue_6_deq_ready & readData_readDataQueue_6_deq_valid;
  assign readData_readDataQueue_6_enq_valid = |readData_readResultSelect_6;
  wire [31:0]       readData_data_7;
  wire              isWaiteForThisData_7;
  wire              readData_readDataQueue_7_enq_ready = ~_readData_readDataQueue_fifo_7_full;
  wire              readData_readDataQueue_7_deq_ready;
  wire              readData_readDataQueue_7_enq_valid;
  wire              readData_readDataQueue_7_deq_valid = ~_readData_readDataQueue_fifo_7_empty | readData_readDataQueue_7_enq_valid;
  wire [31:0]       readData_readDataQueue_7_enq_bits;
  wire [31:0]       readData_readDataQueue_7_deq_bits = _readData_readDataQueue_fifo_7_empty ? readData_readDataQueue_7_enq_bits : _readData_readDataQueue_fifo_7_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_7 = {write1HPipe_1[7], write1HPipe_0[7]};
  wire [1:0]        readData_readResultSelect_lo_hi_7 = {write1HPipe_3[7], write1HPipe_2[7]};
  wire [3:0]        readData_readResultSelect_lo_7 = {readData_readResultSelect_lo_hi_7, readData_readResultSelect_lo_lo_7};
  wire [1:0]        readData_readResultSelect_hi_lo_7 = {write1HPipe_5[7], write1HPipe_4[7]};
  wire [1:0]        readData_readResultSelect_hi_hi_7 = {write1HPipe_7[7], write1HPipe_6[7]};
  wire [3:0]        readData_readResultSelect_hi_7 = {readData_readResultSelect_hi_hi_7, readData_readResultSelect_hi_lo_7};
  wire [7:0]        readData_readResultSelect_7 = {readData_readResultSelect_hi_7, readData_readResultSelect_lo_7};
  assign readData_data_7 =
    (readData_readResultSelect_7[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_7[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_7[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_7[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_7[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_7[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_7[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_7[7] ? dataAfterReorderCheck_7 : 32'h0);
  assign readData_readDataQueue_7_enq_bits = readData_data_7;
  wire              readTokenRelease_7 = readData_readDataQueue_7_deq_ready & readData_readDataQueue_7_deq_valid;
  assign readData_readDataQueue_7_enq_valid = |readData_readResultSelect_7;
  reg  [7:0]        waiteReadDataPipeReg_executeGroup;
  reg  [7:0]        waiteReadDataPipeReg_sourceValid;
  reg  [7:0]        waiteReadDataPipeReg_replaceVs1;
  reg  [7:0]        waiteReadDataPipeReg_needRead;
  reg               waiteReadDataPipeReg_last;
  reg  [31:0]       waiteReadData_0;
  reg  [31:0]       waiteReadData_1;
  reg  [31:0]       waiteReadData_2;
  reg  [31:0]       waiteReadData_3;
  reg  [31:0]       waiteReadData_4;
  reg  [31:0]       waiteReadData_5;
  reg  [31:0]       waiteReadData_6;
  reg  [31:0]       waiteReadData_7;
  reg  [7:0]        waiteReadSate;
  reg               waiteReadStageValid;
  wire [1:0]        executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]        executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire              writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_16 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]       _GEN_80 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_80;
  wire [31:0]       writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_80;
  wire [31:0]       writeDataVec_data_unreadData_16;
  assign writeDataVec_data_unreadData_16 = _GEN_80;
  wire [7:0]        writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire              writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_17 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]       _GEN_81 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_81;
  wire [31:0]       writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_81;
  wire [31:0]       writeDataVec_data_unreadData_17;
  assign writeDataVec_data_unreadData_17 = _GEN_81;
  wire [7:0]        writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire              writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_18 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]       _GEN_82 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_82;
  wire [31:0]       writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_82;
  wire [31:0]       writeDataVec_data_unreadData_18;
  assign writeDataVec_data_unreadData_18 = _GEN_82;
  wire [7:0]        writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire              writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_19 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]       _GEN_83 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_83;
  wire [31:0]       writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_83;
  wire [31:0]       writeDataVec_data_unreadData_19;
  assign writeDataVec_data_unreadData_19 = _GEN_83;
  wire [7:0]        writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire              writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[4];
  wire              writeDataVec_data_dataIsRead_12 = waiteReadDataPipeReg_needRead[4];
  wire              writeDataVec_data_dataIsRead_20 = waiteReadDataPipeReg_needRead[4];
  wire [31:0]       _GEN_84 = waiteReadDataPipeReg_replaceVs1[4] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_84;
  wire [31:0]       writeDataVec_data_unreadData_12;
  assign writeDataVec_data_unreadData_12 = _GEN_84;
  wire [31:0]       writeDataVec_data_unreadData_20;
  assign writeDataVec_data_unreadData_20 = _GEN_84;
  wire [7:0]        writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_4[7:0] : writeDataVec_data_unreadData_4[7:0];
  wire              writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[5];
  wire              writeDataVec_data_dataIsRead_13 = waiteReadDataPipeReg_needRead[5];
  wire              writeDataVec_data_dataIsRead_21 = waiteReadDataPipeReg_needRead[5];
  wire [31:0]       _GEN_85 = waiteReadDataPipeReg_replaceVs1[5] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_85;
  wire [31:0]       writeDataVec_data_unreadData_13;
  assign writeDataVec_data_unreadData_13 = _GEN_85;
  wire [31:0]       writeDataVec_data_unreadData_21;
  assign writeDataVec_data_unreadData_21 = _GEN_85;
  wire [7:0]        writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_5[7:0] : writeDataVec_data_unreadData_5[7:0];
  wire              writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[6];
  wire              writeDataVec_data_dataIsRead_14 = waiteReadDataPipeReg_needRead[6];
  wire              writeDataVec_data_dataIsRead_22 = waiteReadDataPipeReg_needRead[6];
  wire [31:0]       _GEN_86 = waiteReadDataPipeReg_replaceVs1[6] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_86;
  wire [31:0]       writeDataVec_data_unreadData_14;
  assign writeDataVec_data_unreadData_14 = _GEN_86;
  wire [31:0]       writeDataVec_data_unreadData_22;
  assign writeDataVec_data_unreadData_22 = _GEN_86;
  wire [7:0]        writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_6[7:0] : writeDataVec_data_unreadData_6[7:0];
  wire              writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[7];
  wire              writeDataVec_data_dataIsRead_15 = waiteReadDataPipeReg_needRead[7];
  wire              writeDataVec_data_dataIsRead_23 = waiteReadDataPipeReg_needRead[7];
  wire [31:0]       _GEN_87 = waiteReadDataPipeReg_replaceVs1[7] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_87;
  wire [31:0]       writeDataVec_data_unreadData_15;
  assign writeDataVec_data_unreadData_15 = _GEN_87;
  wire [31:0]       writeDataVec_data_unreadData_23;
  assign writeDataVec_data_unreadData_23 = _GEN_87;
  wire [7:0]        writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_7[7:0] : writeDataVec_data_unreadData_7[7:0];
  wire [15:0]       writeDataVec_data_lo_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]       writeDataVec_data_lo_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]       writeDataVec_data_lo = {writeDataVec_data_lo_hi, writeDataVec_data_lo_lo};
  wire [15:0]       writeDataVec_data_hi_lo = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [15:0]       writeDataVec_data_hi_hi = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [31:0]       writeDataVec_data_hi = {writeDataVec_data_hi_hi, writeDataVec_data_hi_lo};
  wire [63:0]       writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [318:0]      writeDataVec_shifterData = {255'h0, writeDataVec_data} << {311'h0, executeIndexVec_0, 6'h0};
  wire [255:0]      writeDataVec_0 = writeDataVec_shifterData[255:0];
  wire [15:0]       writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_8[15:0];
  wire [15:0]       writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_9[15:0];
  wire [15:0]       writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_10[15:0];
  wire [15:0]       writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_11[15:0];
  wire [15:0]       writeDataVec_data_dataElement_12 = writeDataVec_data_dataIsRead_12 ? waiteReadData_4[15:0] : writeDataVec_data_unreadData_12[15:0];
  wire [15:0]       writeDataVec_data_dataElement_13 = writeDataVec_data_dataIsRead_13 ? waiteReadData_5[15:0] : writeDataVec_data_unreadData_13[15:0];
  wire [15:0]       writeDataVec_data_dataElement_14 = writeDataVec_data_dataIsRead_14 ? waiteReadData_6[15:0] : writeDataVec_data_unreadData_14[15:0];
  wire [15:0]       writeDataVec_data_dataElement_15 = writeDataVec_data_dataIsRead_15 ? waiteReadData_7[15:0] : writeDataVec_data_unreadData_15[15:0];
  wire [31:0]       writeDataVec_data_lo_lo_1 = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [31:0]       writeDataVec_data_lo_hi_1 = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [63:0]       writeDataVec_data_lo_1 = {writeDataVec_data_lo_hi_1, writeDataVec_data_lo_lo_1};
  wire [31:0]       writeDataVec_data_hi_lo_1 = {writeDataVec_data_dataElement_13, writeDataVec_data_dataElement_12};
  wire [31:0]       writeDataVec_data_hi_hi_1 = {writeDataVec_data_dataElement_15, writeDataVec_data_dataElement_14};
  wire [63:0]       writeDataVec_data_hi_1 = {writeDataVec_data_hi_hi_1, writeDataVec_data_hi_lo_1};
  wire [127:0]      writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [382:0]      writeDataVec_shifterData_1 = {255'h0, writeDataVec_data_1} << {375'h0, executeIndexVec_1, 6'h0};
  wire [255:0]      writeDataVec_1 = writeDataVec_shifterData_1[255:0];
  wire [31:0]       writeDataVec_data_dataElement_16 = writeDataVec_data_dataIsRead_16 ? waiteReadData_0 : writeDataVec_data_unreadData_16;
  wire [31:0]       writeDataVec_data_dataElement_17 = writeDataVec_data_dataIsRead_17 ? waiteReadData_1 : writeDataVec_data_unreadData_17;
  wire [31:0]       writeDataVec_data_dataElement_18 = writeDataVec_data_dataIsRead_18 ? waiteReadData_2 : writeDataVec_data_unreadData_18;
  wire [31:0]       writeDataVec_data_dataElement_19 = writeDataVec_data_dataIsRead_19 ? waiteReadData_3 : writeDataVec_data_unreadData_19;
  wire [31:0]       writeDataVec_data_dataElement_20 = writeDataVec_data_dataIsRead_20 ? waiteReadData_4 : writeDataVec_data_unreadData_20;
  wire [31:0]       writeDataVec_data_dataElement_21 = writeDataVec_data_dataIsRead_21 ? waiteReadData_5 : writeDataVec_data_unreadData_21;
  wire [31:0]       writeDataVec_data_dataElement_22 = writeDataVec_data_dataIsRead_22 ? waiteReadData_6 : writeDataVec_data_unreadData_22;
  wire [31:0]       writeDataVec_data_dataElement_23 = writeDataVec_data_dataIsRead_23 ? waiteReadData_7 : writeDataVec_data_unreadData_23;
  wire [63:0]       writeDataVec_data_lo_lo_2 = {writeDataVec_data_dataElement_17, writeDataVec_data_dataElement_16};
  wire [63:0]       writeDataVec_data_lo_hi_2 = {writeDataVec_data_dataElement_19, writeDataVec_data_dataElement_18};
  wire [127:0]      writeDataVec_data_lo_2 = {writeDataVec_data_lo_hi_2, writeDataVec_data_lo_lo_2};
  wire [63:0]       writeDataVec_data_hi_lo_2 = {writeDataVec_data_dataElement_21, writeDataVec_data_dataElement_20};
  wire [63:0]       writeDataVec_data_hi_hi_2 = {writeDataVec_data_dataElement_23, writeDataVec_data_dataElement_22};
  wire [127:0]      writeDataVec_data_hi_2 = {writeDataVec_data_hi_hi_2, writeDataVec_data_hi_lo_2};
  wire [255:0]      writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [382:0]      writeDataVec_shifterData_2 = {127'h0, writeDataVec_data_2};
  wire [255:0]      writeDataVec_2 = writeDataVec_shifterData_2[255:0];
  wire [255:0]      writeData = (sew1H[0] ? writeDataVec_0 : 256'h0) | (sew1H[1] ? writeDataVec_1 : 256'h0) | (sew1H[2] ? writeDataVec_2 : 256'h0);
  wire [1:0]        writeMaskVec_mask_lo_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]        writeMaskVec_mask_lo_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]        writeMaskVec_mask_lo = {writeMaskVec_mask_lo_hi, writeMaskVec_mask_lo_lo};
  wire [1:0]        writeMaskVec_mask_hi_lo = waiteReadDataPipeReg_sourceValid[5:4];
  wire [1:0]        writeMaskVec_mask_hi_hi = waiteReadDataPipeReg_sourceValid[7:6];
  wire [3:0]        writeMaskVec_mask_hi = {writeMaskVec_mask_hi_hi, writeMaskVec_mask_hi_lo};
  wire [7:0]        writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [38:0]       writeMaskVec_shifterMask = {31'h0, writeMaskVec_mask} << {34'h0, executeIndexVec_0, 3'h0};
  wire [31:0]       writeMaskVec_0 = writeMaskVec_shifterMask[31:0];
  wire [3:0]        writeMaskVec_mask_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]        writeMaskVec_mask_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]        writeMaskVec_mask_lo_1 = {writeMaskVec_mask_lo_hi_1, writeMaskVec_mask_lo_lo_1};
  wire [3:0]        writeMaskVec_mask_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[5]}}, {2{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [3:0]        writeMaskVec_mask_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[7]}}, {2{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [7:0]        writeMaskVec_mask_hi_1 = {writeMaskVec_mask_hi_hi_1, writeMaskVec_mask_hi_lo_1};
  wire [15:0]       writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [46:0]       writeMaskVec_shifterMask_1 = {31'h0, writeMaskVec_mask_1} << {42'h0, executeIndexVec_1, 3'h0};
  wire [31:0]       writeMaskVec_1 = writeMaskVec_shifterMask_1[31:0];
  wire [7:0]        writeMaskVec_mask_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]        writeMaskVec_mask_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]       writeMaskVec_mask_lo_2 = {writeMaskVec_mask_lo_hi_2, writeMaskVec_mask_lo_lo_2};
  wire [7:0]        writeMaskVec_mask_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[5]}}, {4{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [7:0]        writeMaskVec_mask_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[7]}}, {4{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [15:0]       writeMaskVec_mask_hi_2 = {writeMaskVec_mask_hi_hi_2, writeMaskVec_mask_hi_lo_2};
  wire [31:0]       writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [46:0]       writeMaskVec_shifterMask_2 = {15'h0, writeMaskVec_mask_2};
  wire [31:0]       writeMaskVec_2 = writeMaskVec_shifterMask_2[31:0];
  wire [31:0]       writeMask = (sew1H[0] ? writeMaskVec_0 : 32'h0) | (sew1H[1] ? writeMaskVec_1 : 32'h0) | (sew1H[2] ? writeMaskVec_2 : 32'h0);
  wire [10:0]       _writeRequest_res_writeData_groupCounter_T_14 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [5:0]        writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_4_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_5_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_6_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [5:0]        writeRequest_7_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_14[7:2];
  wire [31:0]       writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]       writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]       writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]       writeRequest_3_writeData_data = writeData[127:96];
  wire [31:0]       writeRequest_4_writeData_data = writeData[159:128];
  wire [31:0]       writeRequest_5_writeData_data = writeData[191:160];
  wire [31:0]       writeRequest_6_writeData_data = writeData[223:192];
  wire [31:0]       writeRequest_7_writeData_data = writeData[255:224];
  wire [3:0]        writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]        writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]        writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]        writeRequest_3_writeData_mask = writeMask[15:12];
  wire [3:0]        writeRequest_4_writeData_mask = writeMask[19:16];
  wire [3:0]        writeRequest_5_writeData_mask = writeMask[23:20];
  wire [3:0]        writeRequest_6_writeData_mask = writeMask[27:24];
  wire [3:0]        writeRequest_7_writeData_mask = writeMask[31:28];
  wire [1:0]        WillWriteLane_lo_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]        WillWriteLane_lo_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]        WillWriteLane_lo = {WillWriteLane_lo_hi, WillWriteLane_lo_lo};
  wire [1:0]        WillWriteLane_hi_lo = {|writeRequest_5_writeData_mask, |writeRequest_4_writeData_mask};
  wire [1:0]        WillWriteLane_hi_hi = {|writeRequest_7_writeData_mask, |writeRequest_6_writeData_mask};
  wire [3:0]        WillWriteLane_hi = {WillWriteLane_hi_hi, WillWriteLane_hi_lo};
  wire [7:0]        WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire              waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 8'h0);
  wire              waiteStageDeqReady;
  wire              waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire              waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire              isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  assign isWaiteForThisData_4 = waiteReadDataPipeReg_needRead[4] & ~(waiteReadSate[4]) & waiteReadStageValid;
  assign readData_readDataQueue_4_deq_ready = isWaiteForThisData_4;
  assign isWaiteForThisData_5 = waiteReadDataPipeReg_needRead[5] & ~(waiteReadSate[5]) & waiteReadStageValid;
  assign readData_readDataQueue_5_deq_ready = isWaiteForThisData_5;
  assign isWaiteForThisData_6 = waiteReadDataPipeReg_needRead[6] & ~(waiteReadSate[6]) & waiteReadStageValid;
  assign readData_readDataQueue_6_deq_ready = isWaiteForThisData_6;
  assign isWaiteForThisData_7 = waiteReadDataPipeReg_needRead[7] & ~(waiteReadSate[7]) & waiteReadStageValid;
  assign readData_readDataQueue_7_deq_ready = isWaiteForThisData_7;
  wire [1:0]        readResultValid_lo_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]        readResultValid_lo_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]        readResultValid_lo = {readResultValid_lo_hi, readResultValid_lo_lo};
  wire [1:0]        readResultValid_hi_lo = {readTokenRelease_5, readTokenRelease_4};
  wire [1:0]        readResultValid_hi_hi = {readTokenRelease_7, readTokenRelease_6};
  wire [3:0]        readResultValid_hi = {readResultValid_hi_hi, readResultValid_hi_lo};
  wire [7:0]        readResultValid = {readResultValid_hi, readResultValid_lo};
  wire              executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]       source2_lo_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]       source2_lo_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]      source2_lo = {source2_lo_hi, source2_lo_lo};
  wire [63:0]       source2_hi_lo = {exeReqReg_5_bits_source2, exeReqReg_4_bits_source2};
  wire [63:0]       source2_hi_hi = {exeReqReg_7_bits_source2, exeReqReg_6_bits_source2};
  wire [127:0]      source2_hi = {source2_hi_hi, source2_hi_lo};
  wire [255:0]      source2 = {source2_hi, source2_lo};
  wire [127:0]      source1_lo = {source1_lo_hi, source1_lo_lo};
  wire [127:0]      source1_hi = {source1_hi_hi, source1_hi_lo};
  wire [255:0]      source1 = {source1_hi, source1_lo};
  wire              vs1Split_vs1SetIndex = requestCounter[0];
  wire              vs1Split_1_2 = vs1Split_vs1SetIndex;
  wire              vs1Split_2_2 = &vs1Split_vs1SetIndex_1;
  wire [31:0]       _compressSource1_T_3 = sew1H[0] ? readVS1Reg_data : 32'h0;
  wire [3:0][7:0]   _GEN_91 = {{readVS1Reg_data[31:24]}, {readVS1Reg_data[23:16]}, {readVS1Reg_data[15:8]}, {readVS1Reg_data[7:0]}};
  wire [15:0]       _GEN_92 = _compressSource1_T_3[15:0] | (sew1H[1] ? (vs1Split_vs1SetIndex ? readVS1Reg_data[31:16] : readVS1Reg_data[15:0]) : 16'h0);
  wire [31:0]       compressSource1 = {_compressSource1_T_3[31:16], _GEN_92[15:8], _GEN_92[7:0] | (sew1H[2] ? _GEN_91[vs1Split_vs1SetIndex_1] : 8'h0)};
  wire [31:0]       source1Select = mv ? readVS1Reg_data : compressSource1;
  wire              source1Change = sew1H[0] | sew1H[1] & vs1Split_1_2 | sew1H[2] & vs1Split_2_2;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]        view__in_bits_ffoInput_lo_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_lo_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_lo = {view__in_bits_ffoInput_lo_hi, view__in_bits_ffoInput_lo_lo};
  wire [1:0]        view__in_bits_ffoInput_hi_lo = {exeReqReg_5_bits_ffo, exeReqReg_4_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_hi_hi = {exeReqReg_7_bits_ffo, exeReqReg_6_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_hi = {view__in_bits_ffoInput_hi_hi, view__in_bits_ffoInput_hi_lo};
  wire [3:0]        view__in_bits_validInput_lo = {view__in_bits_validInput_lo_hi, view__in_bits_validInput_lo_lo};
  wire [3:0]        view__in_bits_validInput_hi = {view__in_bits_validInput_hi_hi, view__in_bits_validInput_hi_lo};
  wire              reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire [3:0]        view__in_bits_sourceValid_lo = {view__in_bits_sourceValid_lo_hi, view__in_bits_sourceValid_lo_lo};
  wire [3:0]        view__in_bits_sourceValid_hi = {view__in_bits_sourceValid_hi_hi, view__in_bits_sourceValid_hi_lo};
  wire              _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [1:0]        view__in_bits_fpSourceValid_lo_lo = {exeReqReg_1_bits_fpReduceValid, exeReqReg_0_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_lo_hi = {exeReqReg_3_bits_fpReduceValid, exeReqReg_2_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_lo = {view__in_bits_fpSourceValid_lo_hi, view__in_bits_fpSourceValid_lo_lo};
  wire [1:0]        view__in_bits_fpSourceValid_hi_lo = {exeReqReg_5_bits_fpReduceValid, exeReqReg_4_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_hi_hi = {exeReqReg_7_bits_fpReduceValid, exeReqReg_6_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_hi = {view__in_bits_fpSourceValid_hi_hi, view__in_bits_fpSourceValid_hi_lo};
  wire [7:0]        extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [255:0]      _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 256'h0;
  wire [255:0]      executeResult = {_executeResult_T_4[255:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 256'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  wire [3:0]        compressUnitResultQueue_deq_ready_lo = {compressUnitResultQueue_deq_ready_lo_hi, compressUnitResultQueue_deq_ready_lo_lo};
  wire [3:0]        compressUnitResultQueue_deq_ready_hi = {compressUnitResultQueue_deq_ready_hi_hi, compressUnitResultQueue_deq_ready_hi_lo};
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire              compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire              executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 6'h0) | (unitType[3] ? extendGroupCount[5:0] : 6'h0);
  wire [7:0]        executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 6'h0) | (unitType[2] ? requestCounter : 6'h0)} | (unitType[3] ? extendGroupCount : 8'h0);
  wire [31:0]       executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire              maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire              maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire              maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire              maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  wire              maskFilter_4 = |{~maskDestinationType, currentMaskGroupForDestination[159:128]};
  wire              maskFilter_5 = |{~maskDestinationType, currentMaskGroupForDestination[191:160]};
  wire              maskFilter_6 = |{~maskDestinationType, currentMaskGroupForDestination[223:192]};
  wire              maskFilter_7 = |{~maskDestinationType, currentMaskGroupForDestination[255:224]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire              exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire              writeQueue_dataOut_ffoByOther;
  wire [31:0]       writeQueue_dataOut_writeData_data;
  wire [31:0]       exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_writeData_mask;
  wire [3:0]        exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_dataOut_index;
  wire [5:0]        writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_0_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_0_enq_bits_writeData_data;
  wire [3:0]        writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire              writeQueue_0_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [50:0]       writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[13:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[17:14];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[49:18];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[50];
  wire              writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [5:0]        writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire              writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire              writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire              exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire              writeQueue_dataOut_1_ffoByOther;
  wire [31:0]       writeQueue_dataOut_1_writeData_data;
  wire [31:0]       exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_1_writeData_mask;
  wire [3:0]        exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_dataOut_1_index;
  wire [5:0]        writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_1_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_1_enq_bits_writeData_data;
  wire [3:0]        writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire              writeQueue_1_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [50:0]       writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[13:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[17:14];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[49:18];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[50];
  wire              writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [5:0]        writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire              writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire              writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire              exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire              writeQueue_dataOut_2_ffoByOther;
  wire [31:0]       writeQueue_dataOut_2_writeData_data;
  wire [31:0]       exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_2_writeData_mask;
  wire [3:0]        exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_dataOut_2_index;
  wire [5:0]        writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_2_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_2_enq_bits_writeData_data;
  wire [3:0]        writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire              writeQueue_2_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [50:0]       writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[13:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[17:14];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[49:18];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[50];
  wire              writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [5:0]        writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire              writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire              writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire              exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire              writeQueue_dataOut_3_ffoByOther;
  wire [31:0]       writeQueue_dataOut_3_writeData_data;
  wire [31:0]       exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_3_writeData_mask;
  wire [3:0]        exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_dataOut_3_index;
  wire [5:0]        writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_3_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_3_enq_bits_writeData_data;
  wire [3:0]        writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire              writeQueue_3_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [50:0]       writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[13:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[17:14];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[49:18];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[50];
  wire              writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [5:0]        writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire              writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire              writeQueue_3_enq_valid;
  assign writeQueue_4_deq_valid = ~_writeQueue_fifo_4_empty;
  wire              exeResp_4_valid_0 = writeQueue_4_deq_valid;
  wire              writeQueue_dataOut_4_ffoByOther;
  wire [31:0]       writeQueue_dataOut_4_writeData_data;
  wire [31:0]       exeResp_4_bits_data_0 = writeQueue_4_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_4_writeData_mask;
  wire [3:0]        exeResp_4_bits_mask_0 = writeQueue_4_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_4_writeData_vd;
  wire [2:0]        writeQueue_dataOut_4_index;
  wire [5:0]        writeQueue_4_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_4_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_4 = {writeQueue_4_enq_bits_writeData_groupCounter, writeQueue_4_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_4_enq_bits_writeData_data;
  wire [3:0]        writeQueue_4_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_8 = {writeQueue_4_enq_bits_writeData_data, writeQueue_4_enq_bits_writeData_mask};
  wire              writeQueue_4_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_9 = {writeQueue_4_enq_bits_ffoByOther, writeQueue_dataIn_hi_8, writeQueue_dataIn_lo_4};
  wire [50:0]       writeQueue_dataIn_4 = {writeQueue_dataIn_hi_9, writeQueue_4_enq_bits_index};
  assign writeQueue_dataOut_4_index = _writeQueue_fifo_4_data_out[2:0];
  assign writeQueue_dataOut_4_writeData_vd = _writeQueue_fifo_4_data_out[7:3];
  assign writeQueue_dataOut_4_writeData_groupCounter = _writeQueue_fifo_4_data_out[13:8];
  assign writeQueue_dataOut_4_writeData_mask = _writeQueue_fifo_4_data_out[17:14];
  assign writeQueue_dataOut_4_writeData_data = _writeQueue_fifo_4_data_out[49:18];
  assign writeQueue_dataOut_4_ffoByOther = _writeQueue_fifo_4_data_out[50];
  wire              writeQueue_4_deq_bits_ffoByOther = writeQueue_dataOut_4_ffoByOther;
  assign writeQueue_4_deq_bits_writeData_data = writeQueue_dataOut_4_writeData_data;
  assign writeQueue_4_deq_bits_writeData_mask = writeQueue_dataOut_4_writeData_mask;
  wire [5:0]        writeQueue_4_deq_bits_writeData_groupCounter = writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]        writeQueue_4_deq_bits_writeData_vd = writeQueue_dataOut_4_writeData_vd;
  wire [2:0]        writeQueue_4_deq_bits_index = writeQueue_dataOut_4_index;
  wire              writeQueue_4_enq_ready = ~_writeQueue_fifo_4_full;
  wire              writeQueue_4_enq_valid;
  assign writeQueue_5_deq_valid = ~_writeQueue_fifo_5_empty;
  wire              exeResp_5_valid_0 = writeQueue_5_deq_valid;
  wire              writeQueue_dataOut_5_ffoByOther;
  wire [31:0]       writeQueue_dataOut_5_writeData_data;
  wire [31:0]       exeResp_5_bits_data_0 = writeQueue_5_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_5_writeData_mask;
  wire [3:0]        exeResp_5_bits_mask_0 = writeQueue_5_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_5_writeData_vd;
  wire [2:0]        writeQueue_dataOut_5_index;
  wire [5:0]        writeQueue_5_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_5_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_5 = {writeQueue_5_enq_bits_writeData_groupCounter, writeQueue_5_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_5_enq_bits_writeData_data;
  wire [3:0]        writeQueue_5_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_10 = {writeQueue_5_enq_bits_writeData_data, writeQueue_5_enq_bits_writeData_mask};
  wire              writeQueue_5_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_11 = {writeQueue_5_enq_bits_ffoByOther, writeQueue_dataIn_hi_10, writeQueue_dataIn_lo_5};
  wire [50:0]       writeQueue_dataIn_5 = {writeQueue_dataIn_hi_11, writeQueue_5_enq_bits_index};
  assign writeQueue_dataOut_5_index = _writeQueue_fifo_5_data_out[2:0];
  assign writeQueue_dataOut_5_writeData_vd = _writeQueue_fifo_5_data_out[7:3];
  assign writeQueue_dataOut_5_writeData_groupCounter = _writeQueue_fifo_5_data_out[13:8];
  assign writeQueue_dataOut_5_writeData_mask = _writeQueue_fifo_5_data_out[17:14];
  assign writeQueue_dataOut_5_writeData_data = _writeQueue_fifo_5_data_out[49:18];
  assign writeQueue_dataOut_5_ffoByOther = _writeQueue_fifo_5_data_out[50];
  wire              writeQueue_5_deq_bits_ffoByOther = writeQueue_dataOut_5_ffoByOther;
  assign writeQueue_5_deq_bits_writeData_data = writeQueue_dataOut_5_writeData_data;
  assign writeQueue_5_deq_bits_writeData_mask = writeQueue_dataOut_5_writeData_mask;
  wire [5:0]        writeQueue_5_deq_bits_writeData_groupCounter = writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]        writeQueue_5_deq_bits_writeData_vd = writeQueue_dataOut_5_writeData_vd;
  wire [2:0]        writeQueue_5_deq_bits_index = writeQueue_dataOut_5_index;
  wire              writeQueue_5_enq_ready = ~_writeQueue_fifo_5_full;
  wire              writeQueue_5_enq_valid;
  assign writeQueue_6_deq_valid = ~_writeQueue_fifo_6_empty;
  wire              exeResp_6_valid_0 = writeQueue_6_deq_valid;
  wire              writeQueue_dataOut_6_ffoByOther;
  wire [31:0]       writeQueue_dataOut_6_writeData_data;
  wire [31:0]       exeResp_6_bits_data_0 = writeQueue_6_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_6_writeData_mask;
  wire [3:0]        exeResp_6_bits_mask_0 = writeQueue_6_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_6_writeData_vd;
  wire [2:0]        writeQueue_dataOut_6_index;
  wire [5:0]        writeQueue_6_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_6_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_6 = {writeQueue_6_enq_bits_writeData_groupCounter, writeQueue_6_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_6_enq_bits_writeData_data;
  wire [3:0]        writeQueue_6_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_12 = {writeQueue_6_enq_bits_writeData_data, writeQueue_6_enq_bits_writeData_mask};
  wire              writeQueue_6_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_13 = {writeQueue_6_enq_bits_ffoByOther, writeQueue_dataIn_hi_12, writeQueue_dataIn_lo_6};
  wire [50:0]       writeQueue_dataIn_6 = {writeQueue_dataIn_hi_13, writeQueue_6_enq_bits_index};
  assign writeQueue_dataOut_6_index = _writeQueue_fifo_6_data_out[2:0];
  assign writeQueue_dataOut_6_writeData_vd = _writeQueue_fifo_6_data_out[7:3];
  assign writeQueue_dataOut_6_writeData_groupCounter = _writeQueue_fifo_6_data_out[13:8];
  assign writeQueue_dataOut_6_writeData_mask = _writeQueue_fifo_6_data_out[17:14];
  assign writeQueue_dataOut_6_writeData_data = _writeQueue_fifo_6_data_out[49:18];
  assign writeQueue_dataOut_6_ffoByOther = _writeQueue_fifo_6_data_out[50];
  wire              writeQueue_6_deq_bits_ffoByOther = writeQueue_dataOut_6_ffoByOther;
  assign writeQueue_6_deq_bits_writeData_data = writeQueue_dataOut_6_writeData_data;
  assign writeQueue_6_deq_bits_writeData_mask = writeQueue_dataOut_6_writeData_mask;
  wire [5:0]        writeQueue_6_deq_bits_writeData_groupCounter = writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]        writeQueue_6_deq_bits_writeData_vd = writeQueue_dataOut_6_writeData_vd;
  wire [2:0]        writeQueue_6_deq_bits_index = writeQueue_dataOut_6_index;
  wire              writeQueue_6_enq_ready = ~_writeQueue_fifo_6_full;
  wire              writeQueue_6_enq_valid;
  assign writeQueue_7_deq_valid = ~_writeQueue_fifo_7_empty;
  wire              exeResp_7_valid_0 = writeQueue_7_deq_valid;
  wire              writeQueue_dataOut_7_ffoByOther;
  wire [31:0]       writeQueue_dataOut_7_writeData_data;
  wire [31:0]       exeResp_7_bits_data_0 = writeQueue_7_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_7_writeData_mask;
  wire [3:0]        exeResp_7_bits_mask_0 = writeQueue_7_deq_bits_writeData_mask;
  wire [5:0]        writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_7_writeData_vd;
  wire [2:0]        writeQueue_dataOut_7_index;
  wire [5:0]        writeQueue_7_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_7_enq_bits_writeData_vd;
  wire [10:0]       writeQueue_dataIn_lo_7 = {writeQueue_7_enq_bits_writeData_groupCounter, writeQueue_7_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_7_enq_bits_writeData_data;
  wire [3:0]        writeQueue_7_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_14 = {writeQueue_7_enq_bits_writeData_data, writeQueue_7_enq_bits_writeData_mask};
  wire              writeQueue_7_enq_bits_ffoByOther;
  wire [47:0]       writeQueue_dataIn_hi_15 = {writeQueue_7_enq_bits_ffoByOther, writeQueue_dataIn_hi_14, writeQueue_dataIn_lo_7};
  wire [50:0]       writeQueue_dataIn_7 = {writeQueue_dataIn_hi_15, writeQueue_7_enq_bits_index};
  assign writeQueue_dataOut_7_index = _writeQueue_fifo_7_data_out[2:0];
  assign writeQueue_dataOut_7_writeData_vd = _writeQueue_fifo_7_data_out[7:3];
  assign writeQueue_dataOut_7_writeData_groupCounter = _writeQueue_fifo_7_data_out[13:8];
  assign writeQueue_dataOut_7_writeData_mask = _writeQueue_fifo_7_data_out[17:14];
  assign writeQueue_dataOut_7_writeData_data = _writeQueue_fifo_7_data_out[49:18];
  assign writeQueue_dataOut_7_ffoByOther = _writeQueue_fifo_7_data_out[50];
  wire              writeQueue_7_deq_bits_ffoByOther = writeQueue_dataOut_7_ffoByOther;
  assign writeQueue_7_deq_bits_writeData_data = writeQueue_dataOut_7_writeData_data;
  assign writeQueue_7_deq_bits_writeData_mask = writeQueue_dataOut_7_writeData_mask;
  wire [5:0]        writeQueue_7_deq_bits_writeData_groupCounter = writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]        writeQueue_7_deq_bits_writeData_vd = writeQueue_dataOut_7_writeData_vd;
  wire [2:0]        writeQueue_7_deq_bits_index = writeQueue_dataOut_7_index;
  wire              writeQueue_7_enq_ready = ~_writeQueue_fifo_7_full;
  wire              writeQueue_7_enq_valid;
  wire              dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]        exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter;
  wire              _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]        exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_1;
  wire              _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]        exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_2;
  wire              _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]        exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_3;
  wire              _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_4 = waiteStageDeqFire & WillWriteLane[4];
  assign writeQueue_4_enq_valid = _maskedWrite_out_4_valid | dataNotInShifter_readTypeWriteVrf_4;
  assign writeQueue_4_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_vd : 5'h0;
  assign writeQueue_4_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_groupCounter : _maskedWrite_out_4_bits_writeData_groupCounter;
  assign writeQueue_4_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_mask : _maskedWrite_out_4_bits_writeData_mask;
  assign writeQueue_4_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_data : _maskedWrite_out_4_bits_writeData_data;
  assign writeQueue_4_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_4 & _maskedWrite_out_4_bits_ffoByOther;
  wire [4:0]        exeResp_4_bits_vd_0 = instReg_vd + {1'h0, writeQueue_4_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_4_bits_offset_0 = writeQueue_4_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_4;
  wire              _dataNotInShifter_T_12 = exeResp_4_ready_0 & exeResp_4_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_4 = _dataNotInShifter_T_12 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_5 = waiteStageDeqFire & WillWriteLane[5];
  assign writeQueue_5_enq_valid = _maskedWrite_out_5_valid | dataNotInShifter_readTypeWriteVrf_5;
  assign writeQueue_5_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_vd : 5'h0;
  assign writeQueue_5_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_groupCounter : _maskedWrite_out_5_bits_writeData_groupCounter;
  assign writeQueue_5_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_mask : _maskedWrite_out_5_bits_writeData_mask;
  assign writeQueue_5_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_data : _maskedWrite_out_5_bits_writeData_data;
  assign writeQueue_5_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_5 & _maskedWrite_out_5_bits_ffoByOther;
  wire [4:0]        exeResp_5_bits_vd_0 = instReg_vd + {1'h0, writeQueue_5_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_5_bits_offset_0 = writeQueue_5_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_5;
  wire              _dataNotInShifter_T_15 = exeResp_5_ready_0 & exeResp_5_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_5 = _dataNotInShifter_T_15 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_6 = waiteStageDeqFire & WillWriteLane[6];
  assign writeQueue_6_enq_valid = _maskedWrite_out_6_valid | dataNotInShifter_readTypeWriteVrf_6;
  assign writeQueue_6_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_vd : 5'h0;
  assign writeQueue_6_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_groupCounter : _maskedWrite_out_6_bits_writeData_groupCounter;
  assign writeQueue_6_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_mask : _maskedWrite_out_6_bits_writeData_mask;
  assign writeQueue_6_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_data : _maskedWrite_out_6_bits_writeData_data;
  assign writeQueue_6_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_6 & _maskedWrite_out_6_bits_ffoByOther;
  wire [4:0]        exeResp_6_bits_vd_0 = instReg_vd + {1'h0, writeQueue_6_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_6_bits_offset_0 = writeQueue_6_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_6;
  wire              _dataNotInShifter_T_18 = exeResp_6_ready_0 & exeResp_6_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_6 = _dataNotInShifter_T_18 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_7 = waiteStageDeqFire & WillWriteLane[7];
  assign writeQueue_7_enq_valid = _maskedWrite_out_7_valid | dataNotInShifter_readTypeWriteVrf_7;
  assign writeQueue_7_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_vd : 5'h0;
  assign writeQueue_7_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_groupCounter : _maskedWrite_out_7_bits_writeData_groupCounter;
  assign writeQueue_7_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_mask : _maskedWrite_out_7_bits_writeData_mask;
  assign writeQueue_7_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_data : _maskedWrite_out_7_bits_writeData_data;
  assign writeQueue_7_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_7 & _maskedWrite_out_7_bits_ffoByOther;
  wire [4:0]        exeResp_7_bits_vd_0 = instReg_vd + {1'h0, writeQueue_7_deq_bits_writeData_groupCounter[5:2]};
  wire [1:0]        exeResp_7_bits_offset_0 = writeQueue_7_deq_bits_writeData_groupCounter[1:0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_7;
  wire              _dataNotInShifter_T_21 = exeResp_7_ready_0 & exeResp_7_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_7 = _dataNotInShifter_T_21 ? 3'h1 : 3'h7;
  wire              dataNotInShifter =
    dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0 & dataNotInShifter_writeTokenCounter_4 == 3'h0
    & dataNotInShifter_writeTokenCounter_5 == 3'h0 & dataNotInShifter_writeTokenCounter_6 == 3'h0 & dataNotInShifter_writeTokenCounter_7 == 3'h0;
  assign waiteStageDeqReady =
    (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready)
    & (~(WillWriteLane[4]) | writeQueue_4_enq_ready) & (~(WillWriteLane[5]) | writeQueue_5_enq_ready) & (~(WillWriteLane[6]) | writeQueue_6_enq_ready) & (~(WillWriteLane[7]) | writeQueue_7_enq_ready);
  reg               waiteLastRequest;
  reg               waitQueueClear;
  wire              lastReportValid =
    waitQueueClear & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid | writeQueue_4_deq_valid | writeQueue_5_deq_valid | writeQueue_6_deq_valid | writeQueue_7_deq_valid)
    & dataNotInShifter;
  wire              executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire              executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire              invalidEnq = instReq_valid & instReq_bits_vl == 11'h0 & ~enqMvRD;
  wire [7:0]        _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]       gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 3'h0;
      gatherOffset <= 2'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_orderReduce <= 1'h0;
      instReg_decodeResult_floatMul <= 1'h0;
      instReg_decodeResult_fpExecutionType <= 2'h0;
      instReg_decodeResult_float <= 1'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 11'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 5'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_0_bits_fpReduceValid <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_1_bits_fpReduceValid <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_2_bits_fpReduceValid <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      exeReqReg_3_bits_fpReduceValid <= 1'h0;
      exeReqReg_4_valid <= 1'h0;
      exeReqReg_4_bits_source1 <= 32'h0;
      exeReqReg_4_bits_source2 <= 32'h0;
      exeReqReg_4_bits_index <= 3'h0;
      exeReqReg_4_bits_ffo <= 1'h0;
      exeReqReg_4_bits_fpReduceValid <= 1'h0;
      exeReqReg_5_valid <= 1'h0;
      exeReqReg_5_bits_source1 <= 32'h0;
      exeReqReg_5_bits_source2 <= 32'h0;
      exeReqReg_5_bits_index <= 3'h0;
      exeReqReg_5_bits_ffo <= 1'h0;
      exeReqReg_5_bits_fpReduceValid <= 1'h0;
      exeReqReg_6_valid <= 1'h0;
      exeReqReg_6_bits_source1 <= 32'h0;
      exeReqReg_6_bits_source2 <= 32'h0;
      exeReqReg_6_bits_index <= 3'h0;
      exeReqReg_6_bits_ffo <= 1'h0;
      exeReqReg_6_bits_fpReduceValid <= 1'h0;
      exeReqReg_7_valid <= 1'h0;
      exeReqReg_7_bits_source1 <= 32'h0;
      exeReqReg_7_bits_source2 <= 32'h0;
      exeReqReg_7_bits_index <= 3'h0;
      exeReqReg_7_bits_ffo <= 1'h0;
      exeReqReg_7_bits_fpReduceValid <= 1'h0;
      requestCounter <= 6'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 8'h0;
      readIssueStageState_needRead <= 8'h0;
      readIssueStageState_elementValid <= 8'h0;
      readIssueStageState_replaceVs1 <= 8'h0;
      readIssueStageState_readOffset <= 16'h0;
      readIssueStageState_accessLane_0 <= 3'h0;
      readIssueStageState_accessLane_1 <= 3'h0;
      readIssueStageState_accessLane_2 <= 3'h0;
      readIssueStageState_accessLane_3 <= 3'h0;
      readIssueStageState_accessLane_4 <= 3'h0;
      readIssueStageState_accessLane_5 <= 3'h0;
      readIssueStageState_accessLane_6 <= 3'h0;
      readIssueStageState_accessLane_7 <= 3'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_vsGrowth_4 <= 3'h0;
      readIssueStageState_vsGrowth_5 <= 3'h0;
      readIssueStageState_vsGrowth_6 <= 3'h0;
      readIssueStageState_vsGrowth_7 <= 3'h0;
      readIssueStageState_executeGroup <= 8'h0;
      readIssueStageState_readDataOffset <= 16'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      tokenCheck_counter_4 <= 4'h0;
      tokenCheck_counter_5 <= 4'h0;
      tokenCheck_counter_6 <= 4'h0;
      tokenCheck_counter_7 <= 4'h0;
      reorderQueueAllocate_counter <= 5'h0;
      reorderQueueAllocate_counterWillUpdate <= 5'h0;
      reorderQueueAllocate_counter_1 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 5'h0;
      reorderQueueAllocate_counter_2 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 5'h0;
      reorderQueueAllocate_counter_3 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 5'h0;
      reorderQueueAllocate_counter_4 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_4 <= 5'h0;
      reorderQueueAllocate_counter_5 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_5 <= 5'h0;
      reorderQueueAllocate_counter_6 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_6 <= 5'h0;
      reorderQueueAllocate_counter_7 <= 5'h0;
      reorderQueueAllocate_counterWillUpdate_7 <= 5'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 4'h0;
      reorderStageState_1 <= 4'h0;
      reorderStageState_2 <= 4'h0;
      reorderStageState_3 <= 4'h0;
      reorderStageState_4 <= 4'h0;
      reorderStageState_5 <= 4'h0;
      reorderStageState_6 <= 4'h0;
      reorderStageState_7 <= 4'h0;
      reorderStageNeed_0 <= 4'h0;
      reorderStageNeed_1 <= 4'h0;
      reorderStageNeed_2 <= 4'h0;
      reorderStageNeed_3 <= 4'h0;
      reorderStageNeed_4 <= 4'h0;
      reorderStageNeed_5 <= 4'h0;
      reorderStageNeed_6 <= 4'h0;
      reorderStageNeed_7 <= 4'h0;
      waiteReadDataPipeReg_executeGroup <= 8'h0;
      waiteReadDataPipeReg_sourceValid <= 8'h0;
      waiteReadDataPipeReg_replaceVs1 <= 8'h0;
      waiteReadDataPipeReg_needRead <= 8'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadData_4 <= 32'h0;
      waiteReadData_5 <= 32'h0;
      waiteReadData_6 <= 32'h0;
      waiteReadData_7 <= 32'h0;
      waiteReadSate <= 8'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      dataNotInShifter_writeTokenCounter_4 <= 3'h0;
      dataNotInShifter_writeTokenCounter_5 <= 3'h0;
      dataNotInShifter_writeTokenCounter_6 <= 3'h0;
      dataNotInShifter_writeTokenCounter_7 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_88 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_89;
      automatic logic _GEN_90 = source1Change & viotaCounterAdd;
      _GEN_89 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h0)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h0)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h0)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h0)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h1)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h1)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h1)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h1)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h1)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h1)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h1)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h1)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h2)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h2)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h2)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h2)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h2)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h2)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h2)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h2)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & (&v0UpdateVec_4_bits_offset))
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & (&v0UpdateVec_5_bits_offset))
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & (&v0UpdateVec_6_bits_offset))
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & (&v0UpdateVec_7_bits_offset))
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_7_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_88 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_orderReduce <= instReq_bits_decodeResult_orderReduce;
        instReg_decodeResult_floatMul <= instReq_bits_decodeResult_floatMul;
        instReg_decodeResult_fpExecutionType <= instReq_bits_decodeResult_fpExecutionType;
        instReg_decodeResult_float <= instReq_bits_decodeResult_float;
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_88)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_90 & (readTokenRelease_0 | ~_GEN_89 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_90 & (_tokenCheck_T | ~_GEN_89 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_89 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_90)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 5'h1;
      else if (_GEN_89)
        readVS1Reg_readIndex <= 5'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
        exeReqReg_0_bits_fpReduceValid <= exeRequestQueue_0_deq_bits_fpReduceValid;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
        exeReqReg_1_bits_fpReduceValid <= exeRequestQueue_1_deq_bits_fpReduceValid;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
        exeReqReg_2_bits_fpReduceValid <= exeRequestQueue_2_deq_bits_fpReduceValid;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
        exeReqReg_3_bits_fpReduceValid <= exeRequestQueue_3_deq_bits_fpReduceValid;
      end
      if (tokenIO_4_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_4_valid <= tokenIO_4_maskRequestRelease_0 & ~viota;
      if (tokenIO_4_maskRequestRelease_0) begin
        exeReqReg_4_bits_source1 <= exeRequestQueue_4_deq_bits_source1;
        exeReqReg_4_bits_source2 <= exeRequestQueue_4_deq_bits_source2;
        exeReqReg_4_bits_index <= exeRequestQueue_4_deq_bits_index;
        exeReqReg_4_bits_ffo <= exeRequestQueue_4_deq_bits_ffo;
        exeReqReg_4_bits_fpReduceValid <= exeRequestQueue_4_deq_bits_fpReduceValid;
      end
      if (tokenIO_5_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_5_valid <= tokenIO_5_maskRequestRelease_0 & ~viota;
      if (tokenIO_5_maskRequestRelease_0) begin
        exeReqReg_5_bits_source1 <= exeRequestQueue_5_deq_bits_source1;
        exeReqReg_5_bits_source2 <= exeRequestQueue_5_deq_bits_source2;
        exeReqReg_5_bits_index <= exeRequestQueue_5_deq_bits_index;
        exeReqReg_5_bits_ffo <= exeRequestQueue_5_deq_bits_ffo;
        exeReqReg_5_bits_fpReduceValid <= exeRequestQueue_5_deq_bits_fpReduceValid;
      end
      if (tokenIO_6_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_6_valid <= tokenIO_6_maskRequestRelease_0 & ~viota;
      if (tokenIO_6_maskRequestRelease_0) begin
        exeReqReg_6_bits_source1 <= exeRequestQueue_6_deq_bits_source1;
        exeReqReg_6_bits_source2 <= exeRequestQueue_6_deq_bits_source2;
        exeReqReg_6_bits_index <= exeRequestQueue_6_deq_bits_index;
        exeReqReg_6_bits_ffo <= exeRequestQueue_6_deq_bits_ffo;
        exeReqReg_6_bits_fpReduceValid <= exeRequestQueue_6_deq_bits_fpReduceValid;
      end
      if (tokenIO_7_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_7_valid <= tokenIO_7_maskRequestRelease_0 & ~viota;
      if (tokenIO_7_maskRequestRelease_0) begin
        exeReqReg_7_bits_source1 <= exeRequestQueue_7_deq_bits_source1;
        exeReqReg_7_bits_source2 <= exeRequestQueue_7_deq_bits_source2;
        exeReqReg_7_bits_index <= exeRequestQueue_7_deq_bits_index;
        exeReqReg_7_bits_ffo <= exeRequestQueue_7_deq_bits_ffo;
        exeReqReg_7_bits_fpReduceValid <= exeRequestQueue_7_deq_bits_fpReduceValid;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 6'h0 : requestCounter + 6'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 8'h0;
        readIssueStageState_needRead <= _GEN_78 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_78 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 8'h0;
        readIssueStageState_readOffset <= _GEN_78 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[2:0];
        readIssueStageState_accessLane_1 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[5:3];
        readIssueStageState_accessLane_2 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[8:6];
        readIssueStageState_accessLane_3 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[11:9];
        readIssueStageState_accessLane_4 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_4 : accessLaneSelect[14:12];
        readIssueStageState_accessLane_5 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_5 : accessLaneSelect[17:15];
        readIssueStageState_accessLane_6 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_6 : accessLaneSelect[20:18];
        readIssueStageState_accessLane_7 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_accessLane_7 : accessLaneSelect[23:21];
        readIssueStageState_vsGrowth_0 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_vsGrowth_4 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_4 : growthSelect[14:12];
        readIssueStageState_vsGrowth_5 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_5 : growthSelect[17:15];
        readIssueStageState_vsGrowth_6 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_6 : growthSelect[20:18];
        readIssueStageState_vsGrowth_7 <= _GEN_78 ? _slideAddressGen_indexDeq_bits_vsGrowth_7 : growthSelect[23:21];
        readIssueStageState_executeGroup <= _GEN_78 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_78 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_78 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (pipeReadFire_4 ^ readTokenRelease_4)
        tokenCheck_counter_4 <= tokenCheck_counter_4 + tokenCheck_counterChange_4;
      if (pipeReadFire_5 ^ readTokenRelease_5)
        tokenCheck_counter_5 <= tokenCheck_counter_5 + tokenCheck_counterChange_5;
      if (pipeReadFire_6 ^ readTokenRelease_6)
        tokenCheck_counter_6 <= tokenCheck_counter_6 + tokenCheck_counterChange_6;
      if (pipeReadFire_7 ^ readTokenRelease_7)
        tokenCheck_counter_7 <= tokenCheck_counter_7 + tokenCheck_counterChange_7;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 5'h8;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 5'h8;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 5'h8;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 5'h8;
      end
      if (reorderQueueAllocate_release_4 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_4 <= reorderQueueAllocate_counterUpdate_4;
        reorderQueueAllocate_counterWillUpdate_4 <= reorderQueueAllocate_counterUpdate_4 + 5'h8;
      end
      if (reorderQueueAllocate_release_5 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_5 <= reorderQueueAllocate_counterUpdate_5;
        reorderQueueAllocate_counterWillUpdate_5 <= reorderQueueAllocate_counterUpdate_5 + 5'h8;
      end
      if (reorderQueueAllocate_release_6 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_6 <= reorderQueueAllocate_counterUpdate_6;
        reorderQueueAllocate_counterWillUpdate_6 <= reorderQueueAllocate_counterUpdate_6 + 5'h8;
      end
      if (reorderQueueAllocate_release_7 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_7 <= reorderQueueAllocate_counterUpdate_7;
        reorderQueueAllocate_counterWillUpdate_7 <= reorderQueueAllocate_counterUpdate_7 + 5'h8;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 4'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 4'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 4'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 4'h0;
      if (_write1HPipe_4_T & readType)
        reorderStageState_4 <= reorderStageState_4 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_4 <= 4'h0;
      if (_write1HPipe_5_T & readType)
        reorderStageState_5 <= reorderStageState_5 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_5 <= 4'h0;
      if (_write1HPipe_6_T & readType)
        reorderStageState_6 <= reorderStageState_6 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_6 <= 4'h0;
      if (_write1HPipe_7_T & readType)
        reorderStageState_7 <= reorderStageState_7 + 4'h1;
      else if (reorderStageEnqFire)
        reorderStageState_7 <= 4'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
        reorderStageNeed_4 <= accessCountQueue_deq_bits_4;
        reorderStageNeed_5 <= accessCountQueue_deq_bits_5;
        reorderStageNeed_6 <= accessCountQueue_deq_bits_6;
        reorderStageNeed_7 <= accessCountQueue_deq_bits_7;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (readTokenRelease_4)
        waiteReadData_4 <= readData_readDataQueue_4_deq_bits;
      if (readTokenRelease_5)
        waiteReadData_5 <= readData_readDataQueue_5_deq_bits;
      if (readTokenRelease_6)
        waiteReadData_6 <= readData_readDataQueue_6_deq_bits;
      if (readTokenRelease_7)
        waiteReadData_7 <= readData_readDataQueue_7_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 8'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      if (_dataNotInShifter_T_12 ^ writeRelease_4)
        dataNotInShifter_writeTokenCounter_4 <= dataNotInShifter_writeTokenCounter_4 + dataNotInShifter_writeTokenChange_4;
      if (_dataNotInShifter_T_15 ^ writeRelease_5)
        dataNotInShifter_writeTokenCounter_5 <= dataNotInShifter_writeTokenCounter_5 + dataNotInShifter_writeTokenChange_5;
      if (_dataNotInShifter_T_18 ^ writeRelease_6)
        dataNotInShifter_writeTokenCounter_6 <= dataNotInShifter_writeTokenCounter_6 + dataNotInShifter_writeTokenChange_6;
      if (_dataNotInShifter_T_21 ^ writeRelease_7)
        dataNotInShifter_writeTokenCounter_7 <= dataNotInShifter_writeTokenCounter_7 + dataNotInShifter_writeTokenChange_7;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:75];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h4C; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[7'h0];
        v0_1 = _RANDOM[7'h1];
        v0_2 = _RANDOM[7'h2];
        v0_3 = _RANDOM[7'h3];
        v0_4 = _RANDOM[7'h4];
        v0_5 = _RANDOM[7'h5];
        v0_6 = _RANDOM[7'h6];
        v0_7 = _RANDOM[7'h7];
        v0_8 = _RANDOM[7'h8];
        v0_9 = _RANDOM[7'h9];
        v0_10 = _RANDOM[7'hA];
        v0_11 = _RANDOM[7'hB];
        v0_12 = _RANDOM[7'hC];
        v0_13 = _RANDOM[7'hD];
        v0_14 = _RANDOM[7'hE];
        v0_15 = _RANDOM[7'hF];
        v0_16 = _RANDOM[7'h10];
        v0_17 = _RANDOM[7'h11];
        v0_18 = _RANDOM[7'h12];
        v0_19 = _RANDOM[7'h13];
        v0_20 = _RANDOM[7'h14];
        v0_21 = _RANDOM[7'h15];
        v0_22 = _RANDOM[7'h16];
        v0_23 = _RANDOM[7'h17];
        v0_24 = _RANDOM[7'h18];
        v0_25 = _RANDOM[7'h19];
        v0_26 = _RANDOM[7'h1A];
        v0_27 = _RANDOM[7'h1B];
        v0_28 = _RANDOM[7'h1C];
        v0_29 = _RANDOM[7'h1D];
        v0_30 = _RANDOM[7'h1E];
        v0_31 = _RANDOM[7'h1F];
        gatherReadState = _RANDOM[7'h20][1:0];
        gatherDatOffset = _RANDOM[7'h20][3:2];
        gatherLane = _RANDOM[7'h20][6:4];
        gatherOffset = _RANDOM[7'h20][8:7];
        gatherGrowth = _RANDOM[7'h20][11:9];
        instReg_instructionIndex = _RANDOM[7'h20][14:12];
        instReg_decodeResult_orderReduce = _RANDOM[7'h20][15];
        instReg_decodeResult_floatMul = _RANDOM[7'h20][16];
        instReg_decodeResult_fpExecutionType = _RANDOM[7'h20][18:17];
        instReg_decodeResult_float = _RANDOM[7'h20][19];
        instReg_decodeResult_specialSlot = _RANDOM[7'h20][20];
        instReg_decodeResult_topUop = _RANDOM[7'h20][25:21];
        instReg_decodeResult_popCount = _RANDOM[7'h20][26];
        instReg_decodeResult_ffo = _RANDOM[7'h20][27];
        instReg_decodeResult_average = _RANDOM[7'h20][28];
        instReg_decodeResult_reverse = _RANDOM[7'h20][29];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[7'h20][30];
        instReg_decodeResult_scheduler = _RANDOM[7'h20][31];
        instReg_decodeResult_sReadVD = _RANDOM[7'h21][0];
        instReg_decodeResult_vtype = _RANDOM[7'h21][1];
        instReg_decodeResult_sWrite = _RANDOM[7'h21][2];
        instReg_decodeResult_crossRead = _RANDOM[7'h21][3];
        instReg_decodeResult_crossWrite = _RANDOM[7'h21][4];
        instReg_decodeResult_maskUnit = _RANDOM[7'h21][5];
        instReg_decodeResult_special = _RANDOM[7'h21][6];
        instReg_decodeResult_saturate = _RANDOM[7'h21][7];
        instReg_decodeResult_vwmacc = _RANDOM[7'h21][8];
        instReg_decodeResult_readOnly = _RANDOM[7'h21][9];
        instReg_decodeResult_maskSource = _RANDOM[7'h21][10];
        instReg_decodeResult_maskDestination = _RANDOM[7'h21][11];
        instReg_decodeResult_maskLogic = _RANDOM[7'h21][12];
        instReg_decodeResult_uop = _RANDOM[7'h21][16:13];
        instReg_decodeResult_iota = _RANDOM[7'h21][17];
        instReg_decodeResult_mv = _RANDOM[7'h21][18];
        instReg_decodeResult_extend = _RANDOM[7'h21][19];
        instReg_decodeResult_unOrderWrite = _RANDOM[7'h21][20];
        instReg_decodeResult_compress = _RANDOM[7'h21][21];
        instReg_decodeResult_gather16 = _RANDOM[7'h21][22];
        instReg_decodeResult_gather = _RANDOM[7'h21][23];
        instReg_decodeResult_slid = _RANDOM[7'h21][24];
        instReg_decodeResult_targetRd = _RANDOM[7'h21][25];
        instReg_decodeResult_widenReduce = _RANDOM[7'h21][26];
        instReg_decodeResult_red = _RANDOM[7'h21][27];
        instReg_decodeResult_nr = _RANDOM[7'h21][28];
        instReg_decodeResult_itype = _RANDOM[7'h21][29];
        instReg_decodeResult_unsigned1 = _RANDOM[7'h21][30];
        instReg_decodeResult_unsigned0 = _RANDOM[7'h21][31];
        instReg_decodeResult_other = _RANDOM[7'h22][0];
        instReg_decodeResult_multiCycle = _RANDOM[7'h22][1];
        instReg_decodeResult_divider = _RANDOM[7'h22][2];
        instReg_decodeResult_multiplier = _RANDOM[7'h22][3];
        instReg_decodeResult_shift = _RANDOM[7'h22][4];
        instReg_decodeResult_adder = _RANDOM[7'h22][5];
        instReg_decodeResult_logic = _RANDOM[7'h22][6];
        instReg_readFromScala = {_RANDOM[7'h22][31:7], _RANDOM[7'h23][6:0]};
        instReg_sew = _RANDOM[7'h23][8:7];
        instReg_vlmul = _RANDOM[7'h23][11:9];
        instReg_maskType = _RANDOM[7'h23][12];
        instReg_vxrm = _RANDOM[7'h23][15:13];
        instReg_vs2 = _RANDOM[7'h23][20:16];
        instReg_vs1 = _RANDOM[7'h23][25:21];
        instReg_vd = _RANDOM[7'h23][30:26];
        instReg_vl = {_RANDOM[7'h23][31], _RANDOM[7'h24][9:0]};
        instVlValid = _RANDOM[7'h24][10];
        readVS1Reg_dataValid = _RANDOM[7'h24][11];
        readVS1Reg_requestSend = _RANDOM[7'h24][12];
        readVS1Reg_sendToExecution = _RANDOM[7'h24][13];
        readVS1Reg_data = {_RANDOM[7'h24][31:14], _RANDOM[7'h25][13:0]};
        readVS1Reg_readIndex = _RANDOM[7'h25][18:14];
        exeReqReg_0_valid = _RANDOM[7'h25][27];
        exeReqReg_0_bits_source1 = {_RANDOM[7'h25][31:28], _RANDOM[7'h26][27:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[7'h26][31:28], _RANDOM[7'h27][27:0]};
        exeReqReg_0_bits_index = _RANDOM[7'h27][30:28];
        exeReqReg_0_bits_ffo = _RANDOM[7'h27][31];
        exeReqReg_0_bits_fpReduceValid = _RANDOM[7'h28][0];
        exeReqReg_1_valid = _RANDOM[7'h28][1];
        exeReqReg_1_bits_source1 = {_RANDOM[7'h28][31:2], _RANDOM[7'h29][1:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[7'h29][31:2], _RANDOM[7'h2A][1:0]};
        exeReqReg_1_bits_index = _RANDOM[7'h2A][4:2];
        exeReqReg_1_bits_ffo = _RANDOM[7'h2A][5];
        exeReqReg_1_bits_fpReduceValid = _RANDOM[7'h2A][6];
        exeReqReg_2_valid = _RANDOM[7'h2A][7];
        exeReqReg_2_bits_source1 = {_RANDOM[7'h2A][31:8], _RANDOM[7'h2B][7:0]};
        exeReqReg_2_bits_source2 = {_RANDOM[7'h2B][31:8], _RANDOM[7'h2C][7:0]};
        exeReqReg_2_bits_index = _RANDOM[7'h2C][10:8];
        exeReqReg_2_bits_ffo = _RANDOM[7'h2C][11];
        exeReqReg_2_bits_fpReduceValid = _RANDOM[7'h2C][12];
        exeReqReg_3_valid = _RANDOM[7'h2C][13];
        exeReqReg_3_bits_source1 = {_RANDOM[7'h2C][31:14], _RANDOM[7'h2D][13:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[7'h2D][31:14], _RANDOM[7'h2E][13:0]};
        exeReqReg_3_bits_index = _RANDOM[7'h2E][16:14];
        exeReqReg_3_bits_ffo = _RANDOM[7'h2E][17];
        exeReqReg_3_bits_fpReduceValid = _RANDOM[7'h2E][18];
        exeReqReg_4_valid = _RANDOM[7'h2E][19];
        exeReqReg_4_bits_source1 = {_RANDOM[7'h2E][31:20], _RANDOM[7'h2F][19:0]};
        exeReqReg_4_bits_source2 = {_RANDOM[7'h2F][31:20], _RANDOM[7'h30][19:0]};
        exeReqReg_4_bits_index = _RANDOM[7'h30][22:20];
        exeReqReg_4_bits_ffo = _RANDOM[7'h30][23];
        exeReqReg_4_bits_fpReduceValid = _RANDOM[7'h30][24];
        exeReqReg_5_valid = _RANDOM[7'h30][25];
        exeReqReg_5_bits_source1 = {_RANDOM[7'h30][31:26], _RANDOM[7'h31][25:0]};
        exeReqReg_5_bits_source2 = {_RANDOM[7'h31][31:26], _RANDOM[7'h32][25:0]};
        exeReqReg_5_bits_index = _RANDOM[7'h32][28:26];
        exeReqReg_5_bits_ffo = _RANDOM[7'h32][29];
        exeReqReg_5_bits_fpReduceValid = _RANDOM[7'h32][30];
        exeReqReg_6_valid = _RANDOM[7'h32][31];
        exeReqReg_6_bits_source1 = _RANDOM[7'h33];
        exeReqReg_6_bits_source2 = _RANDOM[7'h34];
        exeReqReg_6_bits_index = _RANDOM[7'h35][2:0];
        exeReqReg_6_bits_ffo = _RANDOM[7'h35][3];
        exeReqReg_6_bits_fpReduceValid = _RANDOM[7'h35][4];
        exeReqReg_7_valid = _RANDOM[7'h35][5];
        exeReqReg_7_bits_source1 = {_RANDOM[7'h35][31:6], _RANDOM[7'h36][5:0]};
        exeReqReg_7_bits_source2 = {_RANDOM[7'h36][31:6], _RANDOM[7'h37][5:0]};
        exeReqReg_7_bits_index = _RANDOM[7'h37][8:6];
        exeReqReg_7_bits_ffo = _RANDOM[7'h37][9];
        exeReqReg_7_bits_fpReduceValid = _RANDOM[7'h37][10];
        requestCounter = _RANDOM[7'h37][16:11];
        executeIndex = _RANDOM[7'h37][18:17];
        readIssueStageState_groupReadState = _RANDOM[7'h37][26:19];
        readIssueStageState_needRead = {_RANDOM[7'h37][31:27], _RANDOM[7'h38][2:0]};
        readIssueStageState_elementValid = _RANDOM[7'h38][10:3];
        readIssueStageState_replaceVs1 = _RANDOM[7'h38][18:11];
        readIssueStageState_readOffset = {_RANDOM[7'h38][31:19], _RANDOM[7'h39][2:0]};
        readIssueStageState_accessLane_0 = _RANDOM[7'h39][5:3];
        readIssueStageState_accessLane_1 = _RANDOM[7'h39][8:6];
        readIssueStageState_accessLane_2 = _RANDOM[7'h39][11:9];
        readIssueStageState_accessLane_3 = _RANDOM[7'h39][14:12];
        readIssueStageState_accessLane_4 = _RANDOM[7'h39][17:15];
        readIssueStageState_accessLane_5 = _RANDOM[7'h39][20:18];
        readIssueStageState_accessLane_6 = _RANDOM[7'h39][23:21];
        readIssueStageState_accessLane_7 = _RANDOM[7'h39][26:24];
        readIssueStageState_vsGrowth_0 = _RANDOM[7'h39][29:27];
        readIssueStageState_vsGrowth_1 = {_RANDOM[7'h39][31:30], _RANDOM[7'h3A][0]};
        readIssueStageState_vsGrowth_2 = _RANDOM[7'h3A][3:1];
        readIssueStageState_vsGrowth_3 = _RANDOM[7'h3A][6:4];
        readIssueStageState_vsGrowth_4 = _RANDOM[7'h3A][9:7];
        readIssueStageState_vsGrowth_5 = _RANDOM[7'h3A][12:10];
        readIssueStageState_vsGrowth_6 = _RANDOM[7'h3A][15:13];
        readIssueStageState_vsGrowth_7 = _RANDOM[7'h3A][18:16];
        readIssueStageState_executeGroup = _RANDOM[7'h3A][26:19];
        readIssueStageState_readDataOffset = {_RANDOM[7'h3A][31:27], _RANDOM[7'h3B][10:0]};
        readIssueStageState_last = _RANDOM[7'h3B][11];
        readIssueStageValid = _RANDOM[7'h3B][12];
        tokenCheck_counter = _RANDOM[7'h3B][16:13];
        tokenCheck_counter_1 = _RANDOM[7'h3B][20:17];
        tokenCheck_counter_2 = _RANDOM[7'h3B][24:21];
        tokenCheck_counter_3 = _RANDOM[7'h3B][28:25];
        tokenCheck_counter_4 = {_RANDOM[7'h3B][31:29], _RANDOM[7'h3C][0]};
        tokenCheck_counter_5 = _RANDOM[7'h3C][4:1];
        tokenCheck_counter_6 = _RANDOM[7'h3C][8:5];
        tokenCheck_counter_7 = _RANDOM[7'h3C][12:9];
        reorderQueueAllocate_counter = _RANDOM[7'h3C][17:13];
        reorderQueueAllocate_counterWillUpdate = _RANDOM[7'h3C][22:18];
        reorderQueueAllocate_counter_1 = _RANDOM[7'h3C][27:23];
        reorderQueueAllocate_counterWillUpdate_1 = {_RANDOM[7'h3C][31:28], _RANDOM[7'h3D][0]};
        reorderQueueAllocate_counter_2 = _RANDOM[7'h3D][5:1];
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[7'h3D][10:6];
        reorderQueueAllocate_counter_3 = _RANDOM[7'h3D][15:11];
        reorderQueueAllocate_counterWillUpdate_3 = _RANDOM[7'h3D][20:16];
        reorderQueueAllocate_counter_4 = _RANDOM[7'h3D][25:21];
        reorderQueueAllocate_counterWillUpdate_4 = _RANDOM[7'h3D][30:26];
        reorderQueueAllocate_counter_5 = {_RANDOM[7'h3D][31], _RANDOM[7'h3E][3:0]};
        reorderQueueAllocate_counterWillUpdate_5 = _RANDOM[7'h3E][8:4];
        reorderQueueAllocate_counter_6 = _RANDOM[7'h3E][13:9];
        reorderQueueAllocate_counterWillUpdate_6 = _RANDOM[7'h3E][18:14];
        reorderQueueAllocate_counter_7 = _RANDOM[7'h3E][23:19];
        reorderQueueAllocate_counterWillUpdate_7 = _RANDOM[7'h3E][28:24];
        reorderStageValid = _RANDOM[7'h3E][29];
        reorderStageState_0 = {_RANDOM[7'h3E][31:30], _RANDOM[7'h3F][1:0]};
        reorderStageState_1 = _RANDOM[7'h3F][5:2];
        reorderStageState_2 = _RANDOM[7'h3F][9:6];
        reorderStageState_3 = _RANDOM[7'h3F][13:10];
        reorderStageState_4 = _RANDOM[7'h3F][17:14];
        reorderStageState_5 = _RANDOM[7'h3F][21:18];
        reorderStageState_6 = _RANDOM[7'h3F][25:22];
        reorderStageState_7 = _RANDOM[7'h3F][29:26];
        reorderStageNeed_0 = {_RANDOM[7'h3F][31:30], _RANDOM[7'h40][1:0]};
        reorderStageNeed_1 = _RANDOM[7'h40][5:2];
        reorderStageNeed_2 = _RANDOM[7'h40][9:6];
        reorderStageNeed_3 = _RANDOM[7'h40][13:10];
        reorderStageNeed_4 = _RANDOM[7'h40][17:14];
        reorderStageNeed_5 = _RANDOM[7'h40][21:18];
        reorderStageNeed_6 = _RANDOM[7'h40][25:22];
        reorderStageNeed_7 = _RANDOM[7'h40][29:26];
        waiteReadDataPipeReg_executeGroup = {_RANDOM[7'h40][31:30], _RANDOM[7'h41][5:0]};
        waiteReadDataPipeReg_sourceValid = _RANDOM[7'h41][13:6];
        waiteReadDataPipeReg_replaceVs1 = _RANDOM[7'h41][21:14];
        waiteReadDataPipeReg_needRead = _RANDOM[7'h41][29:22];
        waiteReadDataPipeReg_last = _RANDOM[7'h41][30];
        waiteReadData_0 = {_RANDOM[7'h41][31], _RANDOM[7'h42][30:0]};
        waiteReadData_1 = {_RANDOM[7'h42][31], _RANDOM[7'h43][30:0]};
        waiteReadData_2 = {_RANDOM[7'h43][31], _RANDOM[7'h44][30:0]};
        waiteReadData_3 = {_RANDOM[7'h44][31], _RANDOM[7'h45][30:0]};
        waiteReadData_4 = {_RANDOM[7'h45][31], _RANDOM[7'h46][30:0]};
        waiteReadData_5 = {_RANDOM[7'h46][31], _RANDOM[7'h47][30:0]};
        waiteReadData_6 = {_RANDOM[7'h47][31], _RANDOM[7'h48][30:0]};
        waiteReadData_7 = {_RANDOM[7'h48][31], _RANDOM[7'h49][30:0]};
        waiteReadSate = {_RANDOM[7'h49][31], _RANDOM[7'h4A][6:0]};
        waiteReadStageValid = _RANDOM[7'h4A][7];
        dataNotInShifter_writeTokenCounter = _RANDOM[7'h4A][10:8];
        dataNotInShifter_writeTokenCounter_1 = _RANDOM[7'h4A][13:11];
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[7'h4A][16:14];
        dataNotInShifter_writeTokenCounter_3 = _RANDOM[7'h4A][19:17];
        dataNotInShifter_writeTokenCounter_4 = _RANDOM[7'h4A][22:20];
        dataNotInShifter_writeTokenCounter_5 = _RANDOM[7'h4A][25:23];
        dataNotInShifter_writeTokenCounter_6 = _RANDOM[7'h4A][28:26];
        dataNotInShifter_writeTokenCounter_7 = _RANDOM[7'h4A][31:29];
        waiteLastRequest = _RANDOM[7'h4B][0];
        waitQueueClear = _RANDOM[7'h4B][1];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire              exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire              exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire              exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire              exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire              exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire              exeRequestQueue_4_empty;
  assign exeRequestQueue_4_empty = _exeRequestQueue_queue_fifo_4_empty;
  wire              exeRequestQueue_4_full;
  assign exeRequestQueue_4_full = _exeRequestQueue_queue_fifo_4_full;
  wire              exeRequestQueue_5_empty;
  assign exeRequestQueue_5_empty = _exeRequestQueue_queue_fifo_5_empty;
  wire              exeRequestQueue_5_full;
  assign exeRequestQueue_5_full = _exeRequestQueue_queue_fifo_5_full;
  wire              exeRequestQueue_6_empty;
  assign exeRequestQueue_6_empty = _exeRequestQueue_queue_fifo_6_empty;
  wire              exeRequestQueue_6_full;
  assign exeRequestQueue_6_full = _exeRequestQueue_queue_fifo_6_full;
  wire              exeRequestQueue_7_empty;
  assign exeRequestQueue_7_empty = _exeRequestQueue_queue_fifo_7_empty;
  wire              exeRequestQueue_7_full;
  assign exeRequestQueue_7_full = _exeRequestQueue_queue_fifo_7_full;
  wire              accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire              accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire              readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire              readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire              compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire              reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire              reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire              reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire              reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire              reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire              reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire              reorderQueueVec_4_empty;
  assign reorderQueueVec_4_empty = _reorderQueueVec_fifo_4_empty;
  wire              reorderQueueVec_4_full;
  assign reorderQueueVec_4_full = _reorderQueueVec_fifo_4_full;
  wire              reorderQueueVec_5_empty;
  assign reorderQueueVec_5_empty = _reorderQueueVec_fifo_5_empty;
  wire              reorderQueueVec_5_full;
  assign reorderQueueVec_5_full = _reorderQueueVec_fifo_5_full;
  wire              reorderQueueVec_6_empty;
  assign reorderQueueVec_6_empty = _reorderQueueVec_fifo_6_empty;
  wire              reorderQueueVec_6_full;
  assign reorderQueueVec_6_full = _reorderQueueVec_fifo_6_full;
  wire              reorderQueueVec_7_empty;
  assign reorderQueueVec_7_empty = _reorderQueueVec_fifo_7_empty;
  wire              reorderQueueVec_7_full;
  assign reorderQueueVec_7_full = _reorderQueueVec_fifo_7_full;
  wire              readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire              readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire              readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire              readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire              readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire              readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire              readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire              readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire              readMessageQueue_4_empty;
  assign readMessageQueue_4_empty = _readMessageQueue_fifo_4_empty;
  wire              readMessageQueue_4_full;
  assign readMessageQueue_4_full = _readMessageQueue_fifo_4_full;
  wire              readMessageQueue_5_empty;
  assign readMessageQueue_5_empty = _readMessageQueue_fifo_5_empty;
  wire              readMessageQueue_5_full;
  assign readMessageQueue_5_full = _readMessageQueue_fifo_5_full;
  wire              readMessageQueue_6_empty;
  assign readMessageQueue_6_empty = _readMessageQueue_fifo_6_empty;
  wire              readMessageQueue_6_full;
  assign readMessageQueue_6_full = _readMessageQueue_fifo_6_full;
  wire              readMessageQueue_7_empty;
  assign readMessageQueue_7_empty = _readMessageQueue_fifo_7_empty;
  wire              readMessageQueue_7_full;
  assign readMessageQueue_7_full = _readMessageQueue_fifo_7_full;
  wire              readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire              readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire              readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire              readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire              readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  wire              readData_readDataQueue_4_empty;
  assign readData_readDataQueue_4_empty = _readData_readDataQueue_fifo_4_empty;
  wire              readData_readDataQueue_4_full;
  assign readData_readDataQueue_4_full = _readData_readDataQueue_fifo_4_full;
  wire              readData_readDataQueue_5_empty;
  assign readData_readDataQueue_5_empty = _readData_readDataQueue_fifo_5_empty;
  wire              readData_readDataQueue_5_full;
  assign readData_readDataQueue_5_full = _readData_readDataQueue_fifo_5_full;
  wire              readData_readDataQueue_6_empty;
  assign readData_readDataQueue_6_empty = _readData_readDataQueue_fifo_6_empty;
  wire              readData_readDataQueue_6_full;
  assign readData_readDataQueue_6_full = _readData_readDataQueue_fifo_6_full;
  wire              readData_readDataQueue_7_empty;
  assign readData_readDataQueue_7_empty = _readData_readDataQueue_fifo_7_empty;
  wire              readData_readDataQueue_7_full;
  assign readData_readDataQueue_7_full = _readData_readDataQueue_fifo_7_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire              writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire              writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire              writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire              writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire              writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire              writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire              writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire              writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  wire              writeQueue_4_empty;
  assign writeQueue_4_empty = _writeQueue_fifo_4_empty;
  wire              writeQueue_4_full;
  assign writeQueue_4_full = _writeQueue_fifo_4_full;
  wire              writeQueue_5_empty;
  assign writeQueue_5_empty = _writeQueue_fifo_5_empty;
  wire              writeQueue_5_full;
  assign writeQueue_5_full = _writeQueue_fifo_5_full;
  wire              writeQueue_6_empty;
  assign writeQueue_6_empty = _writeQueue_fifo_6_empty;
  wire              writeQueue_6_full;
  assign writeQueue_6_full = _writeQueue_fifo_6_full;
  wire              writeQueue_7_empty;
  assign writeQueue_7_empty = _writeQueue_fifo_7_empty;
  wire              writeQueue_7_full;
  assign writeQueue_7_full = _writeQueue_fifo_7_full;
  BitLevelMaskWrite maskedWrite (
    .clock                             (clock),
    .reset                             (reset),
    .needWAR                           (maskDestinationType),
    .vd                                (instReg_vd),
    .in_0_ready                        (_maskedWrite_in_0_ready),
    .in_0_valid                        (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                    (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                 (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                    (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter            (unitType[2] ? 6'h0 : executeDeqGroupCounter[5:0]),
    .in_0_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                        (_maskedWrite_in_1_ready),
    .in_1_valid                        (executeValid & maskFilter_1),
    .in_1_bits_data                    (executeResult[63:32]),
    .in_1_bits_bitMask                 (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                    (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_1_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                        (_maskedWrite_in_2_ready),
    .in_2_valid                        (executeValid & maskFilter_2),
    .in_2_bits_data                    (executeResult[95:64]),
    .in_2_bits_bitMask                 (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                    (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_2_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                        (_maskedWrite_in_3_ready),
    .in_3_valid                        (executeValid & maskFilter_3),
    .in_3_bits_data                    (executeResult[127:96]),
    .in_3_bits_bitMask                 (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                    (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_3_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .in_4_ready                        (_maskedWrite_in_4_ready),
    .in_4_valid                        (executeValid & maskFilter_4),
    .in_4_bits_data                    (executeResult[159:128]),
    .in_4_bits_bitMask                 (currentMaskGroupForDestination[159:128]),
    .in_4_bits_mask                    (executeWriteByteMask[19:16]),
    .in_4_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_4_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[4] & ffo),
    .in_5_ready                        (_maskedWrite_in_5_ready),
    .in_5_valid                        (executeValid & maskFilter_5),
    .in_5_bits_data                    (executeResult[191:160]),
    .in_5_bits_bitMask                 (currentMaskGroupForDestination[191:160]),
    .in_5_bits_mask                    (executeWriteByteMask[23:20]),
    .in_5_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_5_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[5] & ffo),
    .in_6_ready                        (_maskedWrite_in_6_ready),
    .in_6_valid                        (executeValid & maskFilter_6),
    .in_6_bits_data                    (executeResult[223:192]),
    .in_6_bits_bitMask                 (currentMaskGroupForDestination[223:192]),
    .in_6_bits_mask                    (executeWriteByteMask[27:24]),
    .in_6_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_6_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[6] & ffo),
    .in_7_ready                        (_maskedWrite_in_7_ready),
    .in_7_valid                        (executeValid & maskFilter_7),
    .in_7_bits_data                    (executeResult[255:224]),
    .in_7_bits_bitMask                 (currentMaskGroupForDestination[255:224]),
    .in_7_bits_mask                    (executeWriteByteMask[31:28]),
    .in_7_bits_groupCounter            (executeDeqGroupCounter[5:0]),
    .in_7_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[7] & ffo),
    .out_0_ready                       (writeQueue_0_enq_ready),
    .out_0_valid                       (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther             (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data         (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask         (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                       (writeQueue_1_enq_ready),
    .out_1_valid                       (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther             (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data         (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask         (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                       (writeQueue_2_enq_ready),
    .out_2_valid                       (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther             (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data         (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask         (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                       (writeQueue_3_enq_ready),
    .out_3_valid                       (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther             (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data         (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask         (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter (_maskedWrite_out_3_bits_writeData_groupCounter),
    .out_4_ready                       (writeQueue_4_enq_ready),
    .out_4_valid                       (_maskedWrite_out_4_valid),
    .out_4_bits_ffoByOther             (_maskedWrite_out_4_bits_ffoByOther),
    .out_4_bits_writeData_data         (_maskedWrite_out_4_bits_writeData_data),
    .out_4_bits_writeData_mask         (_maskedWrite_out_4_bits_writeData_mask),
    .out_4_bits_writeData_groupCounter (_maskedWrite_out_4_bits_writeData_groupCounter),
    .out_5_ready                       (writeQueue_5_enq_ready),
    .out_5_valid                       (_maskedWrite_out_5_valid),
    .out_5_bits_ffoByOther             (_maskedWrite_out_5_bits_ffoByOther),
    .out_5_bits_writeData_data         (_maskedWrite_out_5_bits_writeData_data),
    .out_5_bits_writeData_mask         (_maskedWrite_out_5_bits_writeData_mask),
    .out_5_bits_writeData_groupCounter (_maskedWrite_out_5_bits_writeData_groupCounter),
    .out_6_ready                       (writeQueue_6_enq_ready),
    .out_6_valid                       (_maskedWrite_out_6_valid),
    .out_6_bits_ffoByOther             (_maskedWrite_out_6_bits_ffoByOther),
    .out_6_bits_writeData_data         (_maskedWrite_out_6_bits_writeData_data),
    .out_6_bits_writeData_mask         (_maskedWrite_out_6_bits_writeData_mask),
    .out_6_bits_writeData_groupCounter (_maskedWrite_out_6_bits_writeData_groupCounter),
    .out_7_ready                       (writeQueue_7_enq_ready),
    .out_7_valid                       (_maskedWrite_out_7_valid),
    .out_7_bits_ffoByOther             (_maskedWrite_out_7_bits_ffoByOther),
    .out_7_bits_writeData_data         (_maskedWrite_out_7_bits_writeData_data),
    .out_7_bits_writeData_mask         (_maskedWrite_out_7_bits_writeData_mask),
    .out_7_bits_writeData_groupCounter (_maskedWrite_out_7_bits_writeData_groupCounter),
    .readChannel_0_ready               (readChannel_0_ready_0),
    .readChannel_0_valid               (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs             (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset         (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready               (readChannel_1_ready_0),
    .readChannel_1_valid               (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs             (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset         (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready               (readChannel_2_ready_0),
    .readChannel_2_valid               (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs             (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset         (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready               (readChannel_3_ready_0),
    .readChannel_3_valid               (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs             (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset         (_maskedWrite_readChannel_3_bits_offset),
    .readChannel_4_ready               (readChannel_4_ready_0),
    .readChannel_4_valid               (_maskedWrite_readChannel_4_valid),
    .readChannel_4_bits_vs             (_maskedWrite_readChannel_4_bits_vs),
    .readChannel_4_bits_offset         (_maskedWrite_readChannel_4_bits_offset),
    .readChannel_5_ready               (readChannel_5_ready_0),
    .readChannel_5_valid               (_maskedWrite_readChannel_5_valid),
    .readChannel_5_bits_vs             (_maskedWrite_readChannel_5_bits_vs),
    .readChannel_5_bits_offset         (_maskedWrite_readChannel_5_bits_offset),
    .readChannel_6_ready               (readChannel_6_ready_0),
    .readChannel_6_valid               (_maskedWrite_readChannel_6_valid),
    .readChannel_6_bits_vs             (_maskedWrite_readChannel_6_bits_vs),
    .readChannel_6_bits_offset         (_maskedWrite_readChannel_6_bits_offset),
    .readChannel_7_ready               (readChannel_7_ready_0),
    .readChannel_7_valid               (_maskedWrite_readChannel_7_valid),
    .readChannel_7_bits_vs             (_maskedWrite_readChannel_7_bits_vs),
    .readChannel_7_bits_offset         (_maskedWrite_readChannel_7_bits_offset),
    .readResult_0_valid                (readResult_0_valid),
    .readResult_0_bits                 (readResult_0_bits),
    .readResult_1_valid                (readResult_1_valid),
    .readResult_1_bits                 (readResult_1_bits),
    .readResult_2_valid                (readResult_2_valid),
    .readResult_2_bits                 (readResult_2_bits),
    .readResult_3_valid                (readResult_3_valid),
    .readResult_3_bits                 (readResult_3_bits),
    .readResult_4_valid                (readResult_4_valid),
    .readResult_4_bits                 (readResult_4_bits),
    .readResult_5_valid                (readResult_5_valid),
    .readResult_5_bits                 (readResult_5_bits),
    .readResult_6_valid                (readResult_6_valid),
    .readResult_6_bits                 (readResult_6_bits),
    .readResult_7_valid                (readResult_7_valid),
    .readResult_7_bits                 (readResult_7_bits),
    .stageClear                        (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_4_enq_ready & exeRequestQueue_4_enq_valid & ~(_exeRequestQueue_queue_fifo_4_empty & exeRequestQueue_4_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_4_deq_ready & ~_exeRequestQueue_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_4),
    .empty        (_exeRequestQueue_queue_fifo_4_empty),
    .almost_empty (exeRequestQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_4_almostFull),
    .full         (_exeRequestQueue_queue_fifo_4_full),
    .error        (_exeRequestQueue_queue_fifo_4_error),
    .data_out     (_exeRequestQueue_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_5_enq_ready & exeRequestQueue_5_enq_valid & ~(_exeRequestQueue_queue_fifo_5_empty & exeRequestQueue_5_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_5_deq_ready & ~_exeRequestQueue_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_5),
    .empty        (_exeRequestQueue_queue_fifo_5_empty),
    .almost_empty (exeRequestQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_5_almostFull),
    .full         (_exeRequestQueue_queue_fifo_5_full),
    .error        (_exeRequestQueue_queue_fifo_5_error),
    .data_out     (_exeRequestQueue_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_6_enq_ready & exeRequestQueue_6_enq_valid & ~(_exeRequestQueue_queue_fifo_6_empty & exeRequestQueue_6_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_6_deq_ready & ~_exeRequestQueue_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_6),
    .empty        (_exeRequestQueue_queue_fifo_6_empty),
    .almost_empty (exeRequestQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_6_almostFull),
    .full         (_exeRequestQueue_queue_fifo_6_full),
    .error        (_exeRequestQueue_queue_fifo_6_error),
    .data_out     (_exeRequestQueue_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_7_enq_ready & exeRequestQueue_7_enq_valid & ~(_exeRequestQueue_queue_fifo_7_empty & exeRequestQueue_7_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_7_deq_ready & ~_exeRequestQueue_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_7),
    .empty        (_exeRequestQueue_queue_fifo_7_empty),
    .almost_empty (exeRequestQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_7_almostFull),
    .full         (_exeRequestQueue_queue_fifo_7_full),
    .error        (_exeRequestQueue_queue_fifo_7_error),
    .data_out     (_exeRequestQueue_queue_fifo_7_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_accessLane_4         (_slideAddressGen_indexDeq_bits_accessLane_4),
    .indexDeq_bits_accessLane_5         (_slideAddressGen_indexDeq_bits_accessLane_5),
    .indexDeq_bits_accessLane_6         (_slideAddressGen_indexDeq_bits_accessLane_6),
    .indexDeq_bits_accessLane_7         (_slideAddressGen_indexDeq_bits_accessLane_7),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_vsGrowth_4           (_slideAddressGen_indexDeq_bits_vsGrowth_4),
    .indexDeq_bits_vsGrowth_5           (_slideAddressGen_indexDeq_bits_vsGrowth_5),
    .indexDeq_bits_vsGrowth_6           (_slideAddressGen_indexDeq_bits_vsGrowth_6),
    .indexDeq_bits_vsGrowth_7           (_slideAddressGen_indexDeq_bits_vsGrowth_7),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_40[_slideAddressGen_slideGroupOut[6:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready            (_readCrossBar_input_0_ready),
    .input_0_valid            (readCrossBar_input_0_valid),
    .input_0_bits_vs          (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset      (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane    (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset  (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready            (_readCrossBar_input_1_ready),
    .input_1_valid            (readCrossBar_input_1_valid),
    .input_1_bits_vs          (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset      (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane    (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset  (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready            (_readCrossBar_input_2_ready),
    .input_2_valid            (readCrossBar_input_2_valid),
    .input_2_bits_vs          (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset      (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane    (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset  (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready            (_readCrossBar_input_3_ready),
    .input_3_valid            (readCrossBar_input_3_valid),
    .input_3_bits_vs          (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset      (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane    (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset  (selectExecuteReq_3_bits_dataOffset),
    .input_4_ready            (_readCrossBar_input_4_ready),
    .input_4_valid            (readCrossBar_input_4_valid),
    .input_4_bits_vs          (selectExecuteReq_4_bits_vs),
    .input_4_bits_offset      (selectExecuteReq_4_bits_offset),
    .input_4_bits_readLane    (selectExecuteReq_4_bits_readLane),
    .input_4_bits_dataOffset  (selectExecuteReq_4_bits_dataOffset),
    .input_5_ready            (_readCrossBar_input_5_ready),
    .input_5_valid            (readCrossBar_input_5_valid),
    .input_5_bits_vs          (selectExecuteReq_5_bits_vs),
    .input_5_bits_offset      (selectExecuteReq_5_bits_offset),
    .input_5_bits_readLane    (selectExecuteReq_5_bits_readLane),
    .input_5_bits_dataOffset  (selectExecuteReq_5_bits_dataOffset),
    .input_6_ready            (_readCrossBar_input_6_ready),
    .input_6_valid            (readCrossBar_input_6_valid),
    .input_6_bits_vs          (selectExecuteReq_6_bits_vs),
    .input_6_bits_offset      (selectExecuteReq_6_bits_offset),
    .input_6_bits_readLane    (selectExecuteReq_6_bits_readLane),
    .input_6_bits_dataOffset  (selectExecuteReq_6_bits_dataOffset),
    .input_7_ready            (_readCrossBar_input_7_ready),
    .input_7_valid            (readCrossBar_input_7_valid),
    .input_7_bits_vs          (selectExecuteReq_7_bits_vs),
    .input_7_bits_offset      (selectExecuteReq_7_bits_offset),
    .input_7_bits_readLane    (selectExecuteReq_7_bits_readLane),
    .input_7_bits_dataOffset  (selectExecuteReq_7_bits_dataOffset),
    .output_0_ready           (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid           (_readCrossBar_output_0_valid),
    .output_0_bits_vs         (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset     (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready           (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid           (_readCrossBar_output_1_valid),
    .output_1_bits_vs         (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset     (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready           (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid           (_readCrossBar_output_2_valid),
    .output_2_bits_vs         (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset     (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready           (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid           (_readCrossBar_output_3_valid),
    .output_3_bits_vs         (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset     (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset (readMessageQueue_3_enq_bits_dataOffset),
    .output_4_ready           (readChannel_4_ready_0 & readMessageQueue_4_enq_ready),
    .output_4_valid           (_readCrossBar_output_4_valid),
    .output_4_bits_vs         (_readCrossBar_output_4_bits_vs),
    .output_4_bits_offset     (_readCrossBar_output_4_bits_offset),
    .output_4_bits_writeIndex (_readCrossBar_output_4_bits_writeIndex),
    .output_4_bits_dataOffset (readMessageQueue_4_enq_bits_dataOffset),
    .output_5_ready           (readChannel_5_ready_0 & readMessageQueue_5_enq_ready),
    .output_5_valid           (_readCrossBar_output_5_valid),
    .output_5_bits_vs         (_readCrossBar_output_5_bits_vs),
    .output_5_bits_offset     (_readCrossBar_output_5_bits_offset),
    .output_5_bits_writeIndex (_readCrossBar_output_5_bits_writeIndex),
    .output_5_bits_dataOffset (readMessageQueue_5_enq_bits_dataOffset),
    .output_6_ready           (readChannel_6_ready_0 & readMessageQueue_6_enq_ready),
    .output_6_valid           (_readCrossBar_output_6_valid),
    .output_6_bits_vs         (_readCrossBar_output_6_bits_vs),
    .output_6_bits_offset     (_readCrossBar_output_6_bits_offset),
    .output_6_bits_writeIndex (_readCrossBar_output_6_bits_writeIndex),
    .output_6_bits_dataOffset (readMessageQueue_6_enq_bits_dataOffset),
    .output_7_ready           (readChannel_7_ready_0 & readMessageQueue_7_enq_ready),
    .output_7_valid           (_readCrossBar_output_7_valid),
    .output_7_bits_vs         (_readCrossBar_output_7_bits_vs),
    .output_7_bits_offset     (_readCrossBar_output_7_bits_offset),
    .output_7_bits_writeIndex (_readCrossBar_output_7_bits_writeIndex),
    .output_7_bits_dataOffset (readMessageQueue_7_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(33)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(303)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_4_enq_ready & reorderQueueVec_4_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_4_deq_ready & ~_reorderQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_4),
    .empty        (_reorderQueueVec_fifo_4_empty),
    .almost_empty (reorderQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_4_almostFull),
    .full         (_reorderQueueVec_fifo_4_full),
    .error        (_reorderQueueVec_fifo_4_error),
    .data_out     (_reorderQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_5_enq_ready & reorderQueueVec_5_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_5_deq_ready & ~_reorderQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_5),
    .empty        (_reorderQueueVec_fifo_5_empty),
    .almost_empty (reorderQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_5_almostFull),
    .full         (_reorderQueueVec_fifo_5_full),
    .error        (_reorderQueueVec_fifo_5_error),
    .data_out     (_reorderQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_6_enq_ready & reorderQueueVec_6_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_6_deq_ready & ~_reorderQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_6),
    .empty        (_reorderQueueVec_fifo_6_empty),
    .almost_empty (reorderQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_6_almostFull),
    .full         (_reorderQueueVec_fifo_6_full),
    .error        (_reorderQueueVec_fifo_6_error),
    .data_out     (_reorderQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(16),
    .err_mode(2),
    .rst_mode(3),
    .width(40)
  ) reorderQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_7_enq_ready & reorderQueueVec_7_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_7_deq_ready & ~_reorderQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_7),
    .empty        (_reorderQueueVec_fifo_7_empty),
    .almost_empty (reorderQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_7_almostFull),
    .full         (_reorderQueueVec_fifo_7_full),
    .error        (_reorderQueueVec_fifo_7_error),
    .data_out     (_reorderQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_4_enq_ready & readMessageQueue_4_enq_valid)),
    .pop_req_n    (~(readMessageQueue_4_deq_ready & ~_readMessageQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_4),
    .empty        (_readMessageQueue_fifo_4_empty),
    .almost_empty (readMessageQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_4_almostFull),
    .full         (_readMessageQueue_fifo_4_full),
    .error        (_readMessageQueue_fifo_4_error),
    .data_out     (_readMessageQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_5_enq_ready & readMessageQueue_5_enq_valid)),
    .pop_req_n    (~(readMessageQueue_5_deq_ready & ~_readMessageQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_5),
    .empty        (_readMessageQueue_fifo_5_empty),
    .almost_empty (readMessageQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_5_almostFull),
    .full         (_readMessageQueue_fifo_5_full),
    .error        (_readMessageQueue_fifo_5_error),
    .data_out     (_readMessageQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_6_enq_ready & readMessageQueue_6_enq_valid)),
    .pop_req_n    (~(readMessageQueue_6_deq_ready & ~_readMessageQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_6),
    .empty        (_readMessageQueue_fifo_6_empty),
    .almost_empty (readMessageQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_6_almostFull),
    .full         (_readMessageQueue_fifo_6_full),
    .error        (_readMessageQueue_fifo_6_error),
    .data_out     (_readMessageQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) readMessageQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_7_enq_ready & readMessageQueue_7_enq_valid)),
    .pop_req_n    (~(readMessageQueue_7_deq_ready & ~_readMessageQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_7),
    .empty        (_readMessageQueue_fifo_7_empty),
    .almost_empty (readMessageQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_7_almostFull),
    .full         (_readMessageQueue_fifo_7_full),
    .error        (_readMessageQueue_fifo_7_error),
    .data_out     (_readMessageQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_4_enq_ready & readData_readDataQueue_4_enq_valid & ~(_readData_readDataQueue_fifo_4_empty & readData_readDataQueue_4_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_4_deq_ready & ~_readData_readDataQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_4_enq_bits),
    .empty        (_readData_readDataQueue_fifo_4_empty),
    .almost_empty (readData_readDataQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_4_almostFull),
    .full         (_readData_readDataQueue_fifo_4_full),
    .error        (_readData_readDataQueue_fifo_4_error),
    .data_out     (_readData_readDataQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_5_enq_ready & readData_readDataQueue_5_enq_valid & ~(_readData_readDataQueue_fifo_5_empty & readData_readDataQueue_5_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_5_deq_ready & ~_readData_readDataQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_5_enq_bits),
    .empty        (_readData_readDataQueue_fifo_5_empty),
    .almost_empty (readData_readDataQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_5_almostFull),
    .full         (_readData_readDataQueue_fifo_5_full),
    .error        (_readData_readDataQueue_fifo_5_error),
    .data_out     (_readData_readDataQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_6_enq_ready & readData_readDataQueue_6_enq_valid & ~(_readData_readDataQueue_fifo_6_empty & readData_readDataQueue_6_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_6_deq_ready & ~_readData_readDataQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_6_enq_bits),
    .empty        (_readData_readDataQueue_fifo_6_empty),
    .almost_empty (readData_readDataQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_6_almostFull),
    .full         (_readData_readDataQueue_fifo_6_full),
    .error        (_readData_readDataQueue_fifo_6_error),
    .data_out     (_readData_readDataQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_7_enq_ready & readData_readDataQueue_7_enq_valid & ~(_readData_readDataQueue_fifo_7_empty & readData_readDataQueue_7_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_7_deq_ready & ~_readData_readDataQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_7_enq_bits),
    .empty        (_readData_readDataQueue_fifo_7_empty),
    .almost_empty (readData_readDataQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_7_almostFull),
    .full         (_readData_readDataQueue_fifo_7_full),
    .error        (_readData_readDataQueue_fifo_7_error),
    .data_out     (_readData_readDataQueue_fifo_7_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           (executeElementMask),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock                 (clock),
    .reset                 (reset),
    .in_ready              (_reduceUnit_in_ready),
    .in_valid              (reduceUnit_in_valid),
    .in_bits_maskType      (instReg_maskType),
    .in_bits_eew           (instReg_sew),
    .in_bits_uop           (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1       (readVS1Reg_data),
    .in_bits_source2       (source2),
    .in_bits_sourceValid   ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup     (lastGroup),
    .in_bits_vxrm          (instReg_vxrm),
    .in_bits_aluUop        (instReg_decodeResult_uop),
    .in_bits_sign          (~instReg_decodeResult_unsigned1),
    .in_bits_fpSourceValid ({view__in_bits_fpSourceValid_hi, view__in_bits_fpSourceValid_lo}),
    .out_valid             (_reduceUnit_out_valid),
    .out_bits_data         (_reduceUnit_out_bits_data),
    .out_bits_mask         (_reduceUnit_out_bits_mask),
    .firstGroup            (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction        (instReq_valid),
    .validInst             (|instReg_vl),
    .pop                   (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[5:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_4_enq_ready & writeQueue_4_enq_valid)),
    .pop_req_n    (~(writeQueue_4_deq_ready & ~_writeQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_4),
    .empty        (_writeQueue_fifo_4_empty),
    .almost_empty (writeQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_4_almostFull),
    .full         (_writeQueue_fifo_4_full),
    .error        (_writeQueue_fifo_4_error),
    .data_out     (_writeQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_5_enq_ready & writeQueue_5_enq_valid)),
    .pop_req_n    (~(writeQueue_5_deq_ready & ~_writeQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_5),
    .empty        (_writeQueue_fifo_5_empty),
    .almost_empty (writeQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_5_almostFull),
    .full         (_writeQueue_fifo_5_full),
    .error        (_writeQueue_fifo_5_error),
    .data_out     (_writeQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_6_enq_ready & writeQueue_6_enq_valid)),
    .pop_req_n    (~(writeQueue_6_deq_ready & ~_writeQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_6),
    .empty        (_writeQueue_fifo_6_empty),
    .almost_empty (writeQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_6_almostFull),
    .full         (_writeQueue_fifo_6_full),
    .error        (_writeQueue_fifo_6_error),
    .data_out     (_writeQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) writeQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_7_enq_ready & writeQueue_7_enq_valid)),
    .pop_req_n    (~(writeQueue_7_deq_ready & ~_writeQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_7),
    .empty        (_writeQueue_fifo_7_empty),
    .almost_empty (writeQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_7_almostFull),
    .full         (_writeQueue_fifo_7_full),
    .error        (_writeQueue_fifo_7_error),
    .data_out     (_writeQueue_fifo_7_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign exeResp_4_valid = exeResp_4_valid_0;
  assign exeResp_4_bits_vd = exeResp_4_bits_vd_0;
  assign exeResp_4_bits_offset = exeResp_4_bits_offset_0;
  assign exeResp_4_bits_mask = exeResp_4_bits_mask_0;
  assign exeResp_4_bits_data = exeResp_4_bits_data_0;
  assign exeResp_4_bits_instructionIndex = exeResp_4_bits_instructionIndex_0;
  assign exeResp_5_valid = exeResp_5_valid_0;
  assign exeResp_5_bits_vd = exeResp_5_bits_vd_0;
  assign exeResp_5_bits_offset = exeResp_5_bits_offset_0;
  assign exeResp_5_bits_mask = exeResp_5_bits_mask_0;
  assign exeResp_5_bits_data = exeResp_5_bits_data_0;
  assign exeResp_5_bits_instructionIndex = exeResp_5_bits_instructionIndex_0;
  assign exeResp_6_valid = exeResp_6_valid_0;
  assign exeResp_6_bits_vd = exeResp_6_bits_vd_0;
  assign exeResp_6_bits_offset = exeResp_6_bits_offset_0;
  assign exeResp_6_bits_mask = exeResp_6_bits_mask_0;
  assign exeResp_6_bits_data = exeResp_6_bits_data_0;
  assign exeResp_6_bits_instructionIndex = exeResp_6_bits_instructionIndex_0;
  assign exeResp_7_valid = exeResp_7_valid_0;
  assign exeResp_7_bits_vd = exeResp_7_bits_vd_0;
  assign exeResp_7_bits_offset = exeResp_7_bits_offset_0;
  assign exeResp_7_bits_mask = exeResp_7_bits_mask_0;
  assign exeResp_7_bits_data = exeResp_7_bits_data_0;
  assign exeResp_7_bits_instructionIndex = exeResp_7_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign tokenIO_4_maskRequestRelease = tokenIO_4_maskRequestRelease_0;
  assign tokenIO_5_maskRequestRelease = tokenIO_5_maskRequestRelease_0;
  assign tokenIO_6_maskRequestRelease = tokenIO_6_maskRequestRelease_0;
  assign tokenIO_7_maskRequestRelease = tokenIO_7_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign readChannel_4_valid = readChannel_4_valid_0;
  assign readChannel_4_bits_vs = readChannel_4_bits_vs_0;
  assign readChannel_4_bits_offset = readChannel_4_bits_offset_0;
  assign readChannel_4_bits_instructionIndex = readChannel_4_bits_instructionIndex_0;
  assign readChannel_5_valid = readChannel_5_valid_0;
  assign readChannel_5_bits_vs = readChannel_5_bits_vs_0;
  assign readChannel_5_bits_offset = readChannel_5_bits_offset_0;
  assign readChannel_5_bits_instructionIndex = readChannel_5_bits_instructionIndex_0;
  assign readChannel_6_valid = readChannel_6_valid_0;
  assign readChannel_6_bits_vs = readChannel_6_bits_vs_0;
  assign readChannel_6_bits_offset = readChannel_6_bits_offset_0;
  assign readChannel_6_bits_instructionIndex = readChannel_6_bits_instructionIndex_0;
  assign readChannel_7_valid = readChannel_7_valid_0;
  assign readChannel_7_bits_vs = readChannel_7_bits_vs_0;
  assign readChannel_7_bits_offset = readChannel_7_bits_offset_0;
  assign readChannel_7_bits_instructionIndex = readChannel_7_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = _GEN_15[laneMaskSelect_0[1:0]];
  assign laneMaskInput_1 = _GEN_16[laneMaskSelect_1[1:0]];
  assign laneMaskInput_2 = _GEN_17[laneMaskSelect_2[1:0]];
  assign laneMaskInput_3 = _GEN_18[laneMaskSelect_3[1:0]];
  assign laneMaskInput_4 = _GEN_19[laneMaskSelect_4[1:0]];
  assign laneMaskInput_5 = _GEN_20[laneMaskSelect_5[1:0]];
  assign laneMaskInput_6 = _GEN_21[laneMaskSelect_6[1:0]];
  assign laneMaskInput_7 = _GEN_22[laneMaskSelect_7[1:0]];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

