module MaskUnitReadCrossBar(
  output       input_0_ready,
  input        input_0_valid,
  input  [4:0] input_0_bits_vs,
  input  [1:0] input_0_bits_offset,
  input  [2:0] input_0_bits_readLane,
  input  [1:0] input_0_bits_dataOffset,
  output       input_1_ready,
  input        input_1_valid,
  input  [4:0] input_1_bits_vs,
  input  [1:0] input_1_bits_offset,
  input  [2:0] input_1_bits_readLane,
  input  [1:0] input_1_bits_dataOffset,
  output       input_2_ready,
  input        input_2_valid,
  input  [4:0] input_2_bits_vs,
  input  [1:0] input_2_bits_offset,
  input  [2:0] input_2_bits_readLane,
  input  [1:0] input_2_bits_dataOffset,
  output       input_3_ready,
  input        input_3_valid,
  input  [4:0] input_3_bits_vs,
  input  [1:0] input_3_bits_offset,
  input  [2:0] input_3_bits_readLane,
  input  [1:0] input_3_bits_dataOffset,
  output       input_4_ready,
  input        input_4_valid,
  input  [4:0] input_4_bits_vs,
  input  [1:0] input_4_bits_offset,
  input  [2:0] input_4_bits_readLane,
  input  [1:0] input_4_bits_dataOffset,
  output       input_5_ready,
  input        input_5_valid,
  input  [4:0] input_5_bits_vs,
  input  [1:0] input_5_bits_offset,
  input  [2:0] input_5_bits_readLane,
  input  [1:0] input_5_bits_dataOffset,
  output       input_6_ready,
  input        input_6_valid,
  input  [4:0] input_6_bits_vs,
  input  [1:0] input_6_bits_offset,
  input  [2:0] input_6_bits_readLane,
  input  [1:0] input_6_bits_dataOffset,
  output       input_7_ready,
  input        input_7_valid,
  input  [4:0] input_7_bits_vs,
  input  [1:0] input_7_bits_offset,
  input  [2:0] input_7_bits_readLane,
  input  [1:0] input_7_bits_dataOffset,
  input        output_0_ready,
  output       output_0_valid,
  output [4:0] output_0_bits_vs,
  output [1:0] output_0_bits_offset,
  output [2:0] output_0_bits_writeIndex,
  output [1:0] output_0_bits_dataOffset,
  input        output_1_ready,
  output       output_1_valid,
  output [4:0] output_1_bits_vs,
  output [1:0] output_1_bits_offset,
  output [2:0] output_1_bits_writeIndex,
  output [1:0] output_1_bits_dataOffset,
  input        output_2_ready,
  output       output_2_valid,
  output [4:0] output_2_bits_vs,
  output [1:0] output_2_bits_offset,
  output [2:0] output_2_bits_writeIndex,
  output [1:0] output_2_bits_dataOffset,
  input        output_3_ready,
  output       output_3_valid,
  output [4:0] output_3_bits_vs,
  output [1:0] output_3_bits_offset,
  output [2:0] output_3_bits_writeIndex,
  output [1:0] output_3_bits_dataOffset,
  input        output_4_ready,
  output       output_4_valid,
  output [4:0] output_4_bits_vs,
  output [1:0] output_4_bits_offset,
  output [2:0] output_4_bits_writeIndex,
  output [1:0] output_4_bits_dataOffset,
  input        output_5_ready,
  output       output_5_valid,
  output [4:0] output_5_bits_vs,
  output [1:0] output_5_bits_offset,
  output [2:0] output_5_bits_writeIndex,
  output [1:0] output_5_bits_dataOffset,
  input        output_6_ready,
  output       output_6_valid,
  output [4:0] output_6_bits_vs,
  output [1:0] output_6_bits_offset,
  output [2:0] output_6_bits_writeIndex,
  output [1:0] output_6_bits_dataOffset,
  input        output_7_ready,
  output       output_7_valid,
  output [4:0] output_7_bits_vs,
  output [1:0] output_7_bits_offset,
  output [2:0] output_7_bits_writeIndex,
  output [1:0] output_7_bits_dataOffset
);

  wire       input_0_valid_0 = input_0_valid;
  wire [4:0] input_0_bits_vs_0 = input_0_bits_vs;
  wire [1:0] input_0_bits_offset_0 = input_0_bits_offset;
  wire [2:0] input_0_bits_readLane_0 = input_0_bits_readLane;
  wire [1:0] input_0_bits_dataOffset_0 = input_0_bits_dataOffset;
  wire       input_1_valid_0 = input_1_valid;
  wire [4:0] input_1_bits_vs_0 = input_1_bits_vs;
  wire [1:0] input_1_bits_offset_0 = input_1_bits_offset;
  wire [2:0] input_1_bits_readLane_0 = input_1_bits_readLane;
  wire [1:0] input_1_bits_dataOffset_0 = input_1_bits_dataOffset;
  wire       input_2_valid_0 = input_2_valid;
  wire [4:0] input_2_bits_vs_0 = input_2_bits_vs;
  wire [1:0] input_2_bits_offset_0 = input_2_bits_offset;
  wire [2:0] input_2_bits_readLane_0 = input_2_bits_readLane;
  wire [1:0] input_2_bits_dataOffset_0 = input_2_bits_dataOffset;
  wire       input_3_valid_0 = input_3_valid;
  wire [4:0] input_3_bits_vs_0 = input_3_bits_vs;
  wire [1:0] input_3_bits_offset_0 = input_3_bits_offset;
  wire [2:0] input_3_bits_readLane_0 = input_3_bits_readLane;
  wire [1:0] input_3_bits_dataOffset_0 = input_3_bits_dataOffset;
  wire       input_4_valid_0 = input_4_valid;
  wire [4:0] input_4_bits_vs_0 = input_4_bits_vs;
  wire [1:0] input_4_bits_offset_0 = input_4_bits_offset;
  wire [2:0] input_4_bits_readLane_0 = input_4_bits_readLane;
  wire [1:0] input_4_bits_dataOffset_0 = input_4_bits_dataOffset;
  wire       input_5_valid_0 = input_5_valid;
  wire [4:0] input_5_bits_vs_0 = input_5_bits_vs;
  wire [1:0] input_5_bits_offset_0 = input_5_bits_offset;
  wire [2:0] input_5_bits_readLane_0 = input_5_bits_readLane;
  wire [1:0] input_5_bits_dataOffset_0 = input_5_bits_dataOffset;
  wire       input_6_valid_0 = input_6_valid;
  wire [4:0] input_6_bits_vs_0 = input_6_bits_vs;
  wire [1:0] input_6_bits_offset_0 = input_6_bits_offset;
  wire [2:0] input_6_bits_readLane_0 = input_6_bits_readLane;
  wire [1:0] input_6_bits_dataOffset_0 = input_6_bits_dataOffset;
  wire       input_7_valid_0 = input_7_valid;
  wire [4:0] input_7_bits_vs_0 = input_7_bits_vs;
  wire [1:0] input_7_bits_offset_0 = input_7_bits_offset;
  wire [2:0] input_7_bits_readLane_0 = input_7_bits_readLane;
  wire [1:0] input_7_bits_dataOffset_0 = input_7_bits_dataOffset;
  wire       output_0_ready_0 = output_0_ready;
  wire       output_1_ready_0 = output_1_ready;
  wire       output_2_ready_0 = output_2_ready;
  wire       output_3_ready_0 = output_3_ready;
  wire       output_4_ready_0 = output_4_ready;
  wire       output_5_ready_0 = output_5_ready;
  wire       output_6_ready_0 = output_6_ready;
  wire       output_7_ready_0 = output_7_ready;
  wire [2:0] input_7_bits_requestIndex = 3'h7;
  wire [2:0] input_6_bits_requestIndex = 3'h6;
  wire [2:0] input_5_bits_requestIndex = 3'h5;
  wire [2:0] input_4_bits_requestIndex = 3'h4;
  wire [2:0] input_3_bits_requestIndex = 3'h3;
  wire [2:0] input_2_bits_requestIndex = 3'h2;
  wire [2:0] input_1_bits_requestIndex = 3'h1;
  wire [2:0] input_0_bits_requestIndex = 3'h0;
  wire [4:0] selectReq_bits_vs;
  wire [1:0] selectReq_bits_offset;
  wire [2:0] selectReq_bits_requestIndex;
  wire [1:0] selectReq_bits_dataOffset;
  wire [4:0] selectReq_1_bits_vs;
  wire [1:0] selectReq_1_bits_offset;
  wire [2:0] selectReq_1_bits_requestIndex;
  wire [1:0] selectReq_1_bits_dataOffset;
  wire [4:0] selectReq_2_bits_vs;
  wire [1:0] selectReq_2_bits_offset;
  wire [2:0] selectReq_2_bits_requestIndex;
  wire [1:0] selectReq_2_bits_dataOffset;
  wire [4:0] selectReq_3_bits_vs;
  wire [1:0] selectReq_3_bits_offset;
  wire [2:0] selectReq_3_bits_requestIndex;
  wire [1:0] selectReq_3_bits_dataOffset;
  wire [4:0] selectReq_4_bits_vs;
  wire [1:0] selectReq_4_bits_offset;
  wire [2:0] selectReq_4_bits_requestIndex;
  wire [1:0] selectReq_4_bits_dataOffset;
  wire [4:0] selectReq_5_bits_vs;
  wire [1:0] selectReq_5_bits_offset;
  wire [2:0] selectReq_5_bits_requestIndex;
  wire [1:0] selectReq_5_bits_dataOffset;
  wire [4:0] selectReq_6_bits_vs;
  wire [1:0] selectReq_6_bits_offset;
  wire [2:0] selectReq_6_bits_requestIndex;
  wire [1:0] selectReq_6_bits_dataOffset;
  wire [4:0] selectReq_7_bits_vs;
  wire [1:0] selectReq_7_bits_offset;
  wire [2:0] selectReq_7_bits_requestIndex;
  wire [1:0] selectReq_7_bits_dataOffset;
  wire [7:0] requestReadLane = 8'h1 << input_0_bits_readLane_0;
  wire       free = |requestReadLane;
  wire       outReady =
    requestReadLane[0] & output_0_ready_0 | requestReadLane[1] & output_1_ready_0 | requestReadLane[2] & output_2_ready_0 | requestReadLane[3] & output_3_ready_0 | requestReadLane[4] & output_4_ready_0 | requestReadLane[5]
    & output_5_ready_0 | requestReadLane[6] & output_6_ready_0 | requestReadLane[7] & output_7_ready_0;
  wire       input_0_ready_0 = free & outReady;
  wire [7:0] inputSelect1H_0 = input_0_valid_0 & free ? requestReadLane : 8'h0;
  wire [7:0] requestReadLane_1 = 8'h1 << input_1_bits_readLane_0;
  wire       free_1 = |(requestReadLane_1 & ~inputSelect1H_0);
  wire       outReady_1 =
    requestReadLane_1[0] & output_0_ready_0 | requestReadLane_1[1] & output_1_ready_0 | requestReadLane_1[2] & output_2_ready_0 | requestReadLane_1[3] & output_3_ready_0 | requestReadLane_1[4] & output_4_ready_0 | requestReadLane_1[5]
    & output_5_ready_0 | requestReadLane_1[6] & output_6_ready_0 | requestReadLane_1[7] & output_7_ready_0;
  wire       input_1_ready_0 = free_1 & outReady_1;
  wire [7:0] inputSelect1H_1 = input_1_valid_0 & free_1 ? requestReadLane_1 : 8'h0;
  wire [7:0] _GEN = inputSelect1H_0 | inputSelect1H_1;
  wire [7:0] requestReadLane_2 = 8'h1 << input_2_bits_readLane_0;
  wire       free_2 = |(requestReadLane_2 & ~_GEN);
  wire       outReady_2 =
    requestReadLane_2[0] & output_0_ready_0 | requestReadLane_2[1] & output_1_ready_0 | requestReadLane_2[2] & output_2_ready_0 | requestReadLane_2[3] & output_3_ready_0 | requestReadLane_2[4] & output_4_ready_0 | requestReadLane_2[5]
    & output_5_ready_0 | requestReadLane_2[6] & output_6_ready_0 | requestReadLane_2[7] & output_7_ready_0;
  wire       input_2_ready_0 = free_2 & outReady_2;
  wire [7:0] inputSelect1H_2 = input_2_valid_0 & free_2 ? requestReadLane_2 : 8'h0;
  wire [7:0] _GEN_0 = _GEN | inputSelect1H_2;
  wire [7:0] requestReadLane_3 = 8'h1 << input_3_bits_readLane_0;
  wire       free_3 = |(requestReadLane_3 & ~_GEN_0);
  wire       outReady_3 =
    requestReadLane_3[0] & output_0_ready_0 | requestReadLane_3[1] & output_1_ready_0 | requestReadLane_3[2] & output_2_ready_0 | requestReadLane_3[3] & output_3_ready_0 | requestReadLane_3[4] & output_4_ready_0 | requestReadLane_3[5]
    & output_5_ready_0 | requestReadLane_3[6] & output_6_ready_0 | requestReadLane_3[7] & output_7_ready_0;
  wire       input_3_ready_0 = free_3 & outReady_3;
  wire [7:0] inputSelect1H_3 = input_3_valid_0 & free_3 ? requestReadLane_3 : 8'h0;
  wire [7:0] _GEN_1 = _GEN_0 | inputSelect1H_3;
  wire [7:0] requestReadLane_4 = 8'h1 << input_4_bits_readLane_0;
  wire       free_4 = |(requestReadLane_4 & ~_GEN_1);
  wire       outReady_4 =
    requestReadLane_4[0] & output_0_ready_0 | requestReadLane_4[1] & output_1_ready_0 | requestReadLane_4[2] & output_2_ready_0 | requestReadLane_4[3] & output_3_ready_0 | requestReadLane_4[4] & output_4_ready_0 | requestReadLane_4[5]
    & output_5_ready_0 | requestReadLane_4[6] & output_6_ready_0 | requestReadLane_4[7] & output_7_ready_0;
  wire       input_4_ready_0 = free_4 & outReady_4;
  wire [7:0] inputSelect1H_4 = input_4_valid_0 & free_4 ? requestReadLane_4 : 8'h0;
  wire [7:0] _GEN_2 = _GEN_1 | inputSelect1H_4;
  wire [7:0] requestReadLane_5 = 8'h1 << input_5_bits_readLane_0;
  wire       free_5 = |(requestReadLane_5 & ~_GEN_2);
  wire       outReady_5 =
    requestReadLane_5[0] & output_0_ready_0 | requestReadLane_5[1] & output_1_ready_0 | requestReadLane_5[2] & output_2_ready_0 | requestReadLane_5[3] & output_3_ready_0 | requestReadLane_5[4] & output_4_ready_0 | requestReadLane_5[5]
    & output_5_ready_0 | requestReadLane_5[6] & output_6_ready_0 | requestReadLane_5[7] & output_7_ready_0;
  wire       input_5_ready_0 = free_5 & outReady_5;
  wire [7:0] inputSelect1H_5 = input_5_valid_0 & free_5 ? requestReadLane_5 : 8'h0;
  wire [7:0] _GEN_3 = _GEN_2 | inputSelect1H_5;
  wire [7:0] requestReadLane_6 = 8'h1 << input_6_bits_readLane_0;
  wire       free_6 = |(requestReadLane_6 & ~_GEN_3);
  wire       outReady_6 =
    requestReadLane_6[0] & output_0_ready_0 | requestReadLane_6[1] & output_1_ready_0 | requestReadLane_6[2] & output_2_ready_0 | requestReadLane_6[3] & output_3_ready_0 | requestReadLane_6[4] & output_4_ready_0 | requestReadLane_6[5]
    & output_5_ready_0 | requestReadLane_6[6] & output_6_ready_0 | requestReadLane_6[7] & output_7_ready_0;
  wire       input_6_ready_0 = free_6 & outReady_6;
  wire [7:0] inputSelect1H_6 = input_6_valid_0 & free_6 ? requestReadLane_6 : 8'h0;
  wire [7:0] requestReadLane_7 = 8'h1 << input_7_bits_readLane_0;
  wire       free_7 = |(requestReadLane_7 & ~(_GEN_3 | inputSelect1H_6));
  wire       outReady_7 =
    requestReadLane_7[0] & output_0_ready_0 | requestReadLane_7[1] & output_1_ready_0 | requestReadLane_7[2] & output_2_ready_0 | requestReadLane_7[3] & output_3_ready_0 | requestReadLane_7[4] & output_4_ready_0 | requestReadLane_7[5]
    & output_5_ready_0 | requestReadLane_7[6] & output_6_ready_0 | requestReadLane_7[7] & output_7_ready_0;
  wire       input_7_ready_0 = free_7 & outReady_7;
  wire [7:0] inputSelect1H_7 = input_7_valid_0 & free_7 ? requestReadLane_7 : 8'h0;
  wire [1:0] tryToRead_lo_lo = {inputSelect1H_1[0], inputSelect1H_0[0]};
  wire [1:0] tryToRead_lo_hi = {inputSelect1H_3[0], inputSelect1H_2[0]};
  wire [3:0] tryToRead_lo = {tryToRead_lo_hi, tryToRead_lo_lo};
  wire [1:0] tryToRead_hi_lo = {inputSelect1H_5[0], inputSelect1H_4[0]};
  wire [1:0] tryToRead_hi_hi = {inputSelect1H_7[0], inputSelect1H_6[0]};
  wire [3:0] tryToRead_hi = {tryToRead_hi_hi, tryToRead_hi_lo};
  wire [7:0] tryToRead = {tryToRead_hi, tryToRead_lo};
  wire       output_0_valid_0 = |tryToRead;
  wire [4:0] output_0_bits_vs_0 = selectReq_bits_vs;
  wire [1:0] output_0_bits_offset_0 = selectReq_bits_offset;
  wire [2:0] output_0_bits_writeIndex_0 = selectReq_bits_requestIndex;
  wire [1:0] output_0_bits_dataOffset_0 = selectReq_bits_dataOffset;
  assign selectReq_bits_dataOffset =
    (tryToRead[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_bits_requestIndex = {2'h0, tryToRead[1]} | {1'h0, tryToRead[2], 1'h0} | (tryToRead[3] ? 3'h3 : 3'h0) | {tryToRead[4], 2'h0} | (tryToRead[5] ? 3'h5 : 3'h0) | (tryToRead[6] ? 3'h6 : 3'h0) | {3{tryToRead[7]}};
  wire [2:0] selectReq_bits_readLane =
    (tryToRead[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_bits_offset =
    (tryToRead[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_bits_vs =
    (tryToRead[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_valid =
    tryToRead[0] & input_0_valid_0 | tryToRead[1] & input_1_valid_0 | tryToRead[2] & input_2_valid_0 | tryToRead[3] & input_3_valid_0 | tryToRead[4] & input_4_valid_0 | tryToRead[5] & input_5_valid_0 | tryToRead[6] & input_6_valid_0
    | tryToRead[7] & input_7_valid_0;
  wire       selectReq_ready =
    tryToRead[0] & input_0_ready_0 | tryToRead[1] & input_1_ready_0 | tryToRead[2] & input_2_ready_0 | tryToRead[3] & input_3_ready_0 | tryToRead[4] & input_4_ready_0 | tryToRead[5] & input_5_ready_0 | tryToRead[6] & input_6_ready_0
    | tryToRead[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_1 = {inputSelect1H_1[1], inputSelect1H_0[1]};
  wire [1:0] tryToRead_lo_hi_1 = {inputSelect1H_3[1], inputSelect1H_2[1]};
  wire [3:0] tryToRead_lo_1 = {tryToRead_lo_hi_1, tryToRead_lo_lo_1};
  wire [1:0] tryToRead_hi_lo_1 = {inputSelect1H_5[1], inputSelect1H_4[1]};
  wire [1:0] tryToRead_hi_hi_1 = {inputSelect1H_7[1], inputSelect1H_6[1]};
  wire [3:0] tryToRead_hi_1 = {tryToRead_hi_hi_1, tryToRead_hi_lo_1};
  wire [7:0] tryToRead_1 = {tryToRead_hi_1, tryToRead_lo_1};
  wire       output_1_valid_0 = |tryToRead_1;
  wire [4:0] output_1_bits_vs_0 = selectReq_1_bits_vs;
  wire [1:0] output_1_bits_offset_0 = selectReq_1_bits_offset;
  wire [2:0] output_1_bits_writeIndex_0 = selectReq_1_bits_requestIndex;
  wire [1:0] output_1_bits_dataOffset_0 = selectReq_1_bits_dataOffset;
  assign selectReq_1_bits_dataOffset =
    (tryToRead_1[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_1[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_1[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_1[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_1[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_1[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_1[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_1_bits_requestIndex =
    {2'h0, tryToRead_1[1]} | {1'h0, tryToRead_1[2], 1'h0} | (tryToRead_1[3] ? 3'h3 : 3'h0) | {tryToRead_1[4], 2'h0} | (tryToRead_1[5] ? 3'h5 : 3'h0) | (tryToRead_1[6] ? 3'h6 : 3'h0) | {3{tryToRead_1[7]}};
  wire [2:0] selectReq_1_bits_readLane =
    (tryToRead_1[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_1[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_1[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_1[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_1[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_1[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_1[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_1[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_1_bits_offset =
    (tryToRead_1[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_1[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_1[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_1[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_1[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_1[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_1[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_1[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_1_bits_vs =
    (tryToRead_1[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_1[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_1[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_1[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_1[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_1[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_1[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_1[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_1_valid =
    tryToRead_1[0] & input_0_valid_0 | tryToRead_1[1] & input_1_valid_0 | tryToRead_1[2] & input_2_valid_0 | tryToRead_1[3] & input_3_valid_0 | tryToRead_1[4] & input_4_valid_0 | tryToRead_1[5] & input_5_valid_0 | tryToRead_1[6]
    & input_6_valid_0 | tryToRead_1[7] & input_7_valid_0;
  wire       selectReq_1_ready =
    tryToRead_1[0] & input_0_ready_0 | tryToRead_1[1] & input_1_ready_0 | tryToRead_1[2] & input_2_ready_0 | tryToRead_1[3] & input_3_ready_0 | tryToRead_1[4] & input_4_ready_0 | tryToRead_1[5] & input_5_ready_0 | tryToRead_1[6]
    & input_6_ready_0 | tryToRead_1[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_2 = {inputSelect1H_1[2], inputSelect1H_0[2]};
  wire [1:0] tryToRead_lo_hi_2 = {inputSelect1H_3[2], inputSelect1H_2[2]};
  wire [3:0] tryToRead_lo_2 = {tryToRead_lo_hi_2, tryToRead_lo_lo_2};
  wire [1:0] tryToRead_hi_lo_2 = {inputSelect1H_5[2], inputSelect1H_4[2]};
  wire [1:0] tryToRead_hi_hi_2 = {inputSelect1H_7[2], inputSelect1H_6[2]};
  wire [3:0] tryToRead_hi_2 = {tryToRead_hi_hi_2, tryToRead_hi_lo_2};
  wire [7:0] tryToRead_2 = {tryToRead_hi_2, tryToRead_lo_2};
  wire       output_2_valid_0 = |tryToRead_2;
  wire [4:0] output_2_bits_vs_0 = selectReq_2_bits_vs;
  wire [1:0] output_2_bits_offset_0 = selectReq_2_bits_offset;
  wire [2:0] output_2_bits_writeIndex_0 = selectReq_2_bits_requestIndex;
  wire [1:0] output_2_bits_dataOffset_0 = selectReq_2_bits_dataOffset;
  assign selectReq_2_bits_dataOffset =
    (tryToRead_2[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_2[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_2[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_2[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_2[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_2[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_2[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_2_bits_requestIndex =
    {2'h0, tryToRead_2[1]} | {1'h0, tryToRead_2[2], 1'h0} | (tryToRead_2[3] ? 3'h3 : 3'h0) | {tryToRead_2[4], 2'h0} | (tryToRead_2[5] ? 3'h5 : 3'h0) | (tryToRead_2[6] ? 3'h6 : 3'h0) | {3{tryToRead_2[7]}};
  wire [2:0] selectReq_2_bits_readLane =
    (tryToRead_2[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_2[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_2[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_2[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_2[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_2[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_2[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_2[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_2_bits_offset =
    (tryToRead_2[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_2[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_2[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_2[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_2[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_2[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_2[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_2[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_2_bits_vs =
    (tryToRead_2[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_2[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_2[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_2[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_2[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_2[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_2[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_2[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_2_valid =
    tryToRead_2[0] & input_0_valid_0 | tryToRead_2[1] & input_1_valid_0 | tryToRead_2[2] & input_2_valid_0 | tryToRead_2[3] & input_3_valid_0 | tryToRead_2[4] & input_4_valid_0 | tryToRead_2[5] & input_5_valid_0 | tryToRead_2[6]
    & input_6_valid_0 | tryToRead_2[7] & input_7_valid_0;
  wire       selectReq_2_ready =
    tryToRead_2[0] & input_0_ready_0 | tryToRead_2[1] & input_1_ready_0 | tryToRead_2[2] & input_2_ready_0 | tryToRead_2[3] & input_3_ready_0 | tryToRead_2[4] & input_4_ready_0 | tryToRead_2[5] & input_5_ready_0 | tryToRead_2[6]
    & input_6_ready_0 | tryToRead_2[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_3 = {inputSelect1H_1[3], inputSelect1H_0[3]};
  wire [1:0] tryToRead_lo_hi_3 = {inputSelect1H_3[3], inputSelect1H_2[3]};
  wire [3:0] tryToRead_lo_3 = {tryToRead_lo_hi_3, tryToRead_lo_lo_3};
  wire [1:0] tryToRead_hi_lo_3 = {inputSelect1H_5[3], inputSelect1H_4[3]};
  wire [1:0] tryToRead_hi_hi_3 = {inputSelect1H_7[3], inputSelect1H_6[3]};
  wire [3:0] tryToRead_hi_3 = {tryToRead_hi_hi_3, tryToRead_hi_lo_3};
  wire [7:0] tryToRead_3 = {tryToRead_hi_3, tryToRead_lo_3};
  wire       output_3_valid_0 = |tryToRead_3;
  wire [4:0] output_3_bits_vs_0 = selectReq_3_bits_vs;
  wire [1:0] output_3_bits_offset_0 = selectReq_3_bits_offset;
  wire [2:0] output_3_bits_writeIndex_0 = selectReq_3_bits_requestIndex;
  wire [1:0] output_3_bits_dataOffset_0 = selectReq_3_bits_dataOffset;
  assign selectReq_3_bits_dataOffset =
    (tryToRead_3[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_3[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_3[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_3[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_3[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_3[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_3[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_3_bits_requestIndex =
    {2'h0, tryToRead_3[1]} | {1'h0, tryToRead_3[2], 1'h0} | (tryToRead_3[3] ? 3'h3 : 3'h0) | {tryToRead_3[4], 2'h0} | (tryToRead_3[5] ? 3'h5 : 3'h0) | (tryToRead_3[6] ? 3'h6 : 3'h0) | {3{tryToRead_3[7]}};
  wire [2:0] selectReq_3_bits_readLane =
    (tryToRead_3[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_3[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_3[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_3[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_3[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_3[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_3[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_3[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_3_bits_offset =
    (tryToRead_3[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_3[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_3[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_3[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_3[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_3[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_3[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_3[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_3_bits_vs =
    (tryToRead_3[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_3[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_3[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_3[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_3[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_3[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_3[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_3[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_3_valid =
    tryToRead_3[0] & input_0_valid_0 | tryToRead_3[1] & input_1_valid_0 | tryToRead_3[2] & input_2_valid_0 | tryToRead_3[3] & input_3_valid_0 | tryToRead_3[4] & input_4_valid_0 | tryToRead_3[5] & input_5_valid_0 | tryToRead_3[6]
    & input_6_valid_0 | tryToRead_3[7] & input_7_valid_0;
  wire       selectReq_3_ready =
    tryToRead_3[0] & input_0_ready_0 | tryToRead_3[1] & input_1_ready_0 | tryToRead_3[2] & input_2_ready_0 | tryToRead_3[3] & input_3_ready_0 | tryToRead_3[4] & input_4_ready_0 | tryToRead_3[5] & input_5_ready_0 | tryToRead_3[6]
    & input_6_ready_0 | tryToRead_3[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_4 = {inputSelect1H_1[4], inputSelect1H_0[4]};
  wire [1:0] tryToRead_lo_hi_4 = {inputSelect1H_3[4], inputSelect1H_2[4]};
  wire [3:0] tryToRead_lo_4 = {tryToRead_lo_hi_4, tryToRead_lo_lo_4};
  wire [1:0] tryToRead_hi_lo_4 = {inputSelect1H_5[4], inputSelect1H_4[4]};
  wire [1:0] tryToRead_hi_hi_4 = {inputSelect1H_7[4], inputSelect1H_6[4]};
  wire [3:0] tryToRead_hi_4 = {tryToRead_hi_hi_4, tryToRead_hi_lo_4};
  wire [7:0] tryToRead_4 = {tryToRead_hi_4, tryToRead_lo_4};
  wire       output_4_valid_0 = |tryToRead_4;
  wire [4:0] output_4_bits_vs_0 = selectReq_4_bits_vs;
  wire [1:0] output_4_bits_offset_0 = selectReq_4_bits_offset;
  wire [2:0] output_4_bits_writeIndex_0 = selectReq_4_bits_requestIndex;
  wire [1:0] output_4_bits_dataOffset_0 = selectReq_4_bits_dataOffset;
  assign selectReq_4_bits_dataOffset =
    (tryToRead_4[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_4[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_4[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_4[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_4[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_4[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_4[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_4_bits_requestIndex =
    {2'h0, tryToRead_4[1]} | {1'h0, tryToRead_4[2], 1'h0} | (tryToRead_4[3] ? 3'h3 : 3'h0) | {tryToRead_4[4], 2'h0} | (tryToRead_4[5] ? 3'h5 : 3'h0) | (tryToRead_4[6] ? 3'h6 : 3'h0) | {3{tryToRead_4[7]}};
  wire [2:0] selectReq_4_bits_readLane =
    (tryToRead_4[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_4[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_4[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_4[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_4[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_4[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_4[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_4[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_4_bits_offset =
    (tryToRead_4[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_4[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_4[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_4[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_4[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_4[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_4[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_4[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_4_bits_vs =
    (tryToRead_4[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_4[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_4[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_4[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_4[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_4[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_4[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_4[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_4_valid =
    tryToRead_4[0] & input_0_valid_0 | tryToRead_4[1] & input_1_valid_0 | tryToRead_4[2] & input_2_valid_0 | tryToRead_4[3] & input_3_valid_0 | tryToRead_4[4] & input_4_valid_0 | tryToRead_4[5] & input_5_valid_0 | tryToRead_4[6]
    & input_6_valid_0 | tryToRead_4[7] & input_7_valid_0;
  wire       selectReq_4_ready =
    tryToRead_4[0] & input_0_ready_0 | tryToRead_4[1] & input_1_ready_0 | tryToRead_4[2] & input_2_ready_0 | tryToRead_4[3] & input_3_ready_0 | tryToRead_4[4] & input_4_ready_0 | tryToRead_4[5] & input_5_ready_0 | tryToRead_4[6]
    & input_6_ready_0 | tryToRead_4[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_5 = {inputSelect1H_1[5], inputSelect1H_0[5]};
  wire [1:0] tryToRead_lo_hi_5 = {inputSelect1H_3[5], inputSelect1H_2[5]};
  wire [3:0] tryToRead_lo_5 = {tryToRead_lo_hi_5, tryToRead_lo_lo_5};
  wire [1:0] tryToRead_hi_lo_5 = {inputSelect1H_5[5], inputSelect1H_4[5]};
  wire [1:0] tryToRead_hi_hi_5 = {inputSelect1H_7[5], inputSelect1H_6[5]};
  wire [3:0] tryToRead_hi_5 = {tryToRead_hi_hi_5, tryToRead_hi_lo_5};
  wire [7:0] tryToRead_5 = {tryToRead_hi_5, tryToRead_lo_5};
  wire       output_5_valid_0 = |tryToRead_5;
  wire [4:0] output_5_bits_vs_0 = selectReq_5_bits_vs;
  wire [1:0] output_5_bits_offset_0 = selectReq_5_bits_offset;
  wire [2:0] output_5_bits_writeIndex_0 = selectReq_5_bits_requestIndex;
  wire [1:0] output_5_bits_dataOffset_0 = selectReq_5_bits_dataOffset;
  assign selectReq_5_bits_dataOffset =
    (tryToRead_5[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_5[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_5[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_5[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_5[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_5[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_5[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_5_bits_requestIndex =
    {2'h0, tryToRead_5[1]} | {1'h0, tryToRead_5[2], 1'h0} | (tryToRead_5[3] ? 3'h3 : 3'h0) | {tryToRead_5[4], 2'h0} | (tryToRead_5[5] ? 3'h5 : 3'h0) | (tryToRead_5[6] ? 3'h6 : 3'h0) | {3{tryToRead_5[7]}};
  wire [2:0] selectReq_5_bits_readLane =
    (tryToRead_5[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_5[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_5[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_5[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_5[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_5[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_5[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_5[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_5_bits_offset =
    (tryToRead_5[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_5[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_5[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_5[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_5[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_5[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_5[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_5[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_5_bits_vs =
    (tryToRead_5[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_5[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_5[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_5[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_5[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_5[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_5[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_5[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_5_valid =
    tryToRead_5[0] & input_0_valid_0 | tryToRead_5[1] & input_1_valid_0 | tryToRead_5[2] & input_2_valid_0 | tryToRead_5[3] & input_3_valid_0 | tryToRead_5[4] & input_4_valid_0 | tryToRead_5[5] & input_5_valid_0 | tryToRead_5[6]
    & input_6_valid_0 | tryToRead_5[7] & input_7_valid_0;
  wire       selectReq_5_ready =
    tryToRead_5[0] & input_0_ready_0 | tryToRead_5[1] & input_1_ready_0 | tryToRead_5[2] & input_2_ready_0 | tryToRead_5[3] & input_3_ready_0 | tryToRead_5[4] & input_4_ready_0 | tryToRead_5[5] & input_5_ready_0 | tryToRead_5[6]
    & input_6_ready_0 | tryToRead_5[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_6 = {inputSelect1H_1[6], inputSelect1H_0[6]};
  wire [1:0] tryToRead_lo_hi_6 = {inputSelect1H_3[6], inputSelect1H_2[6]};
  wire [3:0] tryToRead_lo_6 = {tryToRead_lo_hi_6, tryToRead_lo_lo_6};
  wire [1:0] tryToRead_hi_lo_6 = {inputSelect1H_5[6], inputSelect1H_4[6]};
  wire [1:0] tryToRead_hi_hi_6 = {inputSelect1H_7[6], inputSelect1H_6[6]};
  wire [3:0] tryToRead_hi_6 = {tryToRead_hi_hi_6, tryToRead_hi_lo_6};
  wire [7:0] tryToRead_6 = {tryToRead_hi_6, tryToRead_lo_6};
  wire       output_6_valid_0 = |tryToRead_6;
  wire [4:0] output_6_bits_vs_0 = selectReq_6_bits_vs;
  wire [1:0] output_6_bits_offset_0 = selectReq_6_bits_offset;
  wire [2:0] output_6_bits_writeIndex_0 = selectReq_6_bits_requestIndex;
  wire [1:0] output_6_bits_dataOffset_0 = selectReq_6_bits_dataOffset;
  assign selectReq_6_bits_dataOffset =
    (tryToRead_6[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_6[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_6[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_6[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_6[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_6[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_6[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_6_bits_requestIndex =
    {2'h0, tryToRead_6[1]} | {1'h0, tryToRead_6[2], 1'h0} | (tryToRead_6[3] ? 3'h3 : 3'h0) | {tryToRead_6[4], 2'h0} | (tryToRead_6[5] ? 3'h5 : 3'h0) | (tryToRead_6[6] ? 3'h6 : 3'h0) | {3{tryToRead_6[7]}};
  wire [2:0] selectReq_6_bits_readLane =
    (tryToRead_6[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_6[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_6[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_6[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_6[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_6[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_6[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_6[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_6_bits_offset =
    (tryToRead_6[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_6[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_6[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_6[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_6[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_6[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_6[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_6[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_6_bits_vs =
    (tryToRead_6[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_6[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_6[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_6[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_6[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_6[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_6[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_6[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_6_valid =
    tryToRead_6[0] & input_0_valid_0 | tryToRead_6[1] & input_1_valid_0 | tryToRead_6[2] & input_2_valid_0 | tryToRead_6[3] & input_3_valid_0 | tryToRead_6[4] & input_4_valid_0 | tryToRead_6[5] & input_5_valid_0 | tryToRead_6[6]
    & input_6_valid_0 | tryToRead_6[7] & input_7_valid_0;
  wire       selectReq_6_ready =
    tryToRead_6[0] & input_0_ready_0 | tryToRead_6[1] & input_1_ready_0 | tryToRead_6[2] & input_2_ready_0 | tryToRead_6[3] & input_3_ready_0 | tryToRead_6[4] & input_4_ready_0 | tryToRead_6[5] & input_5_ready_0 | tryToRead_6[6]
    & input_6_ready_0 | tryToRead_6[7] & input_7_ready_0;
  wire [1:0] tryToRead_lo_lo_7 = {inputSelect1H_1[7], inputSelect1H_0[7]};
  wire [1:0] tryToRead_lo_hi_7 = {inputSelect1H_3[7], inputSelect1H_2[7]};
  wire [3:0] tryToRead_lo_7 = {tryToRead_lo_hi_7, tryToRead_lo_lo_7};
  wire [1:0] tryToRead_hi_lo_7 = {inputSelect1H_5[7], inputSelect1H_4[7]};
  wire [1:0] tryToRead_hi_hi_7 = {inputSelect1H_7[7], inputSelect1H_6[7]};
  wire [3:0] tryToRead_hi_7 = {tryToRead_hi_hi_7, tryToRead_hi_lo_7};
  wire [7:0] tryToRead_7 = {tryToRead_hi_7, tryToRead_lo_7};
  wire       output_7_valid_0 = |tryToRead_7;
  wire [4:0] output_7_bits_vs_0 = selectReq_7_bits_vs;
  wire [1:0] output_7_bits_offset_0 = selectReq_7_bits_offset;
  wire [2:0] output_7_bits_writeIndex_0 = selectReq_7_bits_requestIndex;
  wire [1:0] output_7_bits_dataOffset_0 = selectReq_7_bits_dataOffset;
  assign selectReq_7_bits_dataOffset =
    (tryToRead_7[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_7[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_7[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_7[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_7[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_7[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_7[7] ? input_7_bits_dataOffset_0 : 2'h0);
  assign selectReq_7_bits_requestIndex =
    {2'h0, tryToRead_7[1]} | {1'h0, tryToRead_7[2], 1'h0} | (tryToRead_7[3] ? 3'h3 : 3'h0) | {tryToRead_7[4], 2'h0} | (tryToRead_7[5] ? 3'h5 : 3'h0) | (tryToRead_7[6] ? 3'h6 : 3'h0) | {3{tryToRead_7[7]}};
  wire [2:0] selectReq_7_bits_readLane =
    (tryToRead_7[0] ? input_0_bits_readLane_0 : 3'h0) | (tryToRead_7[1] ? input_1_bits_readLane_0 : 3'h0) | (tryToRead_7[2] ? input_2_bits_readLane_0 : 3'h0) | (tryToRead_7[3] ? input_3_bits_readLane_0 : 3'h0)
    | (tryToRead_7[4] ? input_4_bits_readLane_0 : 3'h0) | (tryToRead_7[5] ? input_5_bits_readLane_0 : 3'h0) | (tryToRead_7[6] ? input_6_bits_readLane_0 : 3'h0) | (tryToRead_7[7] ? input_7_bits_readLane_0 : 3'h0);
  assign selectReq_7_bits_offset =
    (tryToRead_7[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_7[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_7[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_7[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_7[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_7[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_7[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_7[7] ? input_7_bits_offset_0 : 2'h0);
  assign selectReq_7_bits_vs =
    (tryToRead_7[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_7[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_7[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_7[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_7[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_7[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_7[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_7[7] ? input_7_bits_vs_0 : 5'h0);
  wire       selectReq_7_valid =
    tryToRead_7[0] & input_0_valid_0 | tryToRead_7[1] & input_1_valid_0 | tryToRead_7[2] & input_2_valid_0 | tryToRead_7[3] & input_3_valid_0 | tryToRead_7[4] & input_4_valid_0 | tryToRead_7[5] & input_5_valid_0 | tryToRead_7[6]
    & input_6_valid_0 | tryToRead_7[7] & input_7_valid_0;
  wire       selectReq_7_ready =
    tryToRead_7[0] & input_0_ready_0 | tryToRead_7[1] & input_1_ready_0 | tryToRead_7[2] & input_2_ready_0 | tryToRead_7[3] & input_3_ready_0 | tryToRead_7[4] & input_4_ready_0 | tryToRead_7[5] & input_5_ready_0 | tryToRead_7[6]
    & input_6_ready_0 | tryToRead_7[7] & input_7_ready_0;
  assign input_0_ready = input_0_ready_0;
  assign input_1_ready = input_1_ready_0;
  assign input_2_ready = input_2_ready_0;
  assign input_3_ready = input_3_ready_0;
  assign input_4_ready = input_4_ready_0;
  assign input_5_ready = input_5_ready_0;
  assign input_6_ready = input_6_ready_0;
  assign input_7_ready = input_7_ready_0;
  assign output_0_valid = output_0_valid_0;
  assign output_0_bits_vs = output_0_bits_vs_0;
  assign output_0_bits_offset = output_0_bits_offset_0;
  assign output_0_bits_writeIndex = output_0_bits_writeIndex_0;
  assign output_0_bits_dataOffset = output_0_bits_dataOffset_0;
  assign output_1_valid = output_1_valid_0;
  assign output_1_bits_vs = output_1_bits_vs_0;
  assign output_1_bits_offset = output_1_bits_offset_0;
  assign output_1_bits_writeIndex = output_1_bits_writeIndex_0;
  assign output_1_bits_dataOffset = output_1_bits_dataOffset_0;
  assign output_2_valid = output_2_valid_0;
  assign output_2_bits_vs = output_2_bits_vs_0;
  assign output_2_bits_offset = output_2_bits_offset_0;
  assign output_2_bits_writeIndex = output_2_bits_writeIndex_0;
  assign output_2_bits_dataOffset = output_2_bits_dataOffset_0;
  assign output_3_valid = output_3_valid_0;
  assign output_3_bits_vs = output_3_bits_vs_0;
  assign output_3_bits_offset = output_3_bits_offset_0;
  assign output_3_bits_writeIndex = output_3_bits_writeIndex_0;
  assign output_3_bits_dataOffset = output_3_bits_dataOffset_0;
  assign output_4_valid = output_4_valid_0;
  assign output_4_bits_vs = output_4_bits_vs_0;
  assign output_4_bits_offset = output_4_bits_offset_0;
  assign output_4_bits_writeIndex = output_4_bits_writeIndex_0;
  assign output_4_bits_dataOffset = output_4_bits_dataOffset_0;
  assign output_5_valid = output_5_valid_0;
  assign output_5_bits_vs = output_5_bits_vs_0;
  assign output_5_bits_offset = output_5_bits_offset_0;
  assign output_5_bits_writeIndex = output_5_bits_writeIndex_0;
  assign output_5_bits_dataOffset = output_5_bits_dataOffset_0;
  assign output_6_valid = output_6_valid_0;
  assign output_6_bits_vs = output_6_bits_vs_0;
  assign output_6_bits_offset = output_6_bits_offset_0;
  assign output_6_bits_writeIndex = output_6_bits_writeIndex_0;
  assign output_6_bits_dataOffset = output_6_bits_dataOffset_0;
  assign output_7_valid = output_7_valid_0;
  assign output_7_bits_vs = output_7_bits_vs_0;
  assign output_7_bits_offset = output_7_bits_offset_0;
  assign output_7_bits_writeIndex = output_7_bits_writeIndex_0;
  assign output_7_bits_dataOffset = output_7_bits_dataOffset_0;
endmodule

