
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskedLogic(
  input         clock,
                reset,
                requestIO_valid,
  input  [1:0]  requestIO_bits_tag,
  input  [31:0] requestIO_bits_src_0,
                requestIO_bits_src_1,
                requestIO_bits_src_2,
                requestIO_bits_src_3,
  input  [3:0]  requestIO_bits_opcode,
  output        responseIO_valid,
  output [1:0]  responseIO_bits_tag,
  output [31:0] responseIO_bits_data
);

  wire [31:0]  response_data;
  wire         requestIO_valid_0 = requestIO_valid;
  wire [1:0]   requestIO_bits_tag_0 = requestIO_bits_tag;
  wire [31:0]  requestIO_bits_src_0_0 = requestIO_bits_src_0;
  wire [31:0]  requestIO_bits_src_1_0 = requestIO_bits_src_1;
  wire [31:0]  requestIO_bits_src_2_0 = requestIO_bits_src_2;
  wire [31:0]  requestIO_bits_src_3_0 = requestIO_bits_src_3;
  wire [3:0]   requestIO_bits_opcode_0 = requestIO_bits_opcode;
  wire [1:0]   response_tag = 2'h0;
  wire         requestIO_ready = 1'h1;
  wire         responseIO_ready = 1'h1;
  wire         request_pipeResponse_valid;
  wire [1:0]   request_pipeResponse_bits_tag;
  wire [31:0]  request_pipeResponse_bits_data;
  reg  [1:0]   requestReg_tag;
  wire [1:0]   request_responseWire_tag = requestReg_tag;
  reg  [31:0]  requestReg_src_0;
  reg  [31:0]  requestReg_src_1;
  reg  [31:0]  requestReg_src_2;
  reg  [31:0]  requestReg_src_3;
  reg  [3:0]   requestReg_opcode;
  wire [3:0]   request_opcode = requestReg_opcode;
  reg          requestRegValid;
  wire         vfuRequestFire = requestRegValid;
  wire         request_responseValidWire = requestRegValid;
  wire [31:0]  request_responseWire_data = response_data;
  reg          request_pipeResponse_pipe_v;
  assign request_pipeResponse_valid = request_pipeResponse_pipe_v;
  reg  [1:0]   request_pipeResponse_pipe_b_tag;
  assign request_pipeResponse_bits_tag = request_pipeResponse_pipe_b_tag;
  reg  [31:0]  request_pipeResponse_pipe_b_data;
  assign request_pipeResponse_bits_data = request_pipeResponse_pipe_b_data;
  wire         responseIO_valid_0 = request_pipeResponse_valid;
  wire [1:0]   responseIO_bits_tag_0 = request_pipeResponse_bits_tag;
  wire [31:0]  responseIO_bits_data_0 = request_pipeResponse_bits_data;
  wire [63:0]  request_lo = {requestReg_src_1, requestReg_src_0};
  wire [63:0]  request_hi = {requestReg_src_3, requestReg_src_2};
  wire [129:0] request_hi_1 = {requestReg_tag, request_hi, request_lo};
  wire [31:0]  request_src_0 = request_hi_1[31:0];
  wire [31:0]  request_src_1 = request_hi_1[63:32];
  wire [31:0]  request_src_2 = request_hi_1[95:64];
  wire [31:0]  request_src_3 = request_hi_1[127:96];
  wire [1:0]   request_tag = request_hi_1[129:128];
  wire [4:0]   response_data_plaInput;
  wire [4:0]   response_data_invInputs = ~response_data_plaInput;
  wire         response_data_invMatrixOutputs;
  wire         response_data_andMatrixOutputs_andMatrixInput_0 = response_data_plaInput[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_1 = response_data_plaInput[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_3 = response_data_plaInput[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1 = response_data_plaInput[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_2 = response_data_plaInput[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_4 = response_data_plaInput[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2 = response_data_invInputs[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_1 = response_data_invInputs[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_2 = response_data_invInputs[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3 = response_data_invInputs[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_1 = response_data_invInputs[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_2 = response_data_invInputs[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4 = response_data_invInputs[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_1 = response_data_invInputs[4];
  wire [1:0]   response_data_andMatrixOutputs_lo = {response_data_andMatrixOutputs_andMatrixInput_2, response_data_andMatrixOutputs_andMatrixInput_3};
  wire [1:0]   response_data_andMatrixOutputs_hi = {response_data_andMatrixOutputs_andMatrixInput_0, response_data_andMatrixOutputs_andMatrixInput_1};
  wire         response_data_andMatrixOutputs_4_2 = &{response_data_andMatrixOutputs_hi, response_data_andMatrixOutputs_lo};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_1 = response_data_plaInput[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_2 = response_data_plaInput[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_1 = {response_data_andMatrixOutputs_andMatrixInput_2_1, response_data_andMatrixOutputs_andMatrixInput_3_1};
  wire [1:0]   response_data_andMatrixOutputs_hi_1 = {response_data_andMatrixOutputs_andMatrixInput_0_1, response_data_andMatrixOutputs_andMatrixInput_1_1};
  wire         response_data_andMatrixOutputs_1_2 = &{response_data_andMatrixOutputs_hi_1, response_data_andMatrixOutputs_lo_1};
  wire [1:0]   response_data_andMatrixOutputs_lo_2 = {response_data_andMatrixOutputs_andMatrixInput_2_2, response_data_andMatrixOutputs_andMatrixInput_3_2};
  wire [1:0]   response_data_andMatrixOutputs_hi_2 = {response_data_andMatrixOutputs_andMatrixInput_0_2, response_data_andMatrixOutputs_andMatrixInput_1_2};
  wire         response_data_andMatrixOutputs_3_2 = &{response_data_andMatrixOutputs_hi_2, response_data_andMatrixOutputs_lo_2};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_3 = response_data_invInputs[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_3 = response_data_invInputs[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_4 = response_data_invInputs[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_3 = response_data_plaInput[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_4 = response_data_plaInput[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_3 = {response_data_andMatrixOutputs_andMatrixInput_3_3, response_data_andMatrixOutputs_andMatrixInput_4};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi = {response_data_andMatrixOutputs_andMatrixInput_0_3, response_data_andMatrixOutputs_andMatrixInput_1_3};
  wire [2:0]   response_data_andMatrixOutputs_hi_3 = {response_data_andMatrixOutputs_hi_hi, response_data_andMatrixOutputs_andMatrixInput_2_3};
  wire         response_data_andMatrixOutputs_0_2 = &{response_data_andMatrixOutputs_hi_3, response_data_andMatrixOutputs_lo_3};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_4 = response_data_invInputs[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_4 = {response_data_andMatrixOutputs_andMatrixInput_3_4, response_data_andMatrixOutputs_andMatrixInput_4_1};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_1 = {response_data_andMatrixOutputs_andMatrixInput_0_4, response_data_andMatrixOutputs_andMatrixInput_1_4};
  wire [2:0]   response_data_andMatrixOutputs_hi_4 = {response_data_andMatrixOutputs_hi_hi_1, response_data_andMatrixOutputs_andMatrixInput_2_4};
  wire         response_data_andMatrixOutputs_2_2 = &{response_data_andMatrixOutputs_hi_4, response_data_andMatrixOutputs_lo_4};
  wire [1:0]   response_data_orMatrixOutputs_lo = {response_data_andMatrixOutputs_0_2, response_data_andMatrixOutputs_2_2};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi = {response_data_andMatrixOutputs_4_2, response_data_andMatrixOutputs_1_2};
  wire [2:0]   response_data_orMatrixOutputs_hi = {response_data_orMatrixOutputs_hi_hi, response_data_andMatrixOutputs_3_2};
  wire         response_data_orMatrixOutputs = |{response_data_orMatrixOutputs_hi, response_data_orMatrixOutputs_lo};
  assign response_data_invMatrixOutputs = response_data_orMatrixOutputs;
  wire         response_data_plaOutput = response_data_invMatrixOutputs;
  assign response_data_plaInput = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[0], request_src_1[0]};
  wire [4:0]   response_data_plaInput_1;
  wire [4:0]   response_data_invInputs_1 = ~response_data_plaInput_1;
  wire         response_data_invMatrixOutputs_1;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_5 = response_data_plaInput_1[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_6 = response_data_plaInput_1[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_8 = response_data_plaInput_1[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_5 = response_data_plaInput_1[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_7 = response_data_plaInput_1[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_9 = response_data_plaInput_1[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_5 = response_data_invInputs_1[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_6 = response_data_invInputs_1[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_7 = response_data_invInputs_1[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_5 = response_data_invInputs_1[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_6 = response_data_invInputs_1[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_7 = response_data_invInputs_1[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_2 = response_data_invInputs_1[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_3 = response_data_invInputs_1[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_5 = {response_data_andMatrixOutputs_andMatrixInput_2_5, response_data_andMatrixOutputs_andMatrixInput_3_5};
  wire [1:0]   response_data_andMatrixOutputs_hi_5 = {response_data_andMatrixOutputs_andMatrixInput_0_5, response_data_andMatrixOutputs_andMatrixInput_1_5};
  wire         response_data_andMatrixOutputs_4_2_1 = &{response_data_andMatrixOutputs_hi_5, response_data_andMatrixOutputs_lo_5};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_6 = response_data_plaInput_1[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_7 = response_data_plaInput_1[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_6 = {response_data_andMatrixOutputs_andMatrixInput_2_6, response_data_andMatrixOutputs_andMatrixInput_3_6};
  wire [1:0]   response_data_andMatrixOutputs_hi_6 = {response_data_andMatrixOutputs_andMatrixInput_0_6, response_data_andMatrixOutputs_andMatrixInput_1_6};
  wire         response_data_andMatrixOutputs_1_2_1 = &{response_data_andMatrixOutputs_hi_6, response_data_andMatrixOutputs_lo_6};
  wire [1:0]   response_data_andMatrixOutputs_lo_7 = {response_data_andMatrixOutputs_andMatrixInput_2_7, response_data_andMatrixOutputs_andMatrixInput_3_7};
  wire [1:0]   response_data_andMatrixOutputs_hi_7 = {response_data_andMatrixOutputs_andMatrixInput_0_7, response_data_andMatrixOutputs_andMatrixInput_1_7};
  wire         response_data_andMatrixOutputs_3_2_1 = &{response_data_andMatrixOutputs_hi_7, response_data_andMatrixOutputs_lo_7};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_8 = response_data_invInputs_1[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_8 = response_data_invInputs_1[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_9 = response_data_invInputs_1[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_8 = response_data_plaInput_1[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_9 = response_data_plaInput_1[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_8 = {response_data_andMatrixOutputs_andMatrixInput_3_8, response_data_andMatrixOutputs_andMatrixInput_4_2};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_2 = {response_data_andMatrixOutputs_andMatrixInput_0_8, response_data_andMatrixOutputs_andMatrixInput_1_8};
  wire [2:0]   response_data_andMatrixOutputs_hi_8 = {response_data_andMatrixOutputs_hi_hi_2, response_data_andMatrixOutputs_andMatrixInput_2_8};
  wire         response_data_andMatrixOutputs_0_2_1 = &{response_data_andMatrixOutputs_hi_8, response_data_andMatrixOutputs_lo_8};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_9 = response_data_invInputs_1[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_9 = {response_data_andMatrixOutputs_andMatrixInput_3_9, response_data_andMatrixOutputs_andMatrixInput_4_3};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_3 = {response_data_andMatrixOutputs_andMatrixInput_0_9, response_data_andMatrixOutputs_andMatrixInput_1_9};
  wire [2:0]   response_data_andMatrixOutputs_hi_9 = {response_data_andMatrixOutputs_hi_hi_3, response_data_andMatrixOutputs_andMatrixInput_2_9};
  wire         response_data_andMatrixOutputs_2_2_1 = &{response_data_andMatrixOutputs_hi_9, response_data_andMatrixOutputs_lo_9};
  wire [1:0]   response_data_orMatrixOutputs_lo_1 = {response_data_andMatrixOutputs_0_2_1, response_data_andMatrixOutputs_2_2_1};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_1 = {response_data_andMatrixOutputs_4_2_1, response_data_andMatrixOutputs_1_2_1};
  wire [2:0]   response_data_orMatrixOutputs_hi_1 = {response_data_orMatrixOutputs_hi_hi_1, response_data_andMatrixOutputs_3_2_1};
  wire         response_data_orMatrixOutputs_1 = |{response_data_orMatrixOutputs_hi_1, response_data_orMatrixOutputs_lo_1};
  assign response_data_invMatrixOutputs_1 = response_data_orMatrixOutputs_1;
  wire         response_data_plaOutput_1 = response_data_invMatrixOutputs_1;
  assign response_data_plaInput_1 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[1], request_src_1[1]};
  wire [4:0]   response_data_plaInput_2;
  wire [4:0]   response_data_invInputs_2 = ~response_data_plaInput_2;
  wire         response_data_invMatrixOutputs_2;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_10 = response_data_plaInput_2[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_11 = response_data_plaInput_2[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_13 = response_data_plaInput_2[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_10 = response_data_plaInput_2[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_12 = response_data_plaInput_2[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_14 = response_data_plaInput_2[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_10 = response_data_invInputs_2[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_11 = response_data_invInputs_2[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_12 = response_data_invInputs_2[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_10 = response_data_invInputs_2[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_11 = response_data_invInputs_2[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_12 = response_data_invInputs_2[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_4 = response_data_invInputs_2[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_5 = response_data_invInputs_2[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_10 = {response_data_andMatrixOutputs_andMatrixInput_2_10, response_data_andMatrixOutputs_andMatrixInput_3_10};
  wire [1:0]   response_data_andMatrixOutputs_hi_10 = {response_data_andMatrixOutputs_andMatrixInput_0_10, response_data_andMatrixOutputs_andMatrixInput_1_10};
  wire         response_data_andMatrixOutputs_4_2_2 = &{response_data_andMatrixOutputs_hi_10, response_data_andMatrixOutputs_lo_10};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_11 = response_data_plaInput_2[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_12 = response_data_plaInput_2[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_11 = {response_data_andMatrixOutputs_andMatrixInput_2_11, response_data_andMatrixOutputs_andMatrixInput_3_11};
  wire [1:0]   response_data_andMatrixOutputs_hi_11 = {response_data_andMatrixOutputs_andMatrixInput_0_11, response_data_andMatrixOutputs_andMatrixInput_1_11};
  wire         response_data_andMatrixOutputs_1_2_2 = &{response_data_andMatrixOutputs_hi_11, response_data_andMatrixOutputs_lo_11};
  wire [1:0]   response_data_andMatrixOutputs_lo_12 = {response_data_andMatrixOutputs_andMatrixInput_2_12, response_data_andMatrixOutputs_andMatrixInput_3_12};
  wire [1:0]   response_data_andMatrixOutputs_hi_12 = {response_data_andMatrixOutputs_andMatrixInput_0_12, response_data_andMatrixOutputs_andMatrixInput_1_12};
  wire         response_data_andMatrixOutputs_3_2_2 = &{response_data_andMatrixOutputs_hi_12, response_data_andMatrixOutputs_lo_12};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_13 = response_data_invInputs_2[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_13 = response_data_invInputs_2[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_14 = response_data_invInputs_2[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_13 = response_data_plaInput_2[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_14 = response_data_plaInput_2[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_13 = {response_data_andMatrixOutputs_andMatrixInput_3_13, response_data_andMatrixOutputs_andMatrixInput_4_4};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_4 = {response_data_andMatrixOutputs_andMatrixInput_0_13, response_data_andMatrixOutputs_andMatrixInput_1_13};
  wire [2:0]   response_data_andMatrixOutputs_hi_13 = {response_data_andMatrixOutputs_hi_hi_4, response_data_andMatrixOutputs_andMatrixInput_2_13};
  wire         response_data_andMatrixOutputs_0_2_2 = &{response_data_andMatrixOutputs_hi_13, response_data_andMatrixOutputs_lo_13};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_14 = response_data_invInputs_2[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_14 = {response_data_andMatrixOutputs_andMatrixInput_3_14, response_data_andMatrixOutputs_andMatrixInput_4_5};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_5 = {response_data_andMatrixOutputs_andMatrixInput_0_14, response_data_andMatrixOutputs_andMatrixInput_1_14};
  wire [2:0]   response_data_andMatrixOutputs_hi_14 = {response_data_andMatrixOutputs_hi_hi_5, response_data_andMatrixOutputs_andMatrixInput_2_14};
  wire         response_data_andMatrixOutputs_2_2_2 = &{response_data_andMatrixOutputs_hi_14, response_data_andMatrixOutputs_lo_14};
  wire [1:0]   response_data_orMatrixOutputs_lo_2 = {response_data_andMatrixOutputs_0_2_2, response_data_andMatrixOutputs_2_2_2};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_2 = {response_data_andMatrixOutputs_4_2_2, response_data_andMatrixOutputs_1_2_2};
  wire [2:0]   response_data_orMatrixOutputs_hi_2 = {response_data_orMatrixOutputs_hi_hi_2, response_data_andMatrixOutputs_3_2_2};
  wire         response_data_orMatrixOutputs_2 = |{response_data_orMatrixOutputs_hi_2, response_data_orMatrixOutputs_lo_2};
  assign response_data_invMatrixOutputs_2 = response_data_orMatrixOutputs_2;
  wire         response_data_plaOutput_2 = response_data_invMatrixOutputs_2;
  assign response_data_plaInput_2 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[2], request_src_1[2]};
  wire [4:0]   response_data_plaInput_3;
  wire [4:0]   response_data_invInputs_3 = ~response_data_plaInput_3;
  wire         response_data_invMatrixOutputs_3;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_15 = response_data_plaInput_3[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_16 = response_data_plaInput_3[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_18 = response_data_plaInput_3[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_15 = response_data_plaInput_3[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_17 = response_data_plaInput_3[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_19 = response_data_plaInput_3[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_15 = response_data_invInputs_3[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_16 = response_data_invInputs_3[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_17 = response_data_invInputs_3[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_15 = response_data_invInputs_3[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_16 = response_data_invInputs_3[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_17 = response_data_invInputs_3[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_6 = response_data_invInputs_3[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_7 = response_data_invInputs_3[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_15 = {response_data_andMatrixOutputs_andMatrixInput_2_15, response_data_andMatrixOutputs_andMatrixInput_3_15};
  wire [1:0]   response_data_andMatrixOutputs_hi_15 = {response_data_andMatrixOutputs_andMatrixInput_0_15, response_data_andMatrixOutputs_andMatrixInput_1_15};
  wire         response_data_andMatrixOutputs_4_2_3 = &{response_data_andMatrixOutputs_hi_15, response_data_andMatrixOutputs_lo_15};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_16 = response_data_plaInput_3[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_17 = response_data_plaInput_3[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_16 = {response_data_andMatrixOutputs_andMatrixInput_2_16, response_data_andMatrixOutputs_andMatrixInput_3_16};
  wire [1:0]   response_data_andMatrixOutputs_hi_16 = {response_data_andMatrixOutputs_andMatrixInput_0_16, response_data_andMatrixOutputs_andMatrixInput_1_16};
  wire         response_data_andMatrixOutputs_1_2_3 = &{response_data_andMatrixOutputs_hi_16, response_data_andMatrixOutputs_lo_16};
  wire [1:0]   response_data_andMatrixOutputs_lo_17 = {response_data_andMatrixOutputs_andMatrixInput_2_17, response_data_andMatrixOutputs_andMatrixInput_3_17};
  wire [1:0]   response_data_andMatrixOutputs_hi_17 = {response_data_andMatrixOutputs_andMatrixInput_0_17, response_data_andMatrixOutputs_andMatrixInput_1_17};
  wire         response_data_andMatrixOutputs_3_2_3 = &{response_data_andMatrixOutputs_hi_17, response_data_andMatrixOutputs_lo_17};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_18 = response_data_invInputs_3[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_18 = response_data_invInputs_3[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_19 = response_data_invInputs_3[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_18 = response_data_plaInput_3[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_19 = response_data_plaInput_3[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_18 = {response_data_andMatrixOutputs_andMatrixInput_3_18, response_data_andMatrixOutputs_andMatrixInput_4_6};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_6 = {response_data_andMatrixOutputs_andMatrixInput_0_18, response_data_andMatrixOutputs_andMatrixInput_1_18};
  wire [2:0]   response_data_andMatrixOutputs_hi_18 = {response_data_andMatrixOutputs_hi_hi_6, response_data_andMatrixOutputs_andMatrixInput_2_18};
  wire         response_data_andMatrixOutputs_0_2_3 = &{response_data_andMatrixOutputs_hi_18, response_data_andMatrixOutputs_lo_18};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_19 = response_data_invInputs_3[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_19 = {response_data_andMatrixOutputs_andMatrixInput_3_19, response_data_andMatrixOutputs_andMatrixInput_4_7};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_7 = {response_data_andMatrixOutputs_andMatrixInput_0_19, response_data_andMatrixOutputs_andMatrixInput_1_19};
  wire [2:0]   response_data_andMatrixOutputs_hi_19 = {response_data_andMatrixOutputs_hi_hi_7, response_data_andMatrixOutputs_andMatrixInput_2_19};
  wire         response_data_andMatrixOutputs_2_2_3 = &{response_data_andMatrixOutputs_hi_19, response_data_andMatrixOutputs_lo_19};
  wire [1:0]   response_data_orMatrixOutputs_lo_3 = {response_data_andMatrixOutputs_0_2_3, response_data_andMatrixOutputs_2_2_3};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_3 = {response_data_andMatrixOutputs_4_2_3, response_data_andMatrixOutputs_1_2_3};
  wire [2:0]   response_data_orMatrixOutputs_hi_3 = {response_data_orMatrixOutputs_hi_hi_3, response_data_andMatrixOutputs_3_2_3};
  wire         response_data_orMatrixOutputs_3 = |{response_data_orMatrixOutputs_hi_3, response_data_orMatrixOutputs_lo_3};
  assign response_data_invMatrixOutputs_3 = response_data_orMatrixOutputs_3;
  wire         response_data_plaOutput_3 = response_data_invMatrixOutputs_3;
  assign response_data_plaInput_3 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[3], request_src_1[3]};
  wire [4:0]   response_data_plaInput_4;
  wire [4:0]   response_data_invInputs_4 = ~response_data_plaInput_4;
  wire         response_data_invMatrixOutputs_4;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_20 = response_data_plaInput_4[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_21 = response_data_plaInput_4[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_23 = response_data_plaInput_4[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_20 = response_data_plaInput_4[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_22 = response_data_plaInput_4[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_24 = response_data_plaInput_4[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_20 = response_data_invInputs_4[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_21 = response_data_invInputs_4[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_22 = response_data_invInputs_4[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_20 = response_data_invInputs_4[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_21 = response_data_invInputs_4[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_22 = response_data_invInputs_4[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_8 = response_data_invInputs_4[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_9 = response_data_invInputs_4[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_20 = {response_data_andMatrixOutputs_andMatrixInput_2_20, response_data_andMatrixOutputs_andMatrixInput_3_20};
  wire [1:0]   response_data_andMatrixOutputs_hi_20 = {response_data_andMatrixOutputs_andMatrixInput_0_20, response_data_andMatrixOutputs_andMatrixInput_1_20};
  wire         response_data_andMatrixOutputs_4_2_4 = &{response_data_andMatrixOutputs_hi_20, response_data_andMatrixOutputs_lo_20};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_21 = response_data_plaInput_4[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_22 = response_data_plaInput_4[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_21 = {response_data_andMatrixOutputs_andMatrixInput_2_21, response_data_andMatrixOutputs_andMatrixInput_3_21};
  wire [1:0]   response_data_andMatrixOutputs_hi_21 = {response_data_andMatrixOutputs_andMatrixInput_0_21, response_data_andMatrixOutputs_andMatrixInput_1_21};
  wire         response_data_andMatrixOutputs_1_2_4 = &{response_data_andMatrixOutputs_hi_21, response_data_andMatrixOutputs_lo_21};
  wire [1:0]   response_data_andMatrixOutputs_lo_22 = {response_data_andMatrixOutputs_andMatrixInput_2_22, response_data_andMatrixOutputs_andMatrixInput_3_22};
  wire [1:0]   response_data_andMatrixOutputs_hi_22 = {response_data_andMatrixOutputs_andMatrixInput_0_22, response_data_andMatrixOutputs_andMatrixInput_1_22};
  wire         response_data_andMatrixOutputs_3_2_4 = &{response_data_andMatrixOutputs_hi_22, response_data_andMatrixOutputs_lo_22};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_23 = response_data_invInputs_4[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_23 = response_data_invInputs_4[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_24 = response_data_invInputs_4[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_23 = response_data_plaInput_4[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_24 = response_data_plaInput_4[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_23 = {response_data_andMatrixOutputs_andMatrixInput_3_23, response_data_andMatrixOutputs_andMatrixInput_4_8};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_8 = {response_data_andMatrixOutputs_andMatrixInput_0_23, response_data_andMatrixOutputs_andMatrixInput_1_23};
  wire [2:0]   response_data_andMatrixOutputs_hi_23 = {response_data_andMatrixOutputs_hi_hi_8, response_data_andMatrixOutputs_andMatrixInput_2_23};
  wire         response_data_andMatrixOutputs_0_2_4 = &{response_data_andMatrixOutputs_hi_23, response_data_andMatrixOutputs_lo_23};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_24 = response_data_invInputs_4[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_24 = {response_data_andMatrixOutputs_andMatrixInput_3_24, response_data_andMatrixOutputs_andMatrixInput_4_9};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_9 = {response_data_andMatrixOutputs_andMatrixInput_0_24, response_data_andMatrixOutputs_andMatrixInput_1_24};
  wire [2:0]   response_data_andMatrixOutputs_hi_24 = {response_data_andMatrixOutputs_hi_hi_9, response_data_andMatrixOutputs_andMatrixInput_2_24};
  wire         response_data_andMatrixOutputs_2_2_4 = &{response_data_andMatrixOutputs_hi_24, response_data_andMatrixOutputs_lo_24};
  wire [1:0]   response_data_orMatrixOutputs_lo_4 = {response_data_andMatrixOutputs_0_2_4, response_data_andMatrixOutputs_2_2_4};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_4 = {response_data_andMatrixOutputs_4_2_4, response_data_andMatrixOutputs_1_2_4};
  wire [2:0]   response_data_orMatrixOutputs_hi_4 = {response_data_orMatrixOutputs_hi_hi_4, response_data_andMatrixOutputs_3_2_4};
  wire         response_data_orMatrixOutputs_4 = |{response_data_orMatrixOutputs_hi_4, response_data_orMatrixOutputs_lo_4};
  assign response_data_invMatrixOutputs_4 = response_data_orMatrixOutputs_4;
  wire         response_data_plaOutput_4 = response_data_invMatrixOutputs_4;
  assign response_data_plaInput_4 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[4], request_src_1[4]};
  wire [4:0]   response_data_plaInput_5;
  wire [4:0]   response_data_invInputs_5 = ~response_data_plaInput_5;
  wire         response_data_invMatrixOutputs_5;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_25 = response_data_plaInput_5[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_26 = response_data_plaInput_5[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_28 = response_data_plaInput_5[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_25 = response_data_plaInput_5[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_27 = response_data_plaInput_5[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_29 = response_data_plaInput_5[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_25 = response_data_invInputs_5[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_26 = response_data_invInputs_5[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_27 = response_data_invInputs_5[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_25 = response_data_invInputs_5[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_26 = response_data_invInputs_5[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_27 = response_data_invInputs_5[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_10 = response_data_invInputs_5[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_11 = response_data_invInputs_5[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_25 = {response_data_andMatrixOutputs_andMatrixInput_2_25, response_data_andMatrixOutputs_andMatrixInput_3_25};
  wire [1:0]   response_data_andMatrixOutputs_hi_25 = {response_data_andMatrixOutputs_andMatrixInput_0_25, response_data_andMatrixOutputs_andMatrixInput_1_25};
  wire         response_data_andMatrixOutputs_4_2_5 = &{response_data_andMatrixOutputs_hi_25, response_data_andMatrixOutputs_lo_25};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_26 = response_data_plaInput_5[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_27 = response_data_plaInput_5[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_26 = {response_data_andMatrixOutputs_andMatrixInput_2_26, response_data_andMatrixOutputs_andMatrixInput_3_26};
  wire [1:0]   response_data_andMatrixOutputs_hi_26 = {response_data_andMatrixOutputs_andMatrixInput_0_26, response_data_andMatrixOutputs_andMatrixInput_1_26};
  wire         response_data_andMatrixOutputs_1_2_5 = &{response_data_andMatrixOutputs_hi_26, response_data_andMatrixOutputs_lo_26};
  wire [1:0]   response_data_andMatrixOutputs_lo_27 = {response_data_andMatrixOutputs_andMatrixInput_2_27, response_data_andMatrixOutputs_andMatrixInput_3_27};
  wire [1:0]   response_data_andMatrixOutputs_hi_27 = {response_data_andMatrixOutputs_andMatrixInput_0_27, response_data_andMatrixOutputs_andMatrixInput_1_27};
  wire         response_data_andMatrixOutputs_3_2_5 = &{response_data_andMatrixOutputs_hi_27, response_data_andMatrixOutputs_lo_27};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_28 = response_data_invInputs_5[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_28 = response_data_invInputs_5[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_29 = response_data_invInputs_5[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_28 = response_data_plaInput_5[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_29 = response_data_plaInput_5[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_28 = {response_data_andMatrixOutputs_andMatrixInput_3_28, response_data_andMatrixOutputs_andMatrixInput_4_10};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_10 = {response_data_andMatrixOutputs_andMatrixInput_0_28, response_data_andMatrixOutputs_andMatrixInput_1_28};
  wire [2:0]   response_data_andMatrixOutputs_hi_28 = {response_data_andMatrixOutputs_hi_hi_10, response_data_andMatrixOutputs_andMatrixInput_2_28};
  wire         response_data_andMatrixOutputs_0_2_5 = &{response_data_andMatrixOutputs_hi_28, response_data_andMatrixOutputs_lo_28};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_29 = response_data_invInputs_5[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_29 = {response_data_andMatrixOutputs_andMatrixInput_3_29, response_data_andMatrixOutputs_andMatrixInput_4_11};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_11 = {response_data_andMatrixOutputs_andMatrixInput_0_29, response_data_andMatrixOutputs_andMatrixInput_1_29};
  wire [2:0]   response_data_andMatrixOutputs_hi_29 = {response_data_andMatrixOutputs_hi_hi_11, response_data_andMatrixOutputs_andMatrixInput_2_29};
  wire         response_data_andMatrixOutputs_2_2_5 = &{response_data_andMatrixOutputs_hi_29, response_data_andMatrixOutputs_lo_29};
  wire [1:0]   response_data_orMatrixOutputs_lo_5 = {response_data_andMatrixOutputs_0_2_5, response_data_andMatrixOutputs_2_2_5};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_5 = {response_data_andMatrixOutputs_4_2_5, response_data_andMatrixOutputs_1_2_5};
  wire [2:0]   response_data_orMatrixOutputs_hi_5 = {response_data_orMatrixOutputs_hi_hi_5, response_data_andMatrixOutputs_3_2_5};
  wire         response_data_orMatrixOutputs_5 = |{response_data_orMatrixOutputs_hi_5, response_data_orMatrixOutputs_lo_5};
  assign response_data_invMatrixOutputs_5 = response_data_orMatrixOutputs_5;
  wire         response_data_plaOutput_5 = response_data_invMatrixOutputs_5;
  assign response_data_plaInput_5 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[5], request_src_1[5]};
  wire [4:0]   response_data_plaInput_6;
  wire [4:0]   response_data_invInputs_6 = ~response_data_plaInput_6;
  wire         response_data_invMatrixOutputs_6;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_30 = response_data_plaInput_6[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_31 = response_data_plaInput_6[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_33 = response_data_plaInput_6[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_30 = response_data_plaInput_6[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_32 = response_data_plaInput_6[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_34 = response_data_plaInput_6[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_30 = response_data_invInputs_6[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_31 = response_data_invInputs_6[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_32 = response_data_invInputs_6[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_30 = response_data_invInputs_6[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_31 = response_data_invInputs_6[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_32 = response_data_invInputs_6[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_12 = response_data_invInputs_6[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_13 = response_data_invInputs_6[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_30 = {response_data_andMatrixOutputs_andMatrixInput_2_30, response_data_andMatrixOutputs_andMatrixInput_3_30};
  wire [1:0]   response_data_andMatrixOutputs_hi_30 = {response_data_andMatrixOutputs_andMatrixInput_0_30, response_data_andMatrixOutputs_andMatrixInput_1_30};
  wire         response_data_andMatrixOutputs_4_2_6 = &{response_data_andMatrixOutputs_hi_30, response_data_andMatrixOutputs_lo_30};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_31 = response_data_plaInput_6[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_32 = response_data_plaInput_6[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_31 = {response_data_andMatrixOutputs_andMatrixInput_2_31, response_data_andMatrixOutputs_andMatrixInput_3_31};
  wire [1:0]   response_data_andMatrixOutputs_hi_31 = {response_data_andMatrixOutputs_andMatrixInput_0_31, response_data_andMatrixOutputs_andMatrixInput_1_31};
  wire         response_data_andMatrixOutputs_1_2_6 = &{response_data_andMatrixOutputs_hi_31, response_data_andMatrixOutputs_lo_31};
  wire [1:0]   response_data_andMatrixOutputs_lo_32 = {response_data_andMatrixOutputs_andMatrixInput_2_32, response_data_andMatrixOutputs_andMatrixInput_3_32};
  wire [1:0]   response_data_andMatrixOutputs_hi_32 = {response_data_andMatrixOutputs_andMatrixInput_0_32, response_data_andMatrixOutputs_andMatrixInput_1_32};
  wire         response_data_andMatrixOutputs_3_2_6 = &{response_data_andMatrixOutputs_hi_32, response_data_andMatrixOutputs_lo_32};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_33 = response_data_invInputs_6[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_33 = response_data_invInputs_6[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_34 = response_data_invInputs_6[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_33 = response_data_plaInput_6[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_34 = response_data_plaInput_6[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_33 = {response_data_andMatrixOutputs_andMatrixInput_3_33, response_data_andMatrixOutputs_andMatrixInput_4_12};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_12 = {response_data_andMatrixOutputs_andMatrixInput_0_33, response_data_andMatrixOutputs_andMatrixInput_1_33};
  wire [2:0]   response_data_andMatrixOutputs_hi_33 = {response_data_andMatrixOutputs_hi_hi_12, response_data_andMatrixOutputs_andMatrixInput_2_33};
  wire         response_data_andMatrixOutputs_0_2_6 = &{response_data_andMatrixOutputs_hi_33, response_data_andMatrixOutputs_lo_33};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_34 = response_data_invInputs_6[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_34 = {response_data_andMatrixOutputs_andMatrixInput_3_34, response_data_andMatrixOutputs_andMatrixInput_4_13};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_13 = {response_data_andMatrixOutputs_andMatrixInput_0_34, response_data_andMatrixOutputs_andMatrixInput_1_34};
  wire [2:0]   response_data_andMatrixOutputs_hi_34 = {response_data_andMatrixOutputs_hi_hi_13, response_data_andMatrixOutputs_andMatrixInput_2_34};
  wire         response_data_andMatrixOutputs_2_2_6 = &{response_data_andMatrixOutputs_hi_34, response_data_andMatrixOutputs_lo_34};
  wire [1:0]   response_data_orMatrixOutputs_lo_6 = {response_data_andMatrixOutputs_0_2_6, response_data_andMatrixOutputs_2_2_6};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_6 = {response_data_andMatrixOutputs_4_2_6, response_data_andMatrixOutputs_1_2_6};
  wire [2:0]   response_data_orMatrixOutputs_hi_6 = {response_data_orMatrixOutputs_hi_hi_6, response_data_andMatrixOutputs_3_2_6};
  wire         response_data_orMatrixOutputs_6 = |{response_data_orMatrixOutputs_hi_6, response_data_orMatrixOutputs_lo_6};
  assign response_data_invMatrixOutputs_6 = response_data_orMatrixOutputs_6;
  wire         response_data_plaOutput_6 = response_data_invMatrixOutputs_6;
  assign response_data_plaInput_6 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[6], request_src_1[6]};
  wire [4:0]   response_data_plaInput_7;
  wire [4:0]   response_data_invInputs_7 = ~response_data_plaInput_7;
  wire         response_data_invMatrixOutputs_7;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_35 = response_data_plaInput_7[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_36 = response_data_plaInput_7[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_38 = response_data_plaInput_7[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_35 = response_data_plaInput_7[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_37 = response_data_plaInput_7[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_39 = response_data_plaInput_7[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_35 = response_data_invInputs_7[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_36 = response_data_invInputs_7[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_37 = response_data_invInputs_7[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_35 = response_data_invInputs_7[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_36 = response_data_invInputs_7[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_37 = response_data_invInputs_7[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_14 = response_data_invInputs_7[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_15 = response_data_invInputs_7[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_35 = {response_data_andMatrixOutputs_andMatrixInput_2_35, response_data_andMatrixOutputs_andMatrixInput_3_35};
  wire [1:0]   response_data_andMatrixOutputs_hi_35 = {response_data_andMatrixOutputs_andMatrixInput_0_35, response_data_andMatrixOutputs_andMatrixInput_1_35};
  wire         response_data_andMatrixOutputs_4_2_7 = &{response_data_andMatrixOutputs_hi_35, response_data_andMatrixOutputs_lo_35};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_36 = response_data_plaInput_7[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_37 = response_data_plaInput_7[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_36 = {response_data_andMatrixOutputs_andMatrixInput_2_36, response_data_andMatrixOutputs_andMatrixInput_3_36};
  wire [1:0]   response_data_andMatrixOutputs_hi_36 = {response_data_andMatrixOutputs_andMatrixInput_0_36, response_data_andMatrixOutputs_andMatrixInput_1_36};
  wire         response_data_andMatrixOutputs_1_2_7 = &{response_data_andMatrixOutputs_hi_36, response_data_andMatrixOutputs_lo_36};
  wire [1:0]   response_data_andMatrixOutputs_lo_37 = {response_data_andMatrixOutputs_andMatrixInput_2_37, response_data_andMatrixOutputs_andMatrixInput_3_37};
  wire [1:0]   response_data_andMatrixOutputs_hi_37 = {response_data_andMatrixOutputs_andMatrixInput_0_37, response_data_andMatrixOutputs_andMatrixInput_1_37};
  wire         response_data_andMatrixOutputs_3_2_7 = &{response_data_andMatrixOutputs_hi_37, response_data_andMatrixOutputs_lo_37};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_38 = response_data_invInputs_7[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_38 = response_data_invInputs_7[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_39 = response_data_invInputs_7[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_38 = response_data_plaInput_7[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_39 = response_data_plaInput_7[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_38 = {response_data_andMatrixOutputs_andMatrixInput_3_38, response_data_andMatrixOutputs_andMatrixInput_4_14};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_14 = {response_data_andMatrixOutputs_andMatrixInput_0_38, response_data_andMatrixOutputs_andMatrixInput_1_38};
  wire [2:0]   response_data_andMatrixOutputs_hi_38 = {response_data_andMatrixOutputs_hi_hi_14, response_data_andMatrixOutputs_andMatrixInput_2_38};
  wire         response_data_andMatrixOutputs_0_2_7 = &{response_data_andMatrixOutputs_hi_38, response_data_andMatrixOutputs_lo_38};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_39 = response_data_invInputs_7[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_39 = {response_data_andMatrixOutputs_andMatrixInput_3_39, response_data_andMatrixOutputs_andMatrixInput_4_15};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_15 = {response_data_andMatrixOutputs_andMatrixInput_0_39, response_data_andMatrixOutputs_andMatrixInput_1_39};
  wire [2:0]   response_data_andMatrixOutputs_hi_39 = {response_data_andMatrixOutputs_hi_hi_15, response_data_andMatrixOutputs_andMatrixInput_2_39};
  wire         response_data_andMatrixOutputs_2_2_7 = &{response_data_andMatrixOutputs_hi_39, response_data_andMatrixOutputs_lo_39};
  wire [1:0]   response_data_orMatrixOutputs_lo_7 = {response_data_andMatrixOutputs_0_2_7, response_data_andMatrixOutputs_2_2_7};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_7 = {response_data_andMatrixOutputs_4_2_7, response_data_andMatrixOutputs_1_2_7};
  wire [2:0]   response_data_orMatrixOutputs_hi_7 = {response_data_orMatrixOutputs_hi_hi_7, response_data_andMatrixOutputs_3_2_7};
  wire         response_data_orMatrixOutputs_7 = |{response_data_orMatrixOutputs_hi_7, response_data_orMatrixOutputs_lo_7};
  assign response_data_invMatrixOutputs_7 = response_data_orMatrixOutputs_7;
  wire         response_data_plaOutput_7 = response_data_invMatrixOutputs_7;
  assign response_data_plaInput_7 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[7], request_src_1[7]};
  wire [4:0]   response_data_plaInput_8;
  wire [4:0]   response_data_invInputs_8 = ~response_data_plaInput_8;
  wire         response_data_invMatrixOutputs_8;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_40 = response_data_plaInput_8[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_41 = response_data_plaInput_8[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_43 = response_data_plaInput_8[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_40 = response_data_plaInput_8[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_42 = response_data_plaInput_8[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_44 = response_data_plaInput_8[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_40 = response_data_invInputs_8[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_41 = response_data_invInputs_8[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_42 = response_data_invInputs_8[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_40 = response_data_invInputs_8[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_41 = response_data_invInputs_8[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_42 = response_data_invInputs_8[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_16 = response_data_invInputs_8[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_17 = response_data_invInputs_8[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_40 = {response_data_andMatrixOutputs_andMatrixInput_2_40, response_data_andMatrixOutputs_andMatrixInput_3_40};
  wire [1:0]   response_data_andMatrixOutputs_hi_40 = {response_data_andMatrixOutputs_andMatrixInput_0_40, response_data_andMatrixOutputs_andMatrixInput_1_40};
  wire         response_data_andMatrixOutputs_4_2_8 = &{response_data_andMatrixOutputs_hi_40, response_data_andMatrixOutputs_lo_40};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_41 = response_data_plaInput_8[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_42 = response_data_plaInput_8[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_41 = {response_data_andMatrixOutputs_andMatrixInput_2_41, response_data_andMatrixOutputs_andMatrixInput_3_41};
  wire [1:0]   response_data_andMatrixOutputs_hi_41 = {response_data_andMatrixOutputs_andMatrixInput_0_41, response_data_andMatrixOutputs_andMatrixInput_1_41};
  wire         response_data_andMatrixOutputs_1_2_8 = &{response_data_andMatrixOutputs_hi_41, response_data_andMatrixOutputs_lo_41};
  wire [1:0]   response_data_andMatrixOutputs_lo_42 = {response_data_andMatrixOutputs_andMatrixInput_2_42, response_data_andMatrixOutputs_andMatrixInput_3_42};
  wire [1:0]   response_data_andMatrixOutputs_hi_42 = {response_data_andMatrixOutputs_andMatrixInput_0_42, response_data_andMatrixOutputs_andMatrixInput_1_42};
  wire         response_data_andMatrixOutputs_3_2_8 = &{response_data_andMatrixOutputs_hi_42, response_data_andMatrixOutputs_lo_42};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_43 = response_data_invInputs_8[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_43 = response_data_invInputs_8[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_44 = response_data_invInputs_8[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_43 = response_data_plaInput_8[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_44 = response_data_plaInput_8[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_43 = {response_data_andMatrixOutputs_andMatrixInput_3_43, response_data_andMatrixOutputs_andMatrixInput_4_16};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_16 = {response_data_andMatrixOutputs_andMatrixInput_0_43, response_data_andMatrixOutputs_andMatrixInput_1_43};
  wire [2:0]   response_data_andMatrixOutputs_hi_43 = {response_data_andMatrixOutputs_hi_hi_16, response_data_andMatrixOutputs_andMatrixInput_2_43};
  wire         response_data_andMatrixOutputs_0_2_8 = &{response_data_andMatrixOutputs_hi_43, response_data_andMatrixOutputs_lo_43};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_44 = response_data_invInputs_8[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_44 = {response_data_andMatrixOutputs_andMatrixInput_3_44, response_data_andMatrixOutputs_andMatrixInput_4_17};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_17 = {response_data_andMatrixOutputs_andMatrixInput_0_44, response_data_andMatrixOutputs_andMatrixInput_1_44};
  wire [2:0]   response_data_andMatrixOutputs_hi_44 = {response_data_andMatrixOutputs_hi_hi_17, response_data_andMatrixOutputs_andMatrixInput_2_44};
  wire         response_data_andMatrixOutputs_2_2_8 = &{response_data_andMatrixOutputs_hi_44, response_data_andMatrixOutputs_lo_44};
  wire [1:0]   response_data_orMatrixOutputs_lo_8 = {response_data_andMatrixOutputs_0_2_8, response_data_andMatrixOutputs_2_2_8};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_8 = {response_data_andMatrixOutputs_4_2_8, response_data_andMatrixOutputs_1_2_8};
  wire [2:0]   response_data_orMatrixOutputs_hi_8 = {response_data_orMatrixOutputs_hi_hi_8, response_data_andMatrixOutputs_3_2_8};
  wire         response_data_orMatrixOutputs_8 = |{response_data_orMatrixOutputs_hi_8, response_data_orMatrixOutputs_lo_8};
  assign response_data_invMatrixOutputs_8 = response_data_orMatrixOutputs_8;
  wire         response_data_plaOutput_8 = response_data_invMatrixOutputs_8;
  assign response_data_plaInput_8 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[8], request_src_1[8]};
  wire [4:0]   response_data_plaInput_9;
  wire [4:0]   response_data_invInputs_9 = ~response_data_plaInput_9;
  wire         response_data_invMatrixOutputs_9;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_45 = response_data_plaInput_9[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_46 = response_data_plaInput_9[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_48 = response_data_plaInput_9[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_45 = response_data_plaInput_9[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_47 = response_data_plaInput_9[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_49 = response_data_plaInput_9[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_45 = response_data_invInputs_9[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_46 = response_data_invInputs_9[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_47 = response_data_invInputs_9[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_45 = response_data_invInputs_9[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_46 = response_data_invInputs_9[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_47 = response_data_invInputs_9[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_18 = response_data_invInputs_9[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_19 = response_data_invInputs_9[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_45 = {response_data_andMatrixOutputs_andMatrixInput_2_45, response_data_andMatrixOutputs_andMatrixInput_3_45};
  wire [1:0]   response_data_andMatrixOutputs_hi_45 = {response_data_andMatrixOutputs_andMatrixInput_0_45, response_data_andMatrixOutputs_andMatrixInput_1_45};
  wire         response_data_andMatrixOutputs_4_2_9 = &{response_data_andMatrixOutputs_hi_45, response_data_andMatrixOutputs_lo_45};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_46 = response_data_plaInput_9[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_47 = response_data_plaInput_9[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_46 = {response_data_andMatrixOutputs_andMatrixInput_2_46, response_data_andMatrixOutputs_andMatrixInput_3_46};
  wire [1:0]   response_data_andMatrixOutputs_hi_46 = {response_data_andMatrixOutputs_andMatrixInput_0_46, response_data_andMatrixOutputs_andMatrixInput_1_46};
  wire         response_data_andMatrixOutputs_1_2_9 = &{response_data_andMatrixOutputs_hi_46, response_data_andMatrixOutputs_lo_46};
  wire [1:0]   response_data_andMatrixOutputs_lo_47 = {response_data_andMatrixOutputs_andMatrixInput_2_47, response_data_andMatrixOutputs_andMatrixInput_3_47};
  wire [1:0]   response_data_andMatrixOutputs_hi_47 = {response_data_andMatrixOutputs_andMatrixInput_0_47, response_data_andMatrixOutputs_andMatrixInput_1_47};
  wire         response_data_andMatrixOutputs_3_2_9 = &{response_data_andMatrixOutputs_hi_47, response_data_andMatrixOutputs_lo_47};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_48 = response_data_invInputs_9[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_48 = response_data_invInputs_9[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_49 = response_data_invInputs_9[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_48 = response_data_plaInput_9[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_49 = response_data_plaInput_9[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_48 = {response_data_andMatrixOutputs_andMatrixInput_3_48, response_data_andMatrixOutputs_andMatrixInput_4_18};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_18 = {response_data_andMatrixOutputs_andMatrixInput_0_48, response_data_andMatrixOutputs_andMatrixInput_1_48};
  wire [2:0]   response_data_andMatrixOutputs_hi_48 = {response_data_andMatrixOutputs_hi_hi_18, response_data_andMatrixOutputs_andMatrixInput_2_48};
  wire         response_data_andMatrixOutputs_0_2_9 = &{response_data_andMatrixOutputs_hi_48, response_data_andMatrixOutputs_lo_48};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_49 = response_data_invInputs_9[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_49 = {response_data_andMatrixOutputs_andMatrixInput_3_49, response_data_andMatrixOutputs_andMatrixInput_4_19};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_19 = {response_data_andMatrixOutputs_andMatrixInput_0_49, response_data_andMatrixOutputs_andMatrixInput_1_49};
  wire [2:0]   response_data_andMatrixOutputs_hi_49 = {response_data_andMatrixOutputs_hi_hi_19, response_data_andMatrixOutputs_andMatrixInput_2_49};
  wire         response_data_andMatrixOutputs_2_2_9 = &{response_data_andMatrixOutputs_hi_49, response_data_andMatrixOutputs_lo_49};
  wire [1:0]   response_data_orMatrixOutputs_lo_9 = {response_data_andMatrixOutputs_0_2_9, response_data_andMatrixOutputs_2_2_9};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_9 = {response_data_andMatrixOutputs_4_2_9, response_data_andMatrixOutputs_1_2_9};
  wire [2:0]   response_data_orMatrixOutputs_hi_9 = {response_data_orMatrixOutputs_hi_hi_9, response_data_andMatrixOutputs_3_2_9};
  wire         response_data_orMatrixOutputs_9 = |{response_data_orMatrixOutputs_hi_9, response_data_orMatrixOutputs_lo_9};
  assign response_data_invMatrixOutputs_9 = response_data_orMatrixOutputs_9;
  wire         response_data_plaOutput_9 = response_data_invMatrixOutputs_9;
  assign response_data_plaInput_9 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[9], request_src_1[9]};
  wire [4:0]   response_data_plaInput_10;
  wire [4:0]   response_data_invInputs_10 = ~response_data_plaInput_10;
  wire         response_data_invMatrixOutputs_10;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_50 = response_data_plaInput_10[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_51 = response_data_plaInput_10[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_53 = response_data_plaInput_10[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_50 = response_data_plaInput_10[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_52 = response_data_plaInput_10[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_54 = response_data_plaInput_10[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_50 = response_data_invInputs_10[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_51 = response_data_invInputs_10[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_52 = response_data_invInputs_10[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_50 = response_data_invInputs_10[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_51 = response_data_invInputs_10[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_52 = response_data_invInputs_10[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_20 = response_data_invInputs_10[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_21 = response_data_invInputs_10[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_50 = {response_data_andMatrixOutputs_andMatrixInput_2_50, response_data_andMatrixOutputs_andMatrixInput_3_50};
  wire [1:0]   response_data_andMatrixOutputs_hi_50 = {response_data_andMatrixOutputs_andMatrixInput_0_50, response_data_andMatrixOutputs_andMatrixInput_1_50};
  wire         response_data_andMatrixOutputs_4_2_10 = &{response_data_andMatrixOutputs_hi_50, response_data_andMatrixOutputs_lo_50};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_51 = response_data_plaInput_10[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_52 = response_data_plaInput_10[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_51 = {response_data_andMatrixOutputs_andMatrixInput_2_51, response_data_andMatrixOutputs_andMatrixInput_3_51};
  wire [1:0]   response_data_andMatrixOutputs_hi_51 = {response_data_andMatrixOutputs_andMatrixInput_0_51, response_data_andMatrixOutputs_andMatrixInput_1_51};
  wire         response_data_andMatrixOutputs_1_2_10 = &{response_data_andMatrixOutputs_hi_51, response_data_andMatrixOutputs_lo_51};
  wire [1:0]   response_data_andMatrixOutputs_lo_52 = {response_data_andMatrixOutputs_andMatrixInput_2_52, response_data_andMatrixOutputs_andMatrixInput_3_52};
  wire [1:0]   response_data_andMatrixOutputs_hi_52 = {response_data_andMatrixOutputs_andMatrixInput_0_52, response_data_andMatrixOutputs_andMatrixInput_1_52};
  wire         response_data_andMatrixOutputs_3_2_10 = &{response_data_andMatrixOutputs_hi_52, response_data_andMatrixOutputs_lo_52};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_53 = response_data_invInputs_10[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_53 = response_data_invInputs_10[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_54 = response_data_invInputs_10[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_53 = response_data_plaInput_10[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_54 = response_data_plaInput_10[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_53 = {response_data_andMatrixOutputs_andMatrixInput_3_53, response_data_andMatrixOutputs_andMatrixInput_4_20};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_20 = {response_data_andMatrixOutputs_andMatrixInput_0_53, response_data_andMatrixOutputs_andMatrixInput_1_53};
  wire [2:0]   response_data_andMatrixOutputs_hi_53 = {response_data_andMatrixOutputs_hi_hi_20, response_data_andMatrixOutputs_andMatrixInput_2_53};
  wire         response_data_andMatrixOutputs_0_2_10 = &{response_data_andMatrixOutputs_hi_53, response_data_andMatrixOutputs_lo_53};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_54 = response_data_invInputs_10[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_54 = {response_data_andMatrixOutputs_andMatrixInput_3_54, response_data_andMatrixOutputs_andMatrixInput_4_21};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_21 = {response_data_andMatrixOutputs_andMatrixInput_0_54, response_data_andMatrixOutputs_andMatrixInput_1_54};
  wire [2:0]   response_data_andMatrixOutputs_hi_54 = {response_data_andMatrixOutputs_hi_hi_21, response_data_andMatrixOutputs_andMatrixInput_2_54};
  wire         response_data_andMatrixOutputs_2_2_10 = &{response_data_andMatrixOutputs_hi_54, response_data_andMatrixOutputs_lo_54};
  wire [1:0]   response_data_orMatrixOutputs_lo_10 = {response_data_andMatrixOutputs_0_2_10, response_data_andMatrixOutputs_2_2_10};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_10 = {response_data_andMatrixOutputs_4_2_10, response_data_andMatrixOutputs_1_2_10};
  wire [2:0]   response_data_orMatrixOutputs_hi_10 = {response_data_orMatrixOutputs_hi_hi_10, response_data_andMatrixOutputs_3_2_10};
  wire         response_data_orMatrixOutputs_10 = |{response_data_orMatrixOutputs_hi_10, response_data_orMatrixOutputs_lo_10};
  assign response_data_invMatrixOutputs_10 = response_data_orMatrixOutputs_10;
  wire         response_data_plaOutput_10 = response_data_invMatrixOutputs_10;
  assign response_data_plaInput_10 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[10], request_src_1[10]};
  wire [4:0]   response_data_plaInput_11;
  wire [4:0]   response_data_invInputs_11 = ~response_data_plaInput_11;
  wire         response_data_invMatrixOutputs_11;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_55 = response_data_plaInput_11[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_56 = response_data_plaInput_11[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_58 = response_data_plaInput_11[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_55 = response_data_plaInput_11[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_57 = response_data_plaInput_11[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_59 = response_data_plaInput_11[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_55 = response_data_invInputs_11[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_56 = response_data_invInputs_11[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_57 = response_data_invInputs_11[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_55 = response_data_invInputs_11[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_56 = response_data_invInputs_11[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_57 = response_data_invInputs_11[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_22 = response_data_invInputs_11[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_23 = response_data_invInputs_11[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_55 = {response_data_andMatrixOutputs_andMatrixInput_2_55, response_data_andMatrixOutputs_andMatrixInput_3_55};
  wire [1:0]   response_data_andMatrixOutputs_hi_55 = {response_data_andMatrixOutputs_andMatrixInput_0_55, response_data_andMatrixOutputs_andMatrixInput_1_55};
  wire         response_data_andMatrixOutputs_4_2_11 = &{response_data_andMatrixOutputs_hi_55, response_data_andMatrixOutputs_lo_55};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_56 = response_data_plaInput_11[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_57 = response_data_plaInput_11[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_56 = {response_data_andMatrixOutputs_andMatrixInput_2_56, response_data_andMatrixOutputs_andMatrixInput_3_56};
  wire [1:0]   response_data_andMatrixOutputs_hi_56 = {response_data_andMatrixOutputs_andMatrixInput_0_56, response_data_andMatrixOutputs_andMatrixInput_1_56};
  wire         response_data_andMatrixOutputs_1_2_11 = &{response_data_andMatrixOutputs_hi_56, response_data_andMatrixOutputs_lo_56};
  wire [1:0]   response_data_andMatrixOutputs_lo_57 = {response_data_andMatrixOutputs_andMatrixInput_2_57, response_data_andMatrixOutputs_andMatrixInput_3_57};
  wire [1:0]   response_data_andMatrixOutputs_hi_57 = {response_data_andMatrixOutputs_andMatrixInput_0_57, response_data_andMatrixOutputs_andMatrixInput_1_57};
  wire         response_data_andMatrixOutputs_3_2_11 = &{response_data_andMatrixOutputs_hi_57, response_data_andMatrixOutputs_lo_57};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_58 = response_data_invInputs_11[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_58 = response_data_invInputs_11[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_59 = response_data_invInputs_11[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_58 = response_data_plaInput_11[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_59 = response_data_plaInput_11[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_58 = {response_data_andMatrixOutputs_andMatrixInput_3_58, response_data_andMatrixOutputs_andMatrixInput_4_22};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_22 = {response_data_andMatrixOutputs_andMatrixInput_0_58, response_data_andMatrixOutputs_andMatrixInput_1_58};
  wire [2:0]   response_data_andMatrixOutputs_hi_58 = {response_data_andMatrixOutputs_hi_hi_22, response_data_andMatrixOutputs_andMatrixInput_2_58};
  wire         response_data_andMatrixOutputs_0_2_11 = &{response_data_andMatrixOutputs_hi_58, response_data_andMatrixOutputs_lo_58};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_59 = response_data_invInputs_11[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_59 = {response_data_andMatrixOutputs_andMatrixInput_3_59, response_data_andMatrixOutputs_andMatrixInput_4_23};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_23 = {response_data_andMatrixOutputs_andMatrixInput_0_59, response_data_andMatrixOutputs_andMatrixInput_1_59};
  wire [2:0]   response_data_andMatrixOutputs_hi_59 = {response_data_andMatrixOutputs_hi_hi_23, response_data_andMatrixOutputs_andMatrixInput_2_59};
  wire         response_data_andMatrixOutputs_2_2_11 = &{response_data_andMatrixOutputs_hi_59, response_data_andMatrixOutputs_lo_59};
  wire [1:0]   response_data_orMatrixOutputs_lo_11 = {response_data_andMatrixOutputs_0_2_11, response_data_andMatrixOutputs_2_2_11};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_11 = {response_data_andMatrixOutputs_4_2_11, response_data_andMatrixOutputs_1_2_11};
  wire [2:0]   response_data_orMatrixOutputs_hi_11 = {response_data_orMatrixOutputs_hi_hi_11, response_data_andMatrixOutputs_3_2_11};
  wire         response_data_orMatrixOutputs_11 = |{response_data_orMatrixOutputs_hi_11, response_data_orMatrixOutputs_lo_11};
  assign response_data_invMatrixOutputs_11 = response_data_orMatrixOutputs_11;
  wire         response_data_plaOutput_11 = response_data_invMatrixOutputs_11;
  assign response_data_plaInput_11 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[11], request_src_1[11]};
  wire [4:0]   response_data_plaInput_12;
  wire [4:0]   response_data_invInputs_12 = ~response_data_plaInput_12;
  wire         response_data_invMatrixOutputs_12;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_60 = response_data_plaInput_12[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_61 = response_data_plaInput_12[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_63 = response_data_plaInput_12[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_60 = response_data_plaInput_12[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_62 = response_data_plaInput_12[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_64 = response_data_plaInput_12[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_60 = response_data_invInputs_12[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_61 = response_data_invInputs_12[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_62 = response_data_invInputs_12[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_60 = response_data_invInputs_12[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_61 = response_data_invInputs_12[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_62 = response_data_invInputs_12[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_24 = response_data_invInputs_12[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_25 = response_data_invInputs_12[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_60 = {response_data_andMatrixOutputs_andMatrixInput_2_60, response_data_andMatrixOutputs_andMatrixInput_3_60};
  wire [1:0]   response_data_andMatrixOutputs_hi_60 = {response_data_andMatrixOutputs_andMatrixInput_0_60, response_data_andMatrixOutputs_andMatrixInput_1_60};
  wire         response_data_andMatrixOutputs_4_2_12 = &{response_data_andMatrixOutputs_hi_60, response_data_andMatrixOutputs_lo_60};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_61 = response_data_plaInput_12[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_62 = response_data_plaInput_12[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_61 = {response_data_andMatrixOutputs_andMatrixInput_2_61, response_data_andMatrixOutputs_andMatrixInput_3_61};
  wire [1:0]   response_data_andMatrixOutputs_hi_61 = {response_data_andMatrixOutputs_andMatrixInput_0_61, response_data_andMatrixOutputs_andMatrixInput_1_61};
  wire         response_data_andMatrixOutputs_1_2_12 = &{response_data_andMatrixOutputs_hi_61, response_data_andMatrixOutputs_lo_61};
  wire [1:0]   response_data_andMatrixOutputs_lo_62 = {response_data_andMatrixOutputs_andMatrixInput_2_62, response_data_andMatrixOutputs_andMatrixInput_3_62};
  wire [1:0]   response_data_andMatrixOutputs_hi_62 = {response_data_andMatrixOutputs_andMatrixInput_0_62, response_data_andMatrixOutputs_andMatrixInput_1_62};
  wire         response_data_andMatrixOutputs_3_2_12 = &{response_data_andMatrixOutputs_hi_62, response_data_andMatrixOutputs_lo_62};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_63 = response_data_invInputs_12[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_63 = response_data_invInputs_12[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_64 = response_data_invInputs_12[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_63 = response_data_plaInput_12[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_64 = response_data_plaInput_12[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_63 = {response_data_andMatrixOutputs_andMatrixInput_3_63, response_data_andMatrixOutputs_andMatrixInput_4_24};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_24 = {response_data_andMatrixOutputs_andMatrixInput_0_63, response_data_andMatrixOutputs_andMatrixInput_1_63};
  wire [2:0]   response_data_andMatrixOutputs_hi_63 = {response_data_andMatrixOutputs_hi_hi_24, response_data_andMatrixOutputs_andMatrixInput_2_63};
  wire         response_data_andMatrixOutputs_0_2_12 = &{response_data_andMatrixOutputs_hi_63, response_data_andMatrixOutputs_lo_63};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_64 = response_data_invInputs_12[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_64 = {response_data_andMatrixOutputs_andMatrixInput_3_64, response_data_andMatrixOutputs_andMatrixInput_4_25};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_25 = {response_data_andMatrixOutputs_andMatrixInput_0_64, response_data_andMatrixOutputs_andMatrixInput_1_64};
  wire [2:0]   response_data_andMatrixOutputs_hi_64 = {response_data_andMatrixOutputs_hi_hi_25, response_data_andMatrixOutputs_andMatrixInput_2_64};
  wire         response_data_andMatrixOutputs_2_2_12 = &{response_data_andMatrixOutputs_hi_64, response_data_andMatrixOutputs_lo_64};
  wire [1:0]   response_data_orMatrixOutputs_lo_12 = {response_data_andMatrixOutputs_0_2_12, response_data_andMatrixOutputs_2_2_12};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_12 = {response_data_andMatrixOutputs_4_2_12, response_data_andMatrixOutputs_1_2_12};
  wire [2:0]   response_data_orMatrixOutputs_hi_12 = {response_data_orMatrixOutputs_hi_hi_12, response_data_andMatrixOutputs_3_2_12};
  wire         response_data_orMatrixOutputs_12 = |{response_data_orMatrixOutputs_hi_12, response_data_orMatrixOutputs_lo_12};
  assign response_data_invMatrixOutputs_12 = response_data_orMatrixOutputs_12;
  wire         response_data_plaOutput_12 = response_data_invMatrixOutputs_12;
  assign response_data_plaInput_12 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[12], request_src_1[12]};
  wire [4:0]   response_data_plaInput_13;
  wire [4:0]   response_data_invInputs_13 = ~response_data_plaInput_13;
  wire         response_data_invMatrixOutputs_13;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_65 = response_data_plaInput_13[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_66 = response_data_plaInput_13[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_68 = response_data_plaInput_13[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_65 = response_data_plaInput_13[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_67 = response_data_plaInput_13[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_69 = response_data_plaInput_13[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_65 = response_data_invInputs_13[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_66 = response_data_invInputs_13[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_67 = response_data_invInputs_13[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_65 = response_data_invInputs_13[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_66 = response_data_invInputs_13[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_67 = response_data_invInputs_13[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_26 = response_data_invInputs_13[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_27 = response_data_invInputs_13[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_65 = {response_data_andMatrixOutputs_andMatrixInput_2_65, response_data_andMatrixOutputs_andMatrixInput_3_65};
  wire [1:0]   response_data_andMatrixOutputs_hi_65 = {response_data_andMatrixOutputs_andMatrixInput_0_65, response_data_andMatrixOutputs_andMatrixInput_1_65};
  wire         response_data_andMatrixOutputs_4_2_13 = &{response_data_andMatrixOutputs_hi_65, response_data_andMatrixOutputs_lo_65};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_66 = response_data_plaInput_13[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_67 = response_data_plaInput_13[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_66 = {response_data_andMatrixOutputs_andMatrixInput_2_66, response_data_andMatrixOutputs_andMatrixInput_3_66};
  wire [1:0]   response_data_andMatrixOutputs_hi_66 = {response_data_andMatrixOutputs_andMatrixInput_0_66, response_data_andMatrixOutputs_andMatrixInput_1_66};
  wire         response_data_andMatrixOutputs_1_2_13 = &{response_data_andMatrixOutputs_hi_66, response_data_andMatrixOutputs_lo_66};
  wire [1:0]   response_data_andMatrixOutputs_lo_67 = {response_data_andMatrixOutputs_andMatrixInput_2_67, response_data_andMatrixOutputs_andMatrixInput_3_67};
  wire [1:0]   response_data_andMatrixOutputs_hi_67 = {response_data_andMatrixOutputs_andMatrixInput_0_67, response_data_andMatrixOutputs_andMatrixInput_1_67};
  wire         response_data_andMatrixOutputs_3_2_13 = &{response_data_andMatrixOutputs_hi_67, response_data_andMatrixOutputs_lo_67};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_68 = response_data_invInputs_13[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_68 = response_data_invInputs_13[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_69 = response_data_invInputs_13[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_68 = response_data_plaInput_13[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_69 = response_data_plaInput_13[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_68 = {response_data_andMatrixOutputs_andMatrixInput_3_68, response_data_andMatrixOutputs_andMatrixInput_4_26};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_26 = {response_data_andMatrixOutputs_andMatrixInput_0_68, response_data_andMatrixOutputs_andMatrixInput_1_68};
  wire [2:0]   response_data_andMatrixOutputs_hi_68 = {response_data_andMatrixOutputs_hi_hi_26, response_data_andMatrixOutputs_andMatrixInput_2_68};
  wire         response_data_andMatrixOutputs_0_2_13 = &{response_data_andMatrixOutputs_hi_68, response_data_andMatrixOutputs_lo_68};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_69 = response_data_invInputs_13[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_69 = {response_data_andMatrixOutputs_andMatrixInput_3_69, response_data_andMatrixOutputs_andMatrixInput_4_27};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_27 = {response_data_andMatrixOutputs_andMatrixInput_0_69, response_data_andMatrixOutputs_andMatrixInput_1_69};
  wire [2:0]   response_data_andMatrixOutputs_hi_69 = {response_data_andMatrixOutputs_hi_hi_27, response_data_andMatrixOutputs_andMatrixInput_2_69};
  wire         response_data_andMatrixOutputs_2_2_13 = &{response_data_andMatrixOutputs_hi_69, response_data_andMatrixOutputs_lo_69};
  wire [1:0]   response_data_orMatrixOutputs_lo_13 = {response_data_andMatrixOutputs_0_2_13, response_data_andMatrixOutputs_2_2_13};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_13 = {response_data_andMatrixOutputs_4_2_13, response_data_andMatrixOutputs_1_2_13};
  wire [2:0]   response_data_orMatrixOutputs_hi_13 = {response_data_orMatrixOutputs_hi_hi_13, response_data_andMatrixOutputs_3_2_13};
  wire         response_data_orMatrixOutputs_13 = |{response_data_orMatrixOutputs_hi_13, response_data_orMatrixOutputs_lo_13};
  assign response_data_invMatrixOutputs_13 = response_data_orMatrixOutputs_13;
  wire         response_data_plaOutput_13 = response_data_invMatrixOutputs_13;
  assign response_data_plaInput_13 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[13], request_src_1[13]};
  wire [4:0]   response_data_plaInput_14;
  wire [4:0]   response_data_invInputs_14 = ~response_data_plaInput_14;
  wire         response_data_invMatrixOutputs_14;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_70 = response_data_plaInput_14[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_71 = response_data_plaInput_14[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_73 = response_data_plaInput_14[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_70 = response_data_plaInput_14[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_72 = response_data_plaInput_14[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_74 = response_data_plaInput_14[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_70 = response_data_invInputs_14[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_71 = response_data_invInputs_14[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_72 = response_data_invInputs_14[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_70 = response_data_invInputs_14[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_71 = response_data_invInputs_14[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_72 = response_data_invInputs_14[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_28 = response_data_invInputs_14[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_29 = response_data_invInputs_14[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_70 = {response_data_andMatrixOutputs_andMatrixInput_2_70, response_data_andMatrixOutputs_andMatrixInput_3_70};
  wire [1:0]   response_data_andMatrixOutputs_hi_70 = {response_data_andMatrixOutputs_andMatrixInput_0_70, response_data_andMatrixOutputs_andMatrixInput_1_70};
  wire         response_data_andMatrixOutputs_4_2_14 = &{response_data_andMatrixOutputs_hi_70, response_data_andMatrixOutputs_lo_70};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_71 = response_data_plaInput_14[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_72 = response_data_plaInput_14[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_71 = {response_data_andMatrixOutputs_andMatrixInput_2_71, response_data_andMatrixOutputs_andMatrixInput_3_71};
  wire [1:0]   response_data_andMatrixOutputs_hi_71 = {response_data_andMatrixOutputs_andMatrixInput_0_71, response_data_andMatrixOutputs_andMatrixInput_1_71};
  wire         response_data_andMatrixOutputs_1_2_14 = &{response_data_andMatrixOutputs_hi_71, response_data_andMatrixOutputs_lo_71};
  wire [1:0]   response_data_andMatrixOutputs_lo_72 = {response_data_andMatrixOutputs_andMatrixInput_2_72, response_data_andMatrixOutputs_andMatrixInput_3_72};
  wire [1:0]   response_data_andMatrixOutputs_hi_72 = {response_data_andMatrixOutputs_andMatrixInput_0_72, response_data_andMatrixOutputs_andMatrixInput_1_72};
  wire         response_data_andMatrixOutputs_3_2_14 = &{response_data_andMatrixOutputs_hi_72, response_data_andMatrixOutputs_lo_72};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_73 = response_data_invInputs_14[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_73 = response_data_invInputs_14[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_74 = response_data_invInputs_14[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_73 = response_data_plaInput_14[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_74 = response_data_plaInput_14[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_73 = {response_data_andMatrixOutputs_andMatrixInput_3_73, response_data_andMatrixOutputs_andMatrixInput_4_28};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_28 = {response_data_andMatrixOutputs_andMatrixInput_0_73, response_data_andMatrixOutputs_andMatrixInput_1_73};
  wire [2:0]   response_data_andMatrixOutputs_hi_73 = {response_data_andMatrixOutputs_hi_hi_28, response_data_andMatrixOutputs_andMatrixInput_2_73};
  wire         response_data_andMatrixOutputs_0_2_14 = &{response_data_andMatrixOutputs_hi_73, response_data_andMatrixOutputs_lo_73};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_74 = response_data_invInputs_14[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_74 = {response_data_andMatrixOutputs_andMatrixInput_3_74, response_data_andMatrixOutputs_andMatrixInput_4_29};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_29 = {response_data_andMatrixOutputs_andMatrixInput_0_74, response_data_andMatrixOutputs_andMatrixInput_1_74};
  wire [2:0]   response_data_andMatrixOutputs_hi_74 = {response_data_andMatrixOutputs_hi_hi_29, response_data_andMatrixOutputs_andMatrixInput_2_74};
  wire         response_data_andMatrixOutputs_2_2_14 = &{response_data_andMatrixOutputs_hi_74, response_data_andMatrixOutputs_lo_74};
  wire [1:0]   response_data_orMatrixOutputs_lo_14 = {response_data_andMatrixOutputs_0_2_14, response_data_andMatrixOutputs_2_2_14};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_14 = {response_data_andMatrixOutputs_4_2_14, response_data_andMatrixOutputs_1_2_14};
  wire [2:0]   response_data_orMatrixOutputs_hi_14 = {response_data_orMatrixOutputs_hi_hi_14, response_data_andMatrixOutputs_3_2_14};
  wire         response_data_orMatrixOutputs_14 = |{response_data_orMatrixOutputs_hi_14, response_data_orMatrixOutputs_lo_14};
  assign response_data_invMatrixOutputs_14 = response_data_orMatrixOutputs_14;
  wire         response_data_plaOutput_14 = response_data_invMatrixOutputs_14;
  assign response_data_plaInput_14 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[14], request_src_1[14]};
  wire [4:0]   response_data_plaInput_15;
  wire [4:0]   response_data_invInputs_15 = ~response_data_plaInput_15;
  wire         response_data_invMatrixOutputs_15;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_75 = response_data_plaInput_15[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_76 = response_data_plaInput_15[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_78 = response_data_plaInput_15[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_75 = response_data_plaInput_15[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_77 = response_data_plaInput_15[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_79 = response_data_plaInput_15[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_75 = response_data_invInputs_15[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_76 = response_data_invInputs_15[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_77 = response_data_invInputs_15[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_75 = response_data_invInputs_15[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_76 = response_data_invInputs_15[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_77 = response_data_invInputs_15[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_30 = response_data_invInputs_15[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_31 = response_data_invInputs_15[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_75 = {response_data_andMatrixOutputs_andMatrixInput_2_75, response_data_andMatrixOutputs_andMatrixInput_3_75};
  wire [1:0]   response_data_andMatrixOutputs_hi_75 = {response_data_andMatrixOutputs_andMatrixInput_0_75, response_data_andMatrixOutputs_andMatrixInput_1_75};
  wire         response_data_andMatrixOutputs_4_2_15 = &{response_data_andMatrixOutputs_hi_75, response_data_andMatrixOutputs_lo_75};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_76 = response_data_plaInput_15[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_77 = response_data_plaInput_15[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_76 = {response_data_andMatrixOutputs_andMatrixInput_2_76, response_data_andMatrixOutputs_andMatrixInput_3_76};
  wire [1:0]   response_data_andMatrixOutputs_hi_76 = {response_data_andMatrixOutputs_andMatrixInput_0_76, response_data_andMatrixOutputs_andMatrixInput_1_76};
  wire         response_data_andMatrixOutputs_1_2_15 = &{response_data_andMatrixOutputs_hi_76, response_data_andMatrixOutputs_lo_76};
  wire [1:0]   response_data_andMatrixOutputs_lo_77 = {response_data_andMatrixOutputs_andMatrixInput_2_77, response_data_andMatrixOutputs_andMatrixInput_3_77};
  wire [1:0]   response_data_andMatrixOutputs_hi_77 = {response_data_andMatrixOutputs_andMatrixInput_0_77, response_data_andMatrixOutputs_andMatrixInput_1_77};
  wire         response_data_andMatrixOutputs_3_2_15 = &{response_data_andMatrixOutputs_hi_77, response_data_andMatrixOutputs_lo_77};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_78 = response_data_invInputs_15[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_78 = response_data_invInputs_15[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_79 = response_data_invInputs_15[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_78 = response_data_plaInput_15[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_79 = response_data_plaInput_15[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_78 = {response_data_andMatrixOutputs_andMatrixInput_3_78, response_data_andMatrixOutputs_andMatrixInput_4_30};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_30 = {response_data_andMatrixOutputs_andMatrixInput_0_78, response_data_andMatrixOutputs_andMatrixInput_1_78};
  wire [2:0]   response_data_andMatrixOutputs_hi_78 = {response_data_andMatrixOutputs_hi_hi_30, response_data_andMatrixOutputs_andMatrixInput_2_78};
  wire         response_data_andMatrixOutputs_0_2_15 = &{response_data_andMatrixOutputs_hi_78, response_data_andMatrixOutputs_lo_78};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_79 = response_data_invInputs_15[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_79 = {response_data_andMatrixOutputs_andMatrixInput_3_79, response_data_andMatrixOutputs_andMatrixInput_4_31};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_31 = {response_data_andMatrixOutputs_andMatrixInput_0_79, response_data_andMatrixOutputs_andMatrixInput_1_79};
  wire [2:0]   response_data_andMatrixOutputs_hi_79 = {response_data_andMatrixOutputs_hi_hi_31, response_data_andMatrixOutputs_andMatrixInput_2_79};
  wire         response_data_andMatrixOutputs_2_2_15 = &{response_data_andMatrixOutputs_hi_79, response_data_andMatrixOutputs_lo_79};
  wire [1:0]   response_data_orMatrixOutputs_lo_15 = {response_data_andMatrixOutputs_0_2_15, response_data_andMatrixOutputs_2_2_15};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_15 = {response_data_andMatrixOutputs_4_2_15, response_data_andMatrixOutputs_1_2_15};
  wire [2:0]   response_data_orMatrixOutputs_hi_15 = {response_data_orMatrixOutputs_hi_hi_15, response_data_andMatrixOutputs_3_2_15};
  wire         response_data_orMatrixOutputs_15 = |{response_data_orMatrixOutputs_hi_15, response_data_orMatrixOutputs_lo_15};
  assign response_data_invMatrixOutputs_15 = response_data_orMatrixOutputs_15;
  wire         response_data_plaOutput_15 = response_data_invMatrixOutputs_15;
  assign response_data_plaInput_15 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[15], request_src_1[15]};
  wire [4:0]   response_data_plaInput_16;
  wire [4:0]   response_data_invInputs_16 = ~response_data_plaInput_16;
  wire         response_data_invMatrixOutputs_16;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_80 = response_data_plaInput_16[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_81 = response_data_plaInput_16[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_83 = response_data_plaInput_16[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_80 = response_data_plaInput_16[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_82 = response_data_plaInput_16[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_84 = response_data_plaInput_16[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_80 = response_data_invInputs_16[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_81 = response_data_invInputs_16[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_82 = response_data_invInputs_16[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_80 = response_data_invInputs_16[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_81 = response_data_invInputs_16[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_82 = response_data_invInputs_16[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_32 = response_data_invInputs_16[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_33 = response_data_invInputs_16[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_80 = {response_data_andMatrixOutputs_andMatrixInput_2_80, response_data_andMatrixOutputs_andMatrixInput_3_80};
  wire [1:0]   response_data_andMatrixOutputs_hi_80 = {response_data_andMatrixOutputs_andMatrixInput_0_80, response_data_andMatrixOutputs_andMatrixInput_1_80};
  wire         response_data_andMatrixOutputs_4_2_16 = &{response_data_andMatrixOutputs_hi_80, response_data_andMatrixOutputs_lo_80};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_81 = response_data_plaInput_16[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_82 = response_data_plaInput_16[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_81 = {response_data_andMatrixOutputs_andMatrixInput_2_81, response_data_andMatrixOutputs_andMatrixInput_3_81};
  wire [1:0]   response_data_andMatrixOutputs_hi_81 = {response_data_andMatrixOutputs_andMatrixInput_0_81, response_data_andMatrixOutputs_andMatrixInput_1_81};
  wire         response_data_andMatrixOutputs_1_2_16 = &{response_data_andMatrixOutputs_hi_81, response_data_andMatrixOutputs_lo_81};
  wire [1:0]   response_data_andMatrixOutputs_lo_82 = {response_data_andMatrixOutputs_andMatrixInput_2_82, response_data_andMatrixOutputs_andMatrixInput_3_82};
  wire [1:0]   response_data_andMatrixOutputs_hi_82 = {response_data_andMatrixOutputs_andMatrixInput_0_82, response_data_andMatrixOutputs_andMatrixInput_1_82};
  wire         response_data_andMatrixOutputs_3_2_16 = &{response_data_andMatrixOutputs_hi_82, response_data_andMatrixOutputs_lo_82};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_83 = response_data_invInputs_16[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_83 = response_data_invInputs_16[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_84 = response_data_invInputs_16[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_83 = response_data_plaInput_16[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_84 = response_data_plaInput_16[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_83 = {response_data_andMatrixOutputs_andMatrixInput_3_83, response_data_andMatrixOutputs_andMatrixInput_4_32};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_32 = {response_data_andMatrixOutputs_andMatrixInput_0_83, response_data_andMatrixOutputs_andMatrixInput_1_83};
  wire [2:0]   response_data_andMatrixOutputs_hi_83 = {response_data_andMatrixOutputs_hi_hi_32, response_data_andMatrixOutputs_andMatrixInput_2_83};
  wire         response_data_andMatrixOutputs_0_2_16 = &{response_data_andMatrixOutputs_hi_83, response_data_andMatrixOutputs_lo_83};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_84 = response_data_invInputs_16[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_84 = {response_data_andMatrixOutputs_andMatrixInput_3_84, response_data_andMatrixOutputs_andMatrixInput_4_33};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_33 = {response_data_andMatrixOutputs_andMatrixInput_0_84, response_data_andMatrixOutputs_andMatrixInput_1_84};
  wire [2:0]   response_data_andMatrixOutputs_hi_84 = {response_data_andMatrixOutputs_hi_hi_33, response_data_andMatrixOutputs_andMatrixInput_2_84};
  wire         response_data_andMatrixOutputs_2_2_16 = &{response_data_andMatrixOutputs_hi_84, response_data_andMatrixOutputs_lo_84};
  wire [1:0]   response_data_orMatrixOutputs_lo_16 = {response_data_andMatrixOutputs_0_2_16, response_data_andMatrixOutputs_2_2_16};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_16 = {response_data_andMatrixOutputs_4_2_16, response_data_andMatrixOutputs_1_2_16};
  wire [2:0]   response_data_orMatrixOutputs_hi_16 = {response_data_orMatrixOutputs_hi_hi_16, response_data_andMatrixOutputs_3_2_16};
  wire         response_data_orMatrixOutputs_16 = |{response_data_orMatrixOutputs_hi_16, response_data_orMatrixOutputs_lo_16};
  assign response_data_invMatrixOutputs_16 = response_data_orMatrixOutputs_16;
  wire         response_data_plaOutput_16 = response_data_invMatrixOutputs_16;
  assign response_data_plaInput_16 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[16], request_src_1[16]};
  wire [4:0]   response_data_plaInput_17;
  wire [4:0]   response_data_invInputs_17 = ~response_data_plaInput_17;
  wire         response_data_invMatrixOutputs_17;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_85 = response_data_plaInput_17[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_86 = response_data_plaInput_17[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_88 = response_data_plaInput_17[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_85 = response_data_plaInput_17[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_87 = response_data_plaInput_17[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_89 = response_data_plaInput_17[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_85 = response_data_invInputs_17[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_86 = response_data_invInputs_17[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_87 = response_data_invInputs_17[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_85 = response_data_invInputs_17[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_86 = response_data_invInputs_17[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_87 = response_data_invInputs_17[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_34 = response_data_invInputs_17[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_35 = response_data_invInputs_17[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_85 = {response_data_andMatrixOutputs_andMatrixInput_2_85, response_data_andMatrixOutputs_andMatrixInput_3_85};
  wire [1:0]   response_data_andMatrixOutputs_hi_85 = {response_data_andMatrixOutputs_andMatrixInput_0_85, response_data_andMatrixOutputs_andMatrixInput_1_85};
  wire         response_data_andMatrixOutputs_4_2_17 = &{response_data_andMatrixOutputs_hi_85, response_data_andMatrixOutputs_lo_85};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_86 = response_data_plaInput_17[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_87 = response_data_plaInput_17[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_86 = {response_data_andMatrixOutputs_andMatrixInput_2_86, response_data_andMatrixOutputs_andMatrixInput_3_86};
  wire [1:0]   response_data_andMatrixOutputs_hi_86 = {response_data_andMatrixOutputs_andMatrixInput_0_86, response_data_andMatrixOutputs_andMatrixInput_1_86};
  wire         response_data_andMatrixOutputs_1_2_17 = &{response_data_andMatrixOutputs_hi_86, response_data_andMatrixOutputs_lo_86};
  wire [1:0]   response_data_andMatrixOutputs_lo_87 = {response_data_andMatrixOutputs_andMatrixInput_2_87, response_data_andMatrixOutputs_andMatrixInput_3_87};
  wire [1:0]   response_data_andMatrixOutputs_hi_87 = {response_data_andMatrixOutputs_andMatrixInput_0_87, response_data_andMatrixOutputs_andMatrixInput_1_87};
  wire         response_data_andMatrixOutputs_3_2_17 = &{response_data_andMatrixOutputs_hi_87, response_data_andMatrixOutputs_lo_87};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_88 = response_data_invInputs_17[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_88 = response_data_invInputs_17[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_89 = response_data_invInputs_17[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_88 = response_data_plaInput_17[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_89 = response_data_plaInput_17[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_88 = {response_data_andMatrixOutputs_andMatrixInput_3_88, response_data_andMatrixOutputs_andMatrixInput_4_34};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_34 = {response_data_andMatrixOutputs_andMatrixInput_0_88, response_data_andMatrixOutputs_andMatrixInput_1_88};
  wire [2:0]   response_data_andMatrixOutputs_hi_88 = {response_data_andMatrixOutputs_hi_hi_34, response_data_andMatrixOutputs_andMatrixInput_2_88};
  wire         response_data_andMatrixOutputs_0_2_17 = &{response_data_andMatrixOutputs_hi_88, response_data_andMatrixOutputs_lo_88};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_89 = response_data_invInputs_17[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_89 = {response_data_andMatrixOutputs_andMatrixInput_3_89, response_data_andMatrixOutputs_andMatrixInput_4_35};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_35 = {response_data_andMatrixOutputs_andMatrixInput_0_89, response_data_andMatrixOutputs_andMatrixInput_1_89};
  wire [2:0]   response_data_andMatrixOutputs_hi_89 = {response_data_andMatrixOutputs_hi_hi_35, response_data_andMatrixOutputs_andMatrixInput_2_89};
  wire         response_data_andMatrixOutputs_2_2_17 = &{response_data_andMatrixOutputs_hi_89, response_data_andMatrixOutputs_lo_89};
  wire [1:0]   response_data_orMatrixOutputs_lo_17 = {response_data_andMatrixOutputs_0_2_17, response_data_andMatrixOutputs_2_2_17};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_17 = {response_data_andMatrixOutputs_4_2_17, response_data_andMatrixOutputs_1_2_17};
  wire [2:0]   response_data_orMatrixOutputs_hi_17 = {response_data_orMatrixOutputs_hi_hi_17, response_data_andMatrixOutputs_3_2_17};
  wire         response_data_orMatrixOutputs_17 = |{response_data_orMatrixOutputs_hi_17, response_data_orMatrixOutputs_lo_17};
  assign response_data_invMatrixOutputs_17 = response_data_orMatrixOutputs_17;
  wire         response_data_plaOutput_17 = response_data_invMatrixOutputs_17;
  assign response_data_plaInput_17 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[17], request_src_1[17]};
  wire [4:0]   response_data_plaInput_18;
  wire [4:0]   response_data_invInputs_18 = ~response_data_plaInput_18;
  wire         response_data_invMatrixOutputs_18;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_90 = response_data_plaInput_18[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_91 = response_data_plaInput_18[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_93 = response_data_plaInput_18[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_90 = response_data_plaInput_18[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_92 = response_data_plaInput_18[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_94 = response_data_plaInput_18[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_90 = response_data_invInputs_18[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_91 = response_data_invInputs_18[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_92 = response_data_invInputs_18[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_90 = response_data_invInputs_18[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_91 = response_data_invInputs_18[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_92 = response_data_invInputs_18[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_36 = response_data_invInputs_18[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_37 = response_data_invInputs_18[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_90 = {response_data_andMatrixOutputs_andMatrixInput_2_90, response_data_andMatrixOutputs_andMatrixInput_3_90};
  wire [1:0]   response_data_andMatrixOutputs_hi_90 = {response_data_andMatrixOutputs_andMatrixInput_0_90, response_data_andMatrixOutputs_andMatrixInput_1_90};
  wire         response_data_andMatrixOutputs_4_2_18 = &{response_data_andMatrixOutputs_hi_90, response_data_andMatrixOutputs_lo_90};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_91 = response_data_plaInput_18[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_92 = response_data_plaInput_18[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_91 = {response_data_andMatrixOutputs_andMatrixInput_2_91, response_data_andMatrixOutputs_andMatrixInput_3_91};
  wire [1:0]   response_data_andMatrixOutputs_hi_91 = {response_data_andMatrixOutputs_andMatrixInput_0_91, response_data_andMatrixOutputs_andMatrixInput_1_91};
  wire         response_data_andMatrixOutputs_1_2_18 = &{response_data_andMatrixOutputs_hi_91, response_data_andMatrixOutputs_lo_91};
  wire [1:0]   response_data_andMatrixOutputs_lo_92 = {response_data_andMatrixOutputs_andMatrixInput_2_92, response_data_andMatrixOutputs_andMatrixInput_3_92};
  wire [1:0]   response_data_andMatrixOutputs_hi_92 = {response_data_andMatrixOutputs_andMatrixInput_0_92, response_data_andMatrixOutputs_andMatrixInput_1_92};
  wire         response_data_andMatrixOutputs_3_2_18 = &{response_data_andMatrixOutputs_hi_92, response_data_andMatrixOutputs_lo_92};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_93 = response_data_invInputs_18[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_93 = response_data_invInputs_18[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_94 = response_data_invInputs_18[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_93 = response_data_plaInput_18[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_94 = response_data_plaInput_18[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_93 = {response_data_andMatrixOutputs_andMatrixInput_3_93, response_data_andMatrixOutputs_andMatrixInput_4_36};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_36 = {response_data_andMatrixOutputs_andMatrixInput_0_93, response_data_andMatrixOutputs_andMatrixInput_1_93};
  wire [2:0]   response_data_andMatrixOutputs_hi_93 = {response_data_andMatrixOutputs_hi_hi_36, response_data_andMatrixOutputs_andMatrixInput_2_93};
  wire         response_data_andMatrixOutputs_0_2_18 = &{response_data_andMatrixOutputs_hi_93, response_data_andMatrixOutputs_lo_93};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_94 = response_data_invInputs_18[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_94 = {response_data_andMatrixOutputs_andMatrixInput_3_94, response_data_andMatrixOutputs_andMatrixInput_4_37};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_37 = {response_data_andMatrixOutputs_andMatrixInput_0_94, response_data_andMatrixOutputs_andMatrixInput_1_94};
  wire [2:0]   response_data_andMatrixOutputs_hi_94 = {response_data_andMatrixOutputs_hi_hi_37, response_data_andMatrixOutputs_andMatrixInput_2_94};
  wire         response_data_andMatrixOutputs_2_2_18 = &{response_data_andMatrixOutputs_hi_94, response_data_andMatrixOutputs_lo_94};
  wire [1:0]   response_data_orMatrixOutputs_lo_18 = {response_data_andMatrixOutputs_0_2_18, response_data_andMatrixOutputs_2_2_18};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_18 = {response_data_andMatrixOutputs_4_2_18, response_data_andMatrixOutputs_1_2_18};
  wire [2:0]   response_data_orMatrixOutputs_hi_18 = {response_data_orMatrixOutputs_hi_hi_18, response_data_andMatrixOutputs_3_2_18};
  wire         response_data_orMatrixOutputs_18 = |{response_data_orMatrixOutputs_hi_18, response_data_orMatrixOutputs_lo_18};
  assign response_data_invMatrixOutputs_18 = response_data_orMatrixOutputs_18;
  wire         response_data_plaOutput_18 = response_data_invMatrixOutputs_18;
  assign response_data_plaInput_18 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[18], request_src_1[18]};
  wire [4:0]   response_data_plaInput_19;
  wire [4:0]   response_data_invInputs_19 = ~response_data_plaInput_19;
  wire         response_data_invMatrixOutputs_19;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_95 = response_data_plaInput_19[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_96 = response_data_plaInput_19[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_98 = response_data_plaInput_19[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_95 = response_data_plaInput_19[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_97 = response_data_plaInput_19[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_99 = response_data_plaInput_19[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_95 = response_data_invInputs_19[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_96 = response_data_invInputs_19[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_97 = response_data_invInputs_19[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_95 = response_data_invInputs_19[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_96 = response_data_invInputs_19[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_97 = response_data_invInputs_19[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_38 = response_data_invInputs_19[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_39 = response_data_invInputs_19[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_95 = {response_data_andMatrixOutputs_andMatrixInput_2_95, response_data_andMatrixOutputs_andMatrixInput_3_95};
  wire [1:0]   response_data_andMatrixOutputs_hi_95 = {response_data_andMatrixOutputs_andMatrixInput_0_95, response_data_andMatrixOutputs_andMatrixInput_1_95};
  wire         response_data_andMatrixOutputs_4_2_19 = &{response_data_andMatrixOutputs_hi_95, response_data_andMatrixOutputs_lo_95};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_96 = response_data_plaInput_19[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_97 = response_data_plaInput_19[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_96 = {response_data_andMatrixOutputs_andMatrixInput_2_96, response_data_andMatrixOutputs_andMatrixInput_3_96};
  wire [1:0]   response_data_andMatrixOutputs_hi_96 = {response_data_andMatrixOutputs_andMatrixInput_0_96, response_data_andMatrixOutputs_andMatrixInput_1_96};
  wire         response_data_andMatrixOutputs_1_2_19 = &{response_data_andMatrixOutputs_hi_96, response_data_andMatrixOutputs_lo_96};
  wire [1:0]   response_data_andMatrixOutputs_lo_97 = {response_data_andMatrixOutputs_andMatrixInput_2_97, response_data_andMatrixOutputs_andMatrixInput_3_97};
  wire [1:0]   response_data_andMatrixOutputs_hi_97 = {response_data_andMatrixOutputs_andMatrixInput_0_97, response_data_andMatrixOutputs_andMatrixInput_1_97};
  wire         response_data_andMatrixOutputs_3_2_19 = &{response_data_andMatrixOutputs_hi_97, response_data_andMatrixOutputs_lo_97};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_98 = response_data_invInputs_19[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_98 = response_data_invInputs_19[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_99 = response_data_invInputs_19[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_98 = response_data_plaInput_19[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_99 = response_data_plaInput_19[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_98 = {response_data_andMatrixOutputs_andMatrixInput_3_98, response_data_andMatrixOutputs_andMatrixInput_4_38};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_38 = {response_data_andMatrixOutputs_andMatrixInput_0_98, response_data_andMatrixOutputs_andMatrixInput_1_98};
  wire [2:0]   response_data_andMatrixOutputs_hi_98 = {response_data_andMatrixOutputs_hi_hi_38, response_data_andMatrixOutputs_andMatrixInput_2_98};
  wire         response_data_andMatrixOutputs_0_2_19 = &{response_data_andMatrixOutputs_hi_98, response_data_andMatrixOutputs_lo_98};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_99 = response_data_invInputs_19[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_99 = {response_data_andMatrixOutputs_andMatrixInput_3_99, response_data_andMatrixOutputs_andMatrixInput_4_39};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_39 = {response_data_andMatrixOutputs_andMatrixInput_0_99, response_data_andMatrixOutputs_andMatrixInput_1_99};
  wire [2:0]   response_data_andMatrixOutputs_hi_99 = {response_data_andMatrixOutputs_hi_hi_39, response_data_andMatrixOutputs_andMatrixInput_2_99};
  wire         response_data_andMatrixOutputs_2_2_19 = &{response_data_andMatrixOutputs_hi_99, response_data_andMatrixOutputs_lo_99};
  wire [1:0]   response_data_orMatrixOutputs_lo_19 = {response_data_andMatrixOutputs_0_2_19, response_data_andMatrixOutputs_2_2_19};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_19 = {response_data_andMatrixOutputs_4_2_19, response_data_andMatrixOutputs_1_2_19};
  wire [2:0]   response_data_orMatrixOutputs_hi_19 = {response_data_orMatrixOutputs_hi_hi_19, response_data_andMatrixOutputs_3_2_19};
  wire         response_data_orMatrixOutputs_19 = |{response_data_orMatrixOutputs_hi_19, response_data_orMatrixOutputs_lo_19};
  assign response_data_invMatrixOutputs_19 = response_data_orMatrixOutputs_19;
  wire         response_data_plaOutput_19 = response_data_invMatrixOutputs_19;
  assign response_data_plaInput_19 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[19], request_src_1[19]};
  wire [4:0]   response_data_plaInput_20;
  wire [4:0]   response_data_invInputs_20 = ~response_data_plaInput_20;
  wire         response_data_invMatrixOutputs_20;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_100 = response_data_plaInput_20[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_101 = response_data_plaInput_20[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_103 = response_data_plaInput_20[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_100 = response_data_plaInput_20[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_102 = response_data_plaInput_20[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_104 = response_data_plaInput_20[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_100 = response_data_invInputs_20[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_101 = response_data_invInputs_20[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_102 = response_data_invInputs_20[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_100 = response_data_invInputs_20[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_101 = response_data_invInputs_20[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_102 = response_data_invInputs_20[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_40 = response_data_invInputs_20[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_41 = response_data_invInputs_20[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_100 = {response_data_andMatrixOutputs_andMatrixInput_2_100, response_data_andMatrixOutputs_andMatrixInput_3_100};
  wire [1:0]   response_data_andMatrixOutputs_hi_100 = {response_data_andMatrixOutputs_andMatrixInput_0_100, response_data_andMatrixOutputs_andMatrixInput_1_100};
  wire         response_data_andMatrixOutputs_4_2_20 = &{response_data_andMatrixOutputs_hi_100, response_data_andMatrixOutputs_lo_100};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_101 = response_data_plaInput_20[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_102 = response_data_plaInput_20[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_101 = {response_data_andMatrixOutputs_andMatrixInput_2_101, response_data_andMatrixOutputs_andMatrixInput_3_101};
  wire [1:0]   response_data_andMatrixOutputs_hi_101 = {response_data_andMatrixOutputs_andMatrixInput_0_101, response_data_andMatrixOutputs_andMatrixInput_1_101};
  wire         response_data_andMatrixOutputs_1_2_20 = &{response_data_andMatrixOutputs_hi_101, response_data_andMatrixOutputs_lo_101};
  wire [1:0]   response_data_andMatrixOutputs_lo_102 = {response_data_andMatrixOutputs_andMatrixInput_2_102, response_data_andMatrixOutputs_andMatrixInput_3_102};
  wire [1:0]   response_data_andMatrixOutputs_hi_102 = {response_data_andMatrixOutputs_andMatrixInput_0_102, response_data_andMatrixOutputs_andMatrixInput_1_102};
  wire         response_data_andMatrixOutputs_3_2_20 = &{response_data_andMatrixOutputs_hi_102, response_data_andMatrixOutputs_lo_102};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_103 = response_data_invInputs_20[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_103 = response_data_invInputs_20[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_104 = response_data_invInputs_20[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_103 = response_data_plaInput_20[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_104 = response_data_plaInput_20[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_103 = {response_data_andMatrixOutputs_andMatrixInput_3_103, response_data_andMatrixOutputs_andMatrixInput_4_40};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_40 = {response_data_andMatrixOutputs_andMatrixInput_0_103, response_data_andMatrixOutputs_andMatrixInput_1_103};
  wire [2:0]   response_data_andMatrixOutputs_hi_103 = {response_data_andMatrixOutputs_hi_hi_40, response_data_andMatrixOutputs_andMatrixInput_2_103};
  wire         response_data_andMatrixOutputs_0_2_20 = &{response_data_andMatrixOutputs_hi_103, response_data_andMatrixOutputs_lo_103};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_104 = response_data_invInputs_20[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_104 = {response_data_andMatrixOutputs_andMatrixInput_3_104, response_data_andMatrixOutputs_andMatrixInput_4_41};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_41 = {response_data_andMatrixOutputs_andMatrixInput_0_104, response_data_andMatrixOutputs_andMatrixInput_1_104};
  wire [2:0]   response_data_andMatrixOutputs_hi_104 = {response_data_andMatrixOutputs_hi_hi_41, response_data_andMatrixOutputs_andMatrixInput_2_104};
  wire         response_data_andMatrixOutputs_2_2_20 = &{response_data_andMatrixOutputs_hi_104, response_data_andMatrixOutputs_lo_104};
  wire [1:0]   response_data_orMatrixOutputs_lo_20 = {response_data_andMatrixOutputs_0_2_20, response_data_andMatrixOutputs_2_2_20};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_20 = {response_data_andMatrixOutputs_4_2_20, response_data_andMatrixOutputs_1_2_20};
  wire [2:0]   response_data_orMatrixOutputs_hi_20 = {response_data_orMatrixOutputs_hi_hi_20, response_data_andMatrixOutputs_3_2_20};
  wire         response_data_orMatrixOutputs_20 = |{response_data_orMatrixOutputs_hi_20, response_data_orMatrixOutputs_lo_20};
  assign response_data_invMatrixOutputs_20 = response_data_orMatrixOutputs_20;
  wire         response_data_plaOutput_20 = response_data_invMatrixOutputs_20;
  assign response_data_plaInput_20 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[20], request_src_1[20]};
  wire [4:0]   response_data_plaInput_21;
  wire [4:0]   response_data_invInputs_21 = ~response_data_plaInput_21;
  wire         response_data_invMatrixOutputs_21;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_105 = response_data_plaInput_21[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_106 = response_data_plaInput_21[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_108 = response_data_plaInput_21[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_105 = response_data_plaInput_21[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_107 = response_data_plaInput_21[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_109 = response_data_plaInput_21[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_105 = response_data_invInputs_21[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_106 = response_data_invInputs_21[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_107 = response_data_invInputs_21[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_105 = response_data_invInputs_21[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_106 = response_data_invInputs_21[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_107 = response_data_invInputs_21[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_42 = response_data_invInputs_21[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_43 = response_data_invInputs_21[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_105 = {response_data_andMatrixOutputs_andMatrixInput_2_105, response_data_andMatrixOutputs_andMatrixInput_3_105};
  wire [1:0]   response_data_andMatrixOutputs_hi_105 = {response_data_andMatrixOutputs_andMatrixInput_0_105, response_data_andMatrixOutputs_andMatrixInput_1_105};
  wire         response_data_andMatrixOutputs_4_2_21 = &{response_data_andMatrixOutputs_hi_105, response_data_andMatrixOutputs_lo_105};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_106 = response_data_plaInput_21[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_107 = response_data_plaInput_21[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_106 = {response_data_andMatrixOutputs_andMatrixInput_2_106, response_data_andMatrixOutputs_andMatrixInput_3_106};
  wire [1:0]   response_data_andMatrixOutputs_hi_106 = {response_data_andMatrixOutputs_andMatrixInput_0_106, response_data_andMatrixOutputs_andMatrixInput_1_106};
  wire         response_data_andMatrixOutputs_1_2_21 = &{response_data_andMatrixOutputs_hi_106, response_data_andMatrixOutputs_lo_106};
  wire [1:0]   response_data_andMatrixOutputs_lo_107 = {response_data_andMatrixOutputs_andMatrixInput_2_107, response_data_andMatrixOutputs_andMatrixInput_3_107};
  wire [1:0]   response_data_andMatrixOutputs_hi_107 = {response_data_andMatrixOutputs_andMatrixInput_0_107, response_data_andMatrixOutputs_andMatrixInput_1_107};
  wire         response_data_andMatrixOutputs_3_2_21 = &{response_data_andMatrixOutputs_hi_107, response_data_andMatrixOutputs_lo_107};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_108 = response_data_invInputs_21[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_108 = response_data_invInputs_21[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_109 = response_data_invInputs_21[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_108 = response_data_plaInput_21[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_109 = response_data_plaInput_21[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_108 = {response_data_andMatrixOutputs_andMatrixInput_3_108, response_data_andMatrixOutputs_andMatrixInput_4_42};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_42 = {response_data_andMatrixOutputs_andMatrixInput_0_108, response_data_andMatrixOutputs_andMatrixInput_1_108};
  wire [2:0]   response_data_andMatrixOutputs_hi_108 = {response_data_andMatrixOutputs_hi_hi_42, response_data_andMatrixOutputs_andMatrixInput_2_108};
  wire         response_data_andMatrixOutputs_0_2_21 = &{response_data_andMatrixOutputs_hi_108, response_data_andMatrixOutputs_lo_108};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_109 = response_data_invInputs_21[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_109 = {response_data_andMatrixOutputs_andMatrixInput_3_109, response_data_andMatrixOutputs_andMatrixInput_4_43};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_43 = {response_data_andMatrixOutputs_andMatrixInput_0_109, response_data_andMatrixOutputs_andMatrixInput_1_109};
  wire [2:0]   response_data_andMatrixOutputs_hi_109 = {response_data_andMatrixOutputs_hi_hi_43, response_data_andMatrixOutputs_andMatrixInput_2_109};
  wire         response_data_andMatrixOutputs_2_2_21 = &{response_data_andMatrixOutputs_hi_109, response_data_andMatrixOutputs_lo_109};
  wire [1:0]   response_data_orMatrixOutputs_lo_21 = {response_data_andMatrixOutputs_0_2_21, response_data_andMatrixOutputs_2_2_21};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_21 = {response_data_andMatrixOutputs_4_2_21, response_data_andMatrixOutputs_1_2_21};
  wire [2:0]   response_data_orMatrixOutputs_hi_21 = {response_data_orMatrixOutputs_hi_hi_21, response_data_andMatrixOutputs_3_2_21};
  wire         response_data_orMatrixOutputs_21 = |{response_data_orMatrixOutputs_hi_21, response_data_orMatrixOutputs_lo_21};
  assign response_data_invMatrixOutputs_21 = response_data_orMatrixOutputs_21;
  wire         response_data_plaOutput_21 = response_data_invMatrixOutputs_21;
  assign response_data_plaInput_21 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[21], request_src_1[21]};
  wire [4:0]   response_data_plaInput_22;
  wire [4:0]   response_data_invInputs_22 = ~response_data_plaInput_22;
  wire         response_data_invMatrixOutputs_22;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_110 = response_data_plaInput_22[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_111 = response_data_plaInput_22[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_113 = response_data_plaInput_22[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_110 = response_data_plaInput_22[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_112 = response_data_plaInput_22[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_114 = response_data_plaInput_22[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_110 = response_data_invInputs_22[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_111 = response_data_invInputs_22[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_112 = response_data_invInputs_22[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_110 = response_data_invInputs_22[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_111 = response_data_invInputs_22[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_112 = response_data_invInputs_22[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_44 = response_data_invInputs_22[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_45 = response_data_invInputs_22[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_110 = {response_data_andMatrixOutputs_andMatrixInput_2_110, response_data_andMatrixOutputs_andMatrixInput_3_110};
  wire [1:0]   response_data_andMatrixOutputs_hi_110 = {response_data_andMatrixOutputs_andMatrixInput_0_110, response_data_andMatrixOutputs_andMatrixInput_1_110};
  wire         response_data_andMatrixOutputs_4_2_22 = &{response_data_andMatrixOutputs_hi_110, response_data_andMatrixOutputs_lo_110};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_111 = response_data_plaInput_22[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_112 = response_data_plaInput_22[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_111 = {response_data_andMatrixOutputs_andMatrixInput_2_111, response_data_andMatrixOutputs_andMatrixInput_3_111};
  wire [1:0]   response_data_andMatrixOutputs_hi_111 = {response_data_andMatrixOutputs_andMatrixInput_0_111, response_data_andMatrixOutputs_andMatrixInput_1_111};
  wire         response_data_andMatrixOutputs_1_2_22 = &{response_data_andMatrixOutputs_hi_111, response_data_andMatrixOutputs_lo_111};
  wire [1:0]   response_data_andMatrixOutputs_lo_112 = {response_data_andMatrixOutputs_andMatrixInput_2_112, response_data_andMatrixOutputs_andMatrixInput_3_112};
  wire [1:0]   response_data_andMatrixOutputs_hi_112 = {response_data_andMatrixOutputs_andMatrixInput_0_112, response_data_andMatrixOutputs_andMatrixInput_1_112};
  wire         response_data_andMatrixOutputs_3_2_22 = &{response_data_andMatrixOutputs_hi_112, response_data_andMatrixOutputs_lo_112};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_113 = response_data_invInputs_22[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_113 = response_data_invInputs_22[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_114 = response_data_invInputs_22[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_113 = response_data_plaInput_22[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_114 = response_data_plaInput_22[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_113 = {response_data_andMatrixOutputs_andMatrixInput_3_113, response_data_andMatrixOutputs_andMatrixInput_4_44};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_44 = {response_data_andMatrixOutputs_andMatrixInput_0_113, response_data_andMatrixOutputs_andMatrixInput_1_113};
  wire [2:0]   response_data_andMatrixOutputs_hi_113 = {response_data_andMatrixOutputs_hi_hi_44, response_data_andMatrixOutputs_andMatrixInput_2_113};
  wire         response_data_andMatrixOutputs_0_2_22 = &{response_data_andMatrixOutputs_hi_113, response_data_andMatrixOutputs_lo_113};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_114 = response_data_invInputs_22[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_114 = {response_data_andMatrixOutputs_andMatrixInput_3_114, response_data_andMatrixOutputs_andMatrixInput_4_45};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_45 = {response_data_andMatrixOutputs_andMatrixInput_0_114, response_data_andMatrixOutputs_andMatrixInput_1_114};
  wire [2:0]   response_data_andMatrixOutputs_hi_114 = {response_data_andMatrixOutputs_hi_hi_45, response_data_andMatrixOutputs_andMatrixInput_2_114};
  wire         response_data_andMatrixOutputs_2_2_22 = &{response_data_andMatrixOutputs_hi_114, response_data_andMatrixOutputs_lo_114};
  wire [1:0]   response_data_orMatrixOutputs_lo_22 = {response_data_andMatrixOutputs_0_2_22, response_data_andMatrixOutputs_2_2_22};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_22 = {response_data_andMatrixOutputs_4_2_22, response_data_andMatrixOutputs_1_2_22};
  wire [2:0]   response_data_orMatrixOutputs_hi_22 = {response_data_orMatrixOutputs_hi_hi_22, response_data_andMatrixOutputs_3_2_22};
  wire         response_data_orMatrixOutputs_22 = |{response_data_orMatrixOutputs_hi_22, response_data_orMatrixOutputs_lo_22};
  assign response_data_invMatrixOutputs_22 = response_data_orMatrixOutputs_22;
  wire         response_data_plaOutput_22 = response_data_invMatrixOutputs_22;
  assign response_data_plaInput_22 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[22], request_src_1[22]};
  wire [4:0]   response_data_plaInput_23;
  wire [4:0]   response_data_invInputs_23 = ~response_data_plaInput_23;
  wire         response_data_invMatrixOutputs_23;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_115 = response_data_plaInput_23[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_116 = response_data_plaInput_23[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_118 = response_data_plaInput_23[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_115 = response_data_plaInput_23[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_117 = response_data_plaInput_23[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_119 = response_data_plaInput_23[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_115 = response_data_invInputs_23[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_116 = response_data_invInputs_23[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_117 = response_data_invInputs_23[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_115 = response_data_invInputs_23[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_116 = response_data_invInputs_23[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_117 = response_data_invInputs_23[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_46 = response_data_invInputs_23[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_47 = response_data_invInputs_23[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_115 = {response_data_andMatrixOutputs_andMatrixInput_2_115, response_data_andMatrixOutputs_andMatrixInput_3_115};
  wire [1:0]   response_data_andMatrixOutputs_hi_115 = {response_data_andMatrixOutputs_andMatrixInput_0_115, response_data_andMatrixOutputs_andMatrixInput_1_115};
  wire         response_data_andMatrixOutputs_4_2_23 = &{response_data_andMatrixOutputs_hi_115, response_data_andMatrixOutputs_lo_115};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_116 = response_data_plaInput_23[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_117 = response_data_plaInput_23[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_116 = {response_data_andMatrixOutputs_andMatrixInput_2_116, response_data_andMatrixOutputs_andMatrixInput_3_116};
  wire [1:0]   response_data_andMatrixOutputs_hi_116 = {response_data_andMatrixOutputs_andMatrixInput_0_116, response_data_andMatrixOutputs_andMatrixInput_1_116};
  wire         response_data_andMatrixOutputs_1_2_23 = &{response_data_andMatrixOutputs_hi_116, response_data_andMatrixOutputs_lo_116};
  wire [1:0]   response_data_andMatrixOutputs_lo_117 = {response_data_andMatrixOutputs_andMatrixInput_2_117, response_data_andMatrixOutputs_andMatrixInput_3_117};
  wire [1:0]   response_data_andMatrixOutputs_hi_117 = {response_data_andMatrixOutputs_andMatrixInput_0_117, response_data_andMatrixOutputs_andMatrixInput_1_117};
  wire         response_data_andMatrixOutputs_3_2_23 = &{response_data_andMatrixOutputs_hi_117, response_data_andMatrixOutputs_lo_117};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_118 = response_data_invInputs_23[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_118 = response_data_invInputs_23[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_119 = response_data_invInputs_23[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_118 = response_data_plaInput_23[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_119 = response_data_plaInput_23[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_118 = {response_data_andMatrixOutputs_andMatrixInput_3_118, response_data_andMatrixOutputs_andMatrixInput_4_46};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_46 = {response_data_andMatrixOutputs_andMatrixInput_0_118, response_data_andMatrixOutputs_andMatrixInput_1_118};
  wire [2:0]   response_data_andMatrixOutputs_hi_118 = {response_data_andMatrixOutputs_hi_hi_46, response_data_andMatrixOutputs_andMatrixInput_2_118};
  wire         response_data_andMatrixOutputs_0_2_23 = &{response_data_andMatrixOutputs_hi_118, response_data_andMatrixOutputs_lo_118};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_119 = response_data_invInputs_23[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_119 = {response_data_andMatrixOutputs_andMatrixInput_3_119, response_data_andMatrixOutputs_andMatrixInput_4_47};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_47 = {response_data_andMatrixOutputs_andMatrixInput_0_119, response_data_andMatrixOutputs_andMatrixInput_1_119};
  wire [2:0]   response_data_andMatrixOutputs_hi_119 = {response_data_andMatrixOutputs_hi_hi_47, response_data_andMatrixOutputs_andMatrixInput_2_119};
  wire         response_data_andMatrixOutputs_2_2_23 = &{response_data_andMatrixOutputs_hi_119, response_data_andMatrixOutputs_lo_119};
  wire [1:0]   response_data_orMatrixOutputs_lo_23 = {response_data_andMatrixOutputs_0_2_23, response_data_andMatrixOutputs_2_2_23};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_23 = {response_data_andMatrixOutputs_4_2_23, response_data_andMatrixOutputs_1_2_23};
  wire [2:0]   response_data_orMatrixOutputs_hi_23 = {response_data_orMatrixOutputs_hi_hi_23, response_data_andMatrixOutputs_3_2_23};
  wire         response_data_orMatrixOutputs_23 = |{response_data_orMatrixOutputs_hi_23, response_data_orMatrixOutputs_lo_23};
  assign response_data_invMatrixOutputs_23 = response_data_orMatrixOutputs_23;
  wire         response_data_plaOutput_23 = response_data_invMatrixOutputs_23;
  assign response_data_plaInput_23 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[23], request_src_1[23]};
  wire [4:0]   response_data_plaInput_24;
  wire [4:0]   response_data_invInputs_24 = ~response_data_plaInput_24;
  wire         response_data_invMatrixOutputs_24;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_120 = response_data_plaInput_24[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_121 = response_data_plaInput_24[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_123 = response_data_plaInput_24[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_120 = response_data_plaInput_24[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_122 = response_data_plaInput_24[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_124 = response_data_plaInput_24[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_120 = response_data_invInputs_24[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_121 = response_data_invInputs_24[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_122 = response_data_invInputs_24[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_120 = response_data_invInputs_24[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_121 = response_data_invInputs_24[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_122 = response_data_invInputs_24[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_48 = response_data_invInputs_24[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_49 = response_data_invInputs_24[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_120 = {response_data_andMatrixOutputs_andMatrixInput_2_120, response_data_andMatrixOutputs_andMatrixInput_3_120};
  wire [1:0]   response_data_andMatrixOutputs_hi_120 = {response_data_andMatrixOutputs_andMatrixInput_0_120, response_data_andMatrixOutputs_andMatrixInput_1_120};
  wire         response_data_andMatrixOutputs_4_2_24 = &{response_data_andMatrixOutputs_hi_120, response_data_andMatrixOutputs_lo_120};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_121 = response_data_plaInput_24[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_122 = response_data_plaInput_24[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_121 = {response_data_andMatrixOutputs_andMatrixInput_2_121, response_data_andMatrixOutputs_andMatrixInput_3_121};
  wire [1:0]   response_data_andMatrixOutputs_hi_121 = {response_data_andMatrixOutputs_andMatrixInput_0_121, response_data_andMatrixOutputs_andMatrixInput_1_121};
  wire         response_data_andMatrixOutputs_1_2_24 = &{response_data_andMatrixOutputs_hi_121, response_data_andMatrixOutputs_lo_121};
  wire [1:0]   response_data_andMatrixOutputs_lo_122 = {response_data_andMatrixOutputs_andMatrixInput_2_122, response_data_andMatrixOutputs_andMatrixInput_3_122};
  wire [1:0]   response_data_andMatrixOutputs_hi_122 = {response_data_andMatrixOutputs_andMatrixInput_0_122, response_data_andMatrixOutputs_andMatrixInput_1_122};
  wire         response_data_andMatrixOutputs_3_2_24 = &{response_data_andMatrixOutputs_hi_122, response_data_andMatrixOutputs_lo_122};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_123 = response_data_invInputs_24[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_123 = response_data_invInputs_24[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_124 = response_data_invInputs_24[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_123 = response_data_plaInput_24[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_124 = response_data_plaInput_24[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_123 = {response_data_andMatrixOutputs_andMatrixInput_3_123, response_data_andMatrixOutputs_andMatrixInput_4_48};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_48 = {response_data_andMatrixOutputs_andMatrixInput_0_123, response_data_andMatrixOutputs_andMatrixInput_1_123};
  wire [2:0]   response_data_andMatrixOutputs_hi_123 = {response_data_andMatrixOutputs_hi_hi_48, response_data_andMatrixOutputs_andMatrixInput_2_123};
  wire         response_data_andMatrixOutputs_0_2_24 = &{response_data_andMatrixOutputs_hi_123, response_data_andMatrixOutputs_lo_123};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_124 = response_data_invInputs_24[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_124 = {response_data_andMatrixOutputs_andMatrixInput_3_124, response_data_andMatrixOutputs_andMatrixInput_4_49};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_49 = {response_data_andMatrixOutputs_andMatrixInput_0_124, response_data_andMatrixOutputs_andMatrixInput_1_124};
  wire [2:0]   response_data_andMatrixOutputs_hi_124 = {response_data_andMatrixOutputs_hi_hi_49, response_data_andMatrixOutputs_andMatrixInput_2_124};
  wire         response_data_andMatrixOutputs_2_2_24 = &{response_data_andMatrixOutputs_hi_124, response_data_andMatrixOutputs_lo_124};
  wire [1:0]   response_data_orMatrixOutputs_lo_24 = {response_data_andMatrixOutputs_0_2_24, response_data_andMatrixOutputs_2_2_24};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_24 = {response_data_andMatrixOutputs_4_2_24, response_data_andMatrixOutputs_1_2_24};
  wire [2:0]   response_data_orMatrixOutputs_hi_24 = {response_data_orMatrixOutputs_hi_hi_24, response_data_andMatrixOutputs_3_2_24};
  wire         response_data_orMatrixOutputs_24 = |{response_data_orMatrixOutputs_hi_24, response_data_orMatrixOutputs_lo_24};
  assign response_data_invMatrixOutputs_24 = response_data_orMatrixOutputs_24;
  wire         response_data_plaOutput_24 = response_data_invMatrixOutputs_24;
  assign response_data_plaInput_24 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[24], request_src_1[24]};
  wire [4:0]   response_data_plaInput_25;
  wire [4:0]   response_data_invInputs_25 = ~response_data_plaInput_25;
  wire         response_data_invMatrixOutputs_25;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_125 = response_data_plaInput_25[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_126 = response_data_plaInput_25[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_128 = response_data_plaInput_25[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_125 = response_data_plaInput_25[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_127 = response_data_plaInput_25[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_129 = response_data_plaInput_25[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_125 = response_data_invInputs_25[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_126 = response_data_invInputs_25[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_127 = response_data_invInputs_25[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_125 = response_data_invInputs_25[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_126 = response_data_invInputs_25[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_127 = response_data_invInputs_25[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_50 = response_data_invInputs_25[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_51 = response_data_invInputs_25[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_125 = {response_data_andMatrixOutputs_andMatrixInput_2_125, response_data_andMatrixOutputs_andMatrixInput_3_125};
  wire [1:0]   response_data_andMatrixOutputs_hi_125 = {response_data_andMatrixOutputs_andMatrixInput_0_125, response_data_andMatrixOutputs_andMatrixInput_1_125};
  wire         response_data_andMatrixOutputs_4_2_25 = &{response_data_andMatrixOutputs_hi_125, response_data_andMatrixOutputs_lo_125};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_126 = response_data_plaInput_25[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_127 = response_data_plaInput_25[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_126 = {response_data_andMatrixOutputs_andMatrixInput_2_126, response_data_andMatrixOutputs_andMatrixInput_3_126};
  wire [1:0]   response_data_andMatrixOutputs_hi_126 = {response_data_andMatrixOutputs_andMatrixInput_0_126, response_data_andMatrixOutputs_andMatrixInput_1_126};
  wire         response_data_andMatrixOutputs_1_2_25 = &{response_data_andMatrixOutputs_hi_126, response_data_andMatrixOutputs_lo_126};
  wire [1:0]   response_data_andMatrixOutputs_lo_127 = {response_data_andMatrixOutputs_andMatrixInput_2_127, response_data_andMatrixOutputs_andMatrixInput_3_127};
  wire [1:0]   response_data_andMatrixOutputs_hi_127 = {response_data_andMatrixOutputs_andMatrixInput_0_127, response_data_andMatrixOutputs_andMatrixInput_1_127};
  wire         response_data_andMatrixOutputs_3_2_25 = &{response_data_andMatrixOutputs_hi_127, response_data_andMatrixOutputs_lo_127};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_128 = response_data_invInputs_25[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_128 = response_data_invInputs_25[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_129 = response_data_invInputs_25[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_128 = response_data_plaInput_25[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_129 = response_data_plaInput_25[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_128 = {response_data_andMatrixOutputs_andMatrixInput_3_128, response_data_andMatrixOutputs_andMatrixInput_4_50};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_50 = {response_data_andMatrixOutputs_andMatrixInput_0_128, response_data_andMatrixOutputs_andMatrixInput_1_128};
  wire [2:0]   response_data_andMatrixOutputs_hi_128 = {response_data_andMatrixOutputs_hi_hi_50, response_data_andMatrixOutputs_andMatrixInput_2_128};
  wire         response_data_andMatrixOutputs_0_2_25 = &{response_data_andMatrixOutputs_hi_128, response_data_andMatrixOutputs_lo_128};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_129 = response_data_invInputs_25[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_129 = {response_data_andMatrixOutputs_andMatrixInput_3_129, response_data_andMatrixOutputs_andMatrixInput_4_51};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_51 = {response_data_andMatrixOutputs_andMatrixInput_0_129, response_data_andMatrixOutputs_andMatrixInput_1_129};
  wire [2:0]   response_data_andMatrixOutputs_hi_129 = {response_data_andMatrixOutputs_hi_hi_51, response_data_andMatrixOutputs_andMatrixInput_2_129};
  wire         response_data_andMatrixOutputs_2_2_25 = &{response_data_andMatrixOutputs_hi_129, response_data_andMatrixOutputs_lo_129};
  wire [1:0]   response_data_orMatrixOutputs_lo_25 = {response_data_andMatrixOutputs_0_2_25, response_data_andMatrixOutputs_2_2_25};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_25 = {response_data_andMatrixOutputs_4_2_25, response_data_andMatrixOutputs_1_2_25};
  wire [2:0]   response_data_orMatrixOutputs_hi_25 = {response_data_orMatrixOutputs_hi_hi_25, response_data_andMatrixOutputs_3_2_25};
  wire         response_data_orMatrixOutputs_25 = |{response_data_orMatrixOutputs_hi_25, response_data_orMatrixOutputs_lo_25};
  assign response_data_invMatrixOutputs_25 = response_data_orMatrixOutputs_25;
  wire         response_data_plaOutput_25 = response_data_invMatrixOutputs_25;
  assign response_data_plaInput_25 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[25], request_src_1[25]};
  wire [4:0]   response_data_plaInput_26;
  wire [4:0]   response_data_invInputs_26 = ~response_data_plaInput_26;
  wire         response_data_invMatrixOutputs_26;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_130 = response_data_plaInput_26[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_131 = response_data_plaInput_26[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_133 = response_data_plaInput_26[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_130 = response_data_plaInput_26[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_132 = response_data_plaInput_26[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_134 = response_data_plaInput_26[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_130 = response_data_invInputs_26[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_131 = response_data_invInputs_26[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_132 = response_data_invInputs_26[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_130 = response_data_invInputs_26[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_131 = response_data_invInputs_26[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_132 = response_data_invInputs_26[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_52 = response_data_invInputs_26[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_53 = response_data_invInputs_26[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_130 = {response_data_andMatrixOutputs_andMatrixInput_2_130, response_data_andMatrixOutputs_andMatrixInput_3_130};
  wire [1:0]   response_data_andMatrixOutputs_hi_130 = {response_data_andMatrixOutputs_andMatrixInput_0_130, response_data_andMatrixOutputs_andMatrixInput_1_130};
  wire         response_data_andMatrixOutputs_4_2_26 = &{response_data_andMatrixOutputs_hi_130, response_data_andMatrixOutputs_lo_130};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_131 = response_data_plaInput_26[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_132 = response_data_plaInput_26[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_131 = {response_data_andMatrixOutputs_andMatrixInput_2_131, response_data_andMatrixOutputs_andMatrixInput_3_131};
  wire [1:0]   response_data_andMatrixOutputs_hi_131 = {response_data_andMatrixOutputs_andMatrixInput_0_131, response_data_andMatrixOutputs_andMatrixInput_1_131};
  wire         response_data_andMatrixOutputs_1_2_26 = &{response_data_andMatrixOutputs_hi_131, response_data_andMatrixOutputs_lo_131};
  wire [1:0]   response_data_andMatrixOutputs_lo_132 = {response_data_andMatrixOutputs_andMatrixInput_2_132, response_data_andMatrixOutputs_andMatrixInput_3_132};
  wire [1:0]   response_data_andMatrixOutputs_hi_132 = {response_data_andMatrixOutputs_andMatrixInput_0_132, response_data_andMatrixOutputs_andMatrixInput_1_132};
  wire         response_data_andMatrixOutputs_3_2_26 = &{response_data_andMatrixOutputs_hi_132, response_data_andMatrixOutputs_lo_132};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_133 = response_data_invInputs_26[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_133 = response_data_invInputs_26[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_134 = response_data_invInputs_26[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_133 = response_data_plaInput_26[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_134 = response_data_plaInput_26[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_133 = {response_data_andMatrixOutputs_andMatrixInput_3_133, response_data_andMatrixOutputs_andMatrixInput_4_52};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_52 = {response_data_andMatrixOutputs_andMatrixInput_0_133, response_data_andMatrixOutputs_andMatrixInput_1_133};
  wire [2:0]   response_data_andMatrixOutputs_hi_133 = {response_data_andMatrixOutputs_hi_hi_52, response_data_andMatrixOutputs_andMatrixInput_2_133};
  wire         response_data_andMatrixOutputs_0_2_26 = &{response_data_andMatrixOutputs_hi_133, response_data_andMatrixOutputs_lo_133};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_134 = response_data_invInputs_26[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_134 = {response_data_andMatrixOutputs_andMatrixInput_3_134, response_data_andMatrixOutputs_andMatrixInput_4_53};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_53 = {response_data_andMatrixOutputs_andMatrixInput_0_134, response_data_andMatrixOutputs_andMatrixInput_1_134};
  wire [2:0]   response_data_andMatrixOutputs_hi_134 = {response_data_andMatrixOutputs_hi_hi_53, response_data_andMatrixOutputs_andMatrixInput_2_134};
  wire         response_data_andMatrixOutputs_2_2_26 = &{response_data_andMatrixOutputs_hi_134, response_data_andMatrixOutputs_lo_134};
  wire [1:0]   response_data_orMatrixOutputs_lo_26 = {response_data_andMatrixOutputs_0_2_26, response_data_andMatrixOutputs_2_2_26};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_26 = {response_data_andMatrixOutputs_4_2_26, response_data_andMatrixOutputs_1_2_26};
  wire [2:0]   response_data_orMatrixOutputs_hi_26 = {response_data_orMatrixOutputs_hi_hi_26, response_data_andMatrixOutputs_3_2_26};
  wire         response_data_orMatrixOutputs_26 = |{response_data_orMatrixOutputs_hi_26, response_data_orMatrixOutputs_lo_26};
  assign response_data_invMatrixOutputs_26 = response_data_orMatrixOutputs_26;
  wire         response_data_plaOutput_26 = response_data_invMatrixOutputs_26;
  assign response_data_plaInput_26 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[26], request_src_1[26]};
  wire [4:0]   response_data_plaInput_27;
  wire [4:0]   response_data_invInputs_27 = ~response_data_plaInput_27;
  wire         response_data_invMatrixOutputs_27;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_135 = response_data_plaInput_27[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_136 = response_data_plaInput_27[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_138 = response_data_plaInput_27[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_135 = response_data_plaInput_27[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_137 = response_data_plaInput_27[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_139 = response_data_plaInput_27[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_135 = response_data_invInputs_27[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_136 = response_data_invInputs_27[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_137 = response_data_invInputs_27[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_135 = response_data_invInputs_27[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_136 = response_data_invInputs_27[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_137 = response_data_invInputs_27[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_54 = response_data_invInputs_27[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_55 = response_data_invInputs_27[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_135 = {response_data_andMatrixOutputs_andMatrixInput_2_135, response_data_andMatrixOutputs_andMatrixInput_3_135};
  wire [1:0]   response_data_andMatrixOutputs_hi_135 = {response_data_andMatrixOutputs_andMatrixInput_0_135, response_data_andMatrixOutputs_andMatrixInput_1_135};
  wire         response_data_andMatrixOutputs_4_2_27 = &{response_data_andMatrixOutputs_hi_135, response_data_andMatrixOutputs_lo_135};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_136 = response_data_plaInput_27[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_137 = response_data_plaInput_27[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_136 = {response_data_andMatrixOutputs_andMatrixInput_2_136, response_data_andMatrixOutputs_andMatrixInput_3_136};
  wire [1:0]   response_data_andMatrixOutputs_hi_136 = {response_data_andMatrixOutputs_andMatrixInput_0_136, response_data_andMatrixOutputs_andMatrixInput_1_136};
  wire         response_data_andMatrixOutputs_1_2_27 = &{response_data_andMatrixOutputs_hi_136, response_data_andMatrixOutputs_lo_136};
  wire [1:0]   response_data_andMatrixOutputs_lo_137 = {response_data_andMatrixOutputs_andMatrixInput_2_137, response_data_andMatrixOutputs_andMatrixInput_3_137};
  wire [1:0]   response_data_andMatrixOutputs_hi_137 = {response_data_andMatrixOutputs_andMatrixInput_0_137, response_data_andMatrixOutputs_andMatrixInput_1_137};
  wire         response_data_andMatrixOutputs_3_2_27 = &{response_data_andMatrixOutputs_hi_137, response_data_andMatrixOutputs_lo_137};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_138 = response_data_invInputs_27[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_138 = response_data_invInputs_27[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_139 = response_data_invInputs_27[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_138 = response_data_plaInput_27[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_139 = response_data_plaInput_27[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_138 = {response_data_andMatrixOutputs_andMatrixInput_3_138, response_data_andMatrixOutputs_andMatrixInput_4_54};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_54 = {response_data_andMatrixOutputs_andMatrixInput_0_138, response_data_andMatrixOutputs_andMatrixInput_1_138};
  wire [2:0]   response_data_andMatrixOutputs_hi_138 = {response_data_andMatrixOutputs_hi_hi_54, response_data_andMatrixOutputs_andMatrixInput_2_138};
  wire         response_data_andMatrixOutputs_0_2_27 = &{response_data_andMatrixOutputs_hi_138, response_data_andMatrixOutputs_lo_138};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_139 = response_data_invInputs_27[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_139 = {response_data_andMatrixOutputs_andMatrixInput_3_139, response_data_andMatrixOutputs_andMatrixInput_4_55};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_55 = {response_data_andMatrixOutputs_andMatrixInput_0_139, response_data_andMatrixOutputs_andMatrixInput_1_139};
  wire [2:0]   response_data_andMatrixOutputs_hi_139 = {response_data_andMatrixOutputs_hi_hi_55, response_data_andMatrixOutputs_andMatrixInput_2_139};
  wire         response_data_andMatrixOutputs_2_2_27 = &{response_data_andMatrixOutputs_hi_139, response_data_andMatrixOutputs_lo_139};
  wire [1:0]   response_data_orMatrixOutputs_lo_27 = {response_data_andMatrixOutputs_0_2_27, response_data_andMatrixOutputs_2_2_27};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_27 = {response_data_andMatrixOutputs_4_2_27, response_data_andMatrixOutputs_1_2_27};
  wire [2:0]   response_data_orMatrixOutputs_hi_27 = {response_data_orMatrixOutputs_hi_hi_27, response_data_andMatrixOutputs_3_2_27};
  wire         response_data_orMatrixOutputs_27 = |{response_data_orMatrixOutputs_hi_27, response_data_orMatrixOutputs_lo_27};
  assign response_data_invMatrixOutputs_27 = response_data_orMatrixOutputs_27;
  wire         response_data_plaOutput_27 = response_data_invMatrixOutputs_27;
  assign response_data_plaInput_27 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[27], request_src_1[27]};
  wire [4:0]   response_data_plaInput_28;
  wire [4:0]   response_data_invInputs_28 = ~response_data_plaInput_28;
  wire         response_data_invMatrixOutputs_28;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_140 = response_data_plaInput_28[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_141 = response_data_plaInput_28[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_143 = response_data_plaInput_28[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_140 = response_data_plaInput_28[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_142 = response_data_plaInput_28[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_144 = response_data_plaInput_28[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_140 = response_data_invInputs_28[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_141 = response_data_invInputs_28[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_142 = response_data_invInputs_28[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_140 = response_data_invInputs_28[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_141 = response_data_invInputs_28[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_142 = response_data_invInputs_28[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_56 = response_data_invInputs_28[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_57 = response_data_invInputs_28[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_140 = {response_data_andMatrixOutputs_andMatrixInput_2_140, response_data_andMatrixOutputs_andMatrixInput_3_140};
  wire [1:0]   response_data_andMatrixOutputs_hi_140 = {response_data_andMatrixOutputs_andMatrixInput_0_140, response_data_andMatrixOutputs_andMatrixInput_1_140};
  wire         response_data_andMatrixOutputs_4_2_28 = &{response_data_andMatrixOutputs_hi_140, response_data_andMatrixOutputs_lo_140};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_141 = response_data_plaInput_28[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_142 = response_data_plaInput_28[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_141 = {response_data_andMatrixOutputs_andMatrixInput_2_141, response_data_andMatrixOutputs_andMatrixInput_3_141};
  wire [1:0]   response_data_andMatrixOutputs_hi_141 = {response_data_andMatrixOutputs_andMatrixInput_0_141, response_data_andMatrixOutputs_andMatrixInput_1_141};
  wire         response_data_andMatrixOutputs_1_2_28 = &{response_data_andMatrixOutputs_hi_141, response_data_andMatrixOutputs_lo_141};
  wire [1:0]   response_data_andMatrixOutputs_lo_142 = {response_data_andMatrixOutputs_andMatrixInput_2_142, response_data_andMatrixOutputs_andMatrixInput_3_142};
  wire [1:0]   response_data_andMatrixOutputs_hi_142 = {response_data_andMatrixOutputs_andMatrixInput_0_142, response_data_andMatrixOutputs_andMatrixInput_1_142};
  wire         response_data_andMatrixOutputs_3_2_28 = &{response_data_andMatrixOutputs_hi_142, response_data_andMatrixOutputs_lo_142};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_143 = response_data_invInputs_28[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_143 = response_data_invInputs_28[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_144 = response_data_invInputs_28[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_143 = response_data_plaInput_28[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_144 = response_data_plaInput_28[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_143 = {response_data_andMatrixOutputs_andMatrixInput_3_143, response_data_andMatrixOutputs_andMatrixInput_4_56};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_56 = {response_data_andMatrixOutputs_andMatrixInput_0_143, response_data_andMatrixOutputs_andMatrixInput_1_143};
  wire [2:0]   response_data_andMatrixOutputs_hi_143 = {response_data_andMatrixOutputs_hi_hi_56, response_data_andMatrixOutputs_andMatrixInput_2_143};
  wire         response_data_andMatrixOutputs_0_2_28 = &{response_data_andMatrixOutputs_hi_143, response_data_andMatrixOutputs_lo_143};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_144 = response_data_invInputs_28[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_144 = {response_data_andMatrixOutputs_andMatrixInput_3_144, response_data_andMatrixOutputs_andMatrixInput_4_57};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_57 = {response_data_andMatrixOutputs_andMatrixInput_0_144, response_data_andMatrixOutputs_andMatrixInput_1_144};
  wire [2:0]   response_data_andMatrixOutputs_hi_144 = {response_data_andMatrixOutputs_hi_hi_57, response_data_andMatrixOutputs_andMatrixInput_2_144};
  wire         response_data_andMatrixOutputs_2_2_28 = &{response_data_andMatrixOutputs_hi_144, response_data_andMatrixOutputs_lo_144};
  wire [1:0]   response_data_orMatrixOutputs_lo_28 = {response_data_andMatrixOutputs_0_2_28, response_data_andMatrixOutputs_2_2_28};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_28 = {response_data_andMatrixOutputs_4_2_28, response_data_andMatrixOutputs_1_2_28};
  wire [2:0]   response_data_orMatrixOutputs_hi_28 = {response_data_orMatrixOutputs_hi_hi_28, response_data_andMatrixOutputs_3_2_28};
  wire         response_data_orMatrixOutputs_28 = |{response_data_orMatrixOutputs_hi_28, response_data_orMatrixOutputs_lo_28};
  assign response_data_invMatrixOutputs_28 = response_data_orMatrixOutputs_28;
  wire         response_data_plaOutput_28 = response_data_invMatrixOutputs_28;
  assign response_data_plaInput_28 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[28], request_src_1[28]};
  wire [4:0]   response_data_plaInput_29;
  wire [4:0]   response_data_invInputs_29 = ~response_data_plaInput_29;
  wire         response_data_invMatrixOutputs_29;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_145 = response_data_plaInput_29[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_146 = response_data_plaInput_29[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_148 = response_data_plaInput_29[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_145 = response_data_plaInput_29[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_147 = response_data_plaInput_29[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_149 = response_data_plaInput_29[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_145 = response_data_invInputs_29[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_146 = response_data_invInputs_29[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_147 = response_data_invInputs_29[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_145 = response_data_invInputs_29[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_146 = response_data_invInputs_29[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_147 = response_data_invInputs_29[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_58 = response_data_invInputs_29[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_59 = response_data_invInputs_29[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_145 = {response_data_andMatrixOutputs_andMatrixInput_2_145, response_data_andMatrixOutputs_andMatrixInput_3_145};
  wire [1:0]   response_data_andMatrixOutputs_hi_145 = {response_data_andMatrixOutputs_andMatrixInput_0_145, response_data_andMatrixOutputs_andMatrixInput_1_145};
  wire         response_data_andMatrixOutputs_4_2_29 = &{response_data_andMatrixOutputs_hi_145, response_data_andMatrixOutputs_lo_145};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_146 = response_data_plaInput_29[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_147 = response_data_plaInput_29[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_146 = {response_data_andMatrixOutputs_andMatrixInput_2_146, response_data_andMatrixOutputs_andMatrixInput_3_146};
  wire [1:0]   response_data_andMatrixOutputs_hi_146 = {response_data_andMatrixOutputs_andMatrixInput_0_146, response_data_andMatrixOutputs_andMatrixInput_1_146};
  wire         response_data_andMatrixOutputs_1_2_29 = &{response_data_andMatrixOutputs_hi_146, response_data_andMatrixOutputs_lo_146};
  wire [1:0]   response_data_andMatrixOutputs_lo_147 = {response_data_andMatrixOutputs_andMatrixInput_2_147, response_data_andMatrixOutputs_andMatrixInput_3_147};
  wire [1:0]   response_data_andMatrixOutputs_hi_147 = {response_data_andMatrixOutputs_andMatrixInput_0_147, response_data_andMatrixOutputs_andMatrixInput_1_147};
  wire         response_data_andMatrixOutputs_3_2_29 = &{response_data_andMatrixOutputs_hi_147, response_data_andMatrixOutputs_lo_147};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_148 = response_data_invInputs_29[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_148 = response_data_invInputs_29[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_149 = response_data_invInputs_29[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_148 = response_data_plaInput_29[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_149 = response_data_plaInput_29[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_148 = {response_data_andMatrixOutputs_andMatrixInput_3_148, response_data_andMatrixOutputs_andMatrixInput_4_58};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_58 = {response_data_andMatrixOutputs_andMatrixInput_0_148, response_data_andMatrixOutputs_andMatrixInput_1_148};
  wire [2:0]   response_data_andMatrixOutputs_hi_148 = {response_data_andMatrixOutputs_hi_hi_58, response_data_andMatrixOutputs_andMatrixInput_2_148};
  wire         response_data_andMatrixOutputs_0_2_29 = &{response_data_andMatrixOutputs_hi_148, response_data_andMatrixOutputs_lo_148};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_149 = response_data_invInputs_29[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_149 = {response_data_andMatrixOutputs_andMatrixInput_3_149, response_data_andMatrixOutputs_andMatrixInput_4_59};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_59 = {response_data_andMatrixOutputs_andMatrixInput_0_149, response_data_andMatrixOutputs_andMatrixInput_1_149};
  wire [2:0]   response_data_andMatrixOutputs_hi_149 = {response_data_andMatrixOutputs_hi_hi_59, response_data_andMatrixOutputs_andMatrixInput_2_149};
  wire         response_data_andMatrixOutputs_2_2_29 = &{response_data_andMatrixOutputs_hi_149, response_data_andMatrixOutputs_lo_149};
  wire [1:0]   response_data_orMatrixOutputs_lo_29 = {response_data_andMatrixOutputs_0_2_29, response_data_andMatrixOutputs_2_2_29};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_29 = {response_data_andMatrixOutputs_4_2_29, response_data_andMatrixOutputs_1_2_29};
  wire [2:0]   response_data_orMatrixOutputs_hi_29 = {response_data_orMatrixOutputs_hi_hi_29, response_data_andMatrixOutputs_3_2_29};
  wire         response_data_orMatrixOutputs_29 = |{response_data_orMatrixOutputs_hi_29, response_data_orMatrixOutputs_lo_29};
  assign response_data_invMatrixOutputs_29 = response_data_orMatrixOutputs_29;
  wire         response_data_plaOutput_29 = response_data_invMatrixOutputs_29;
  assign response_data_plaInput_29 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[29], request_src_1[29]};
  wire [4:0]   response_data_plaInput_30;
  wire [4:0]   response_data_invInputs_30 = ~response_data_plaInput_30;
  wire         response_data_invMatrixOutputs_30;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_150 = response_data_plaInput_30[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_151 = response_data_plaInput_30[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_153 = response_data_plaInput_30[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_150 = response_data_plaInput_30[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_152 = response_data_plaInput_30[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_154 = response_data_plaInput_30[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_150 = response_data_invInputs_30[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_151 = response_data_invInputs_30[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_152 = response_data_invInputs_30[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_150 = response_data_invInputs_30[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_151 = response_data_invInputs_30[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_152 = response_data_invInputs_30[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_60 = response_data_invInputs_30[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_61 = response_data_invInputs_30[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_150 = {response_data_andMatrixOutputs_andMatrixInput_2_150, response_data_andMatrixOutputs_andMatrixInput_3_150};
  wire [1:0]   response_data_andMatrixOutputs_hi_150 = {response_data_andMatrixOutputs_andMatrixInput_0_150, response_data_andMatrixOutputs_andMatrixInput_1_150};
  wire         response_data_andMatrixOutputs_4_2_30 = &{response_data_andMatrixOutputs_hi_150, response_data_andMatrixOutputs_lo_150};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_151 = response_data_plaInput_30[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_152 = response_data_plaInput_30[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_151 = {response_data_andMatrixOutputs_andMatrixInput_2_151, response_data_andMatrixOutputs_andMatrixInput_3_151};
  wire [1:0]   response_data_andMatrixOutputs_hi_151 = {response_data_andMatrixOutputs_andMatrixInput_0_151, response_data_andMatrixOutputs_andMatrixInput_1_151};
  wire         response_data_andMatrixOutputs_1_2_30 = &{response_data_andMatrixOutputs_hi_151, response_data_andMatrixOutputs_lo_151};
  wire [1:0]   response_data_andMatrixOutputs_lo_152 = {response_data_andMatrixOutputs_andMatrixInput_2_152, response_data_andMatrixOutputs_andMatrixInput_3_152};
  wire [1:0]   response_data_andMatrixOutputs_hi_152 = {response_data_andMatrixOutputs_andMatrixInput_0_152, response_data_andMatrixOutputs_andMatrixInput_1_152};
  wire         response_data_andMatrixOutputs_3_2_30 = &{response_data_andMatrixOutputs_hi_152, response_data_andMatrixOutputs_lo_152};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_153 = response_data_invInputs_30[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_153 = response_data_invInputs_30[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_154 = response_data_invInputs_30[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_153 = response_data_plaInput_30[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_154 = response_data_plaInput_30[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_153 = {response_data_andMatrixOutputs_andMatrixInput_3_153, response_data_andMatrixOutputs_andMatrixInput_4_60};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_60 = {response_data_andMatrixOutputs_andMatrixInput_0_153, response_data_andMatrixOutputs_andMatrixInput_1_153};
  wire [2:0]   response_data_andMatrixOutputs_hi_153 = {response_data_andMatrixOutputs_hi_hi_60, response_data_andMatrixOutputs_andMatrixInput_2_153};
  wire         response_data_andMatrixOutputs_0_2_30 = &{response_data_andMatrixOutputs_hi_153, response_data_andMatrixOutputs_lo_153};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_154 = response_data_invInputs_30[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_154 = {response_data_andMatrixOutputs_andMatrixInput_3_154, response_data_andMatrixOutputs_andMatrixInput_4_61};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_61 = {response_data_andMatrixOutputs_andMatrixInput_0_154, response_data_andMatrixOutputs_andMatrixInput_1_154};
  wire [2:0]   response_data_andMatrixOutputs_hi_154 = {response_data_andMatrixOutputs_hi_hi_61, response_data_andMatrixOutputs_andMatrixInput_2_154};
  wire         response_data_andMatrixOutputs_2_2_30 = &{response_data_andMatrixOutputs_hi_154, response_data_andMatrixOutputs_lo_154};
  wire [1:0]   response_data_orMatrixOutputs_lo_30 = {response_data_andMatrixOutputs_0_2_30, response_data_andMatrixOutputs_2_2_30};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_30 = {response_data_andMatrixOutputs_4_2_30, response_data_andMatrixOutputs_1_2_30};
  wire [2:0]   response_data_orMatrixOutputs_hi_30 = {response_data_orMatrixOutputs_hi_hi_30, response_data_andMatrixOutputs_3_2_30};
  wire         response_data_orMatrixOutputs_30 = |{response_data_orMatrixOutputs_hi_30, response_data_orMatrixOutputs_lo_30};
  assign response_data_invMatrixOutputs_30 = response_data_orMatrixOutputs_30;
  wire         response_data_plaOutput_30 = response_data_invMatrixOutputs_30;
  assign response_data_plaInput_30 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[30], request_src_1[30]};
  wire [4:0]   response_data_plaInput_31;
  wire [4:0]   response_data_invInputs_31 = ~response_data_plaInput_31;
  wire         response_data_invMatrixOutputs_31;
  wire         response_data_andMatrixOutputs_andMatrixInput_0_155 = response_data_plaInput_31[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_156 = response_data_plaInput_31[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_158 = response_data_plaInput_31[0];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_155 = response_data_plaInput_31[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_0_157 = response_data_plaInput_31[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_159 = response_data_plaInput_31[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_155 = response_data_invInputs_31[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_156 = response_data_invInputs_31[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_157 = response_data_invInputs_31[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_155 = response_data_invInputs_31[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_156 = response_data_invInputs_31[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_157 = response_data_invInputs_31[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_62 = response_data_invInputs_31[4];
  wire         response_data_andMatrixOutputs_andMatrixInput_4_63 = response_data_invInputs_31[4];
  wire [1:0]   response_data_andMatrixOutputs_lo_155 = {response_data_andMatrixOutputs_andMatrixInput_2_155, response_data_andMatrixOutputs_andMatrixInput_3_155};
  wire [1:0]   response_data_andMatrixOutputs_hi_155 = {response_data_andMatrixOutputs_andMatrixInput_0_155, response_data_andMatrixOutputs_andMatrixInput_1_155};
  wire         response_data_andMatrixOutputs_4_2_31 = &{response_data_andMatrixOutputs_hi_155, response_data_andMatrixOutputs_lo_155};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_156 = response_data_plaInput_31[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_1_157 = response_data_plaInput_31[2];
  wire [1:0]   response_data_andMatrixOutputs_lo_156 = {response_data_andMatrixOutputs_andMatrixInput_2_156, response_data_andMatrixOutputs_andMatrixInput_3_156};
  wire [1:0]   response_data_andMatrixOutputs_hi_156 = {response_data_andMatrixOutputs_andMatrixInput_0_156, response_data_andMatrixOutputs_andMatrixInput_1_156};
  wire         response_data_andMatrixOutputs_1_2_31 = &{response_data_andMatrixOutputs_hi_156, response_data_andMatrixOutputs_lo_156};
  wire [1:0]   response_data_andMatrixOutputs_lo_157 = {response_data_andMatrixOutputs_andMatrixInput_2_157, response_data_andMatrixOutputs_andMatrixInput_3_157};
  wire [1:0]   response_data_andMatrixOutputs_hi_157 = {response_data_andMatrixOutputs_andMatrixInput_0_157, response_data_andMatrixOutputs_andMatrixInput_1_157};
  wire         response_data_andMatrixOutputs_3_2_31 = &{response_data_andMatrixOutputs_hi_157, response_data_andMatrixOutputs_lo_157};
  wire         response_data_andMatrixOutputs_andMatrixInput_1_158 = response_data_invInputs_31[1];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_158 = response_data_invInputs_31[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_2_159 = response_data_invInputs_31[2];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_158 = response_data_plaInput_31[3];
  wire         response_data_andMatrixOutputs_andMatrixInput_3_159 = response_data_plaInput_31[3];
  wire [1:0]   response_data_andMatrixOutputs_lo_158 = {response_data_andMatrixOutputs_andMatrixInput_3_158, response_data_andMatrixOutputs_andMatrixInput_4_62};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_62 = {response_data_andMatrixOutputs_andMatrixInput_0_158, response_data_andMatrixOutputs_andMatrixInput_1_158};
  wire [2:0]   response_data_andMatrixOutputs_hi_158 = {response_data_andMatrixOutputs_hi_hi_62, response_data_andMatrixOutputs_andMatrixInput_2_158};
  wire         response_data_andMatrixOutputs_0_2_31 = &{response_data_andMatrixOutputs_hi_158, response_data_andMatrixOutputs_lo_158};
  wire         response_data_andMatrixOutputs_andMatrixInput_0_159 = response_data_invInputs_31[0];
  wire [1:0]   response_data_andMatrixOutputs_lo_159 = {response_data_andMatrixOutputs_andMatrixInput_3_159, response_data_andMatrixOutputs_andMatrixInput_4_63};
  wire [1:0]   response_data_andMatrixOutputs_hi_hi_63 = {response_data_andMatrixOutputs_andMatrixInput_0_159, response_data_andMatrixOutputs_andMatrixInput_1_159};
  wire [2:0]   response_data_andMatrixOutputs_hi_159 = {response_data_andMatrixOutputs_hi_hi_63, response_data_andMatrixOutputs_andMatrixInput_2_159};
  wire         response_data_andMatrixOutputs_2_2_31 = &{response_data_andMatrixOutputs_hi_159, response_data_andMatrixOutputs_lo_159};
  wire [1:0]   response_data_orMatrixOutputs_lo_31 = {response_data_andMatrixOutputs_0_2_31, response_data_andMatrixOutputs_2_2_31};
  wire [1:0]   response_data_orMatrixOutputs_hi_hi_31 = {response_data_andMatrixOutputs_4_2_31, response_data_andMatrixOutputs_1_2_31};
  wire [2:0]   response_data_orMatrixOutputs_hi_31 = {response_data_orMatrixOutputs_hi_hi_31, response_data_andMatrixOutputs_3_2_31};
  wire         response_data_orMatrixOutputs_31 = |{response_data_orMatrixOutputs_hi_31, response_data_orMatrixOutputs_lo_31};
  assign response_data_invMatrixOutputs_31 = response_data_orMatrixOutputs_31;
  wire         response_data_plaOutput_31 = response_data_invMatrixOutputs_31;
  assign response_data_plaInput_31 = {1'h0, request_opcode[1:0], request_opcode[2] ^ request_src_0[31], request_src_1[31]};
  wire [1:0]   response_data_lo_lo_lo_lo = {request_src_3[1] ? response_data_plaOutput_1 ^ request_opcode[3] : request_src_2[1], request_src_3[0] ? response_data_plaOutput ^ request_opcode[3] : request_src_2[0]};
  wire [1:0]   response_data_lo_lo_lo_hi = {request_src_3[3] ? response_data_plaOutput_3 ^ request_opcode[3] : request_src_2[3], request_src_3[2] ? response_data_plaOutput_2 ^ request_opcode[3] : request_src_2[2]};
  wire [3:0]   response_data_lo_lo_lo = {response_data_lo_lo_lo_hi, response_data_lo_lo_lo_lo};
  wire [1:0]   response_data_lo_lo_hi_lo = {request_src_3[5] ? response_data_plaOutput_5 ^ request_opcode[3] : request_src_2[5], request_src_3[4] ? response_data_plaOutput_4 ^ request_opcode[3] : request_src_2[4]};
  wire [1:0]   response_data_lo_lo_hi_hi = {request_src_3[7] ? response_data_plaOutput_7 ^ request_opcode[3] : request_src_2[7], request_src_3[6] ? response_data_plaOutput_6 ^ request_opcode[3] : request_src_2[6]};
  wire [3:0]   response_data_lo_lo_hi = {response_data_lo_lo_hi_hi, response_data_lo_lo_hi_lo};
  wire [7:0]   response_data_lo_lo = {response_data_lo_lo_hi, response_data_lo_lo_lo};
  wire [1:0]   response_data_lo_hi_lo_lo = {request_src_3[9] ? response_data_plaOutput_9 ^ request_opcode[3] : request_src_2[9], request_src_3[8] ? response_data_plaOutput_8 ^ request_opcode[3] : request_src_2[8]};
  wire [1:0]   response_data_lo_hi_lo_hi = {request_src_3[11] ? response_data_plaOutput_11 ^ request_opcode[3] : request_src_2[11], request_src_3[10] ? response_data_plaOutput_10 ^ request_opcode[3] : request_src_2[10]};
  wire [3:0]   response_data_lo_hi_lo = {response_data_lo_hi_lo_hi, response_data_lo_hi_lo_lo};
  wire [1:0]   response_data_lo_hi_hi_lo = {request_src_3[13] ? response_data_plaOutput_13 ^ request_opcode[3] : request_src_2[13], request_src_3[12] ? response_data_plaOutput_12 ^ request_opcode[3] : request_src_2[12]};
  wire [1:0]   response_data_lo_hi_hi_hi = {request_src_3[15] ? response_data_plaOutput_15 ^ request_opcode[3] : request_src_2[15], request_src_3[14] ? response_data_plaOutput_14 ^ request_opcode[3] : request_src_2[14]};
  wire [3:0]   response_data_lo_hi_hi = {response_data_lo_hi_hi_hi, response_data_lo_hi_hi_lo};
  wire [7:0]   response_data_lo_hi = {response_data_lo_hi_hi, response_data_lo_hi_lo};
  wire [15:0]  response_data_lo = {response_data_lo_hi, response_data_lo_lo};
  wire [1:0]   response_data_hi_lo_lo_lo = {request_src_3[17] ? response_data_plaOutput_17 ^ request_opcode[3] : request_src_2[17], request_src_3[16] ? response_data_plaOutput_16 ^ request_opcode[3] : request_src_2[16]};
  wire [1:0]   response_data_hi_lo_lo_hi = {request_src_3[19] ? response_data_plaOutput_19 ^ request_opcode[3] : request_src_2[19], request_src_3[18] ? response_data_plaOutput_18 ^ request_opcode[3] : request_src_2[18]};
  wire [3:0]   response_data_hi_lo_lo = {response_data_hi_lo_lo_hi, response_data_hi_lo_lo_lo};
  wire [1:0]   response_data_hi_lo_hi_lo = {request_src_3[21] ? response_data_plaOutput_21 ^ request_opcode[3] : request_src_2[21], request_src_3[20] ? response_data_plaOutput_20 ^ request_opcode[3] : request_src_2[20]};
  wire [1:0]   response_data_hi_lo_hi_hi = {request_src_3[23] ? response_data_plaOutput_23 ^ request_opcode[3] : request_src_2[23], request_src_3[22] ? response_data_plaOutput_22 ^ request_opcode[3] : request_src_2[22]};
  wire [3:0]   response_data_hi_lo_hi = {response_data_hi_lo_hi_hi, response_data_hi_lo_hi_lo};
  wire [7:0]   response_data_hi_lo = {response_data_hi_lo_hi, response_data_hi_lo_lo};
  wire [1:0]   response_data_hi_hi_lo_lo = {request_src_3[25] ? response_data_plaOutput_25 ^ request_opcode[3] : request_src_2[25], request_src_3[24] ? response_data_plaOutput_24 ^ request_opcode[3] : request_src_2[24]};
  wire [1:0]   response_data_hi_hi_lo_hi = {request_src_3[27] ? response_data_plaOutput_27 ^ request_opcode[3] : request_src_2[27], request_src_3[26] ? response_data_plaOutput_26 ^ request_opcode[3] : request_src_2[26]};
  wire [3:0]   response_data_hi_hi_lo = {response_data_hi_hi_lo_hi, response_data_hi_hi_lo_lo};
  wire [1:0]   response_data_hi_hi_hi_lo = {request_src_3[29] ? response_data_plaOutput_29 ^ request_opcode[3] : request_src_2[29], request_src_3[28] ? response_data_plaOutput_28 ^ request_opcode[3] : request_src_2[28]};
  wire [1:0]   response_data_hi_hi_hi_hi = {request_src_3[31] ? response_data_plaOutput_31 ^ request_opcode[3] : request_src_2[31], request_src_3[30] ? response_data_plaOutput_30 ^ request_opcode[3] : request_src_2[30]};
  wire [3:0]   response_data_hi_hi_hi = {response_data_hi_hi_hi_hi, response_data_hi_hi_hi_lo};
  wire [7:0]   response_data_hi_hi = {response_data_hi_hi_hi, response_data_hi_hi_lo};
  wire [15:0]  response_data_hi = {response_data_hi_hi, response_data_hi_lo};
  assign response_data = {response_data_hi, response_data_lo};
  always @(posedge clock) begin
    if (reset) begin
      requestReg_tag <= 2'h0;
      requestReg_src_0 <= 32'h0;
      requestReg_src_1 <= 32'h0;
      requestReg_src_2 <= 32'h0;
      requestReg_src_3 <= 32'h0;
      requestReg_opcode <= 4'h0;
      requestRegValid <= 1'h0;
      request_pipeResponse_pipe_v <= 1'h0;
    end
    else begin
      if (requestIO_valid_0) begin
        requestReg_tag <= requestIO_bits_tag_0;
        requestReg_src_0 <= requestIO_bits_src_0_0;
        requestReg_src_1 <= requestIO_bits_src_1_0;
        requestReg_src_2 <= requestIO_bits_src_2_0;
        requestReg_src_3 <= requestIO_bits_src_3_0;
        requestReg_opcode <= requestIO_bits_opcode_0;
      end
      requestRegValid <= requestIO_valid_0;
      request_pipeResponse_pipe_v <= request_responseValidWire;
    end
    if (request_responseValidWire) begin
      request_pipeResponse_pipe_b_tag <= request_responseWire_tag;
      request_pipeResponse_pipe_b_data <= request_responseWire_data;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:5];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [2:0] i = 3'h0; i < 3'h6; i += 3'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        requestReg_tag = _RANDOM[3'h0][1:0];
        requestReg_src_0 = {_RANDOM[3'h0][31:2], _RANDOM[3'h1][1:0]};
        requestReg_src_1 = {_RANDOM[3'h1][31:2], _RANDOM[3'h2][1:0]};
        requestReg_src_2 = {_RANDOM[3'h2][31:2], _RANDOM[3'h3][1:0]};
        requestReg_src_3 = {_RANDOM[3'h3][31:2], _RANDOM[3'h4][1:0]};
        requestReg_opcode = _RANDOM[3'h4][5:2];
        requestRegValid = _RANDOM[3'h4][6];
        request_pipeResponse_pipe_v = _RANDOM[3'h4][7];
        request_pipeResponse_pipe_b_tag = _RANDOM[3'h4][9:8];
        request_pipeResponse_pipe_b_data = {_RANDOM[3'h4][31:10], _RANDOM[3'h5][9:0]};
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign responseIO_valid = responseIO_valid_0;
  assign responseIO_bits_tag = responseIO_bits_tag_0;
  assign responseIO_bits_data = responseIO_bits_data_0;
endmodule

