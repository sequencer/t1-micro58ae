module MaskUnitReadCrossBar(
  output       input_0_ready,
  input        input_0_valid,
  input  [4:0] input_0_bits_vs,
  input        input_0_bits_offset,
  input  [4:0] input_0_bits_readLane,
  input  [1:0] input_0_bits_dataOffset,
  output       input_1_ready,
  input        input_1_valid,
  input  [4:0] input_1_bits_vs,
  input        input_1_bits_offset,
  input  [4:0] input_1_bits_readLane,
  input  [1:0] input_1_bits_dataOffset,
  output       input_2_ready,
  input        input_2_valid,
  input  [4:0] input_2_bits_vs,
  input        input_2_bits_offset,
  input  [4:0] input_2_bits_readLane,
  input  [1:0] input_2_bits_dataOffset,
  output       input_3_ready,
  input        input_3_valid,
  input  [4:0] input_3_bits_vs,
  input        input_3_bits_offset,
  input  [4:0] input_3_bits_readLane,
  input  [1:0] input_3_bits_dataOffset,
  output       input_4_ready,
  input        input_4_valid,
  input  [4:0] input_4_bits_vs,
  input        input_4_bits_offset,
  input  [4:0] input_4_bits_readLane,
  input  [1:0] input_4_bits_dataOffset,
  output       input_5_ready,
  input        input_5_valid,
  input  [4:0] input_5_bits_vs,
  input        input_5_bits_offset,
  input  [4:0] input_5_bits_readLane,
  input  [1:0] input_5_bits_dataOffset,
  output       input_6_ready,
  input        input_6_valid,
  input  [4:0] input_6_bits_vs,
  input        input_6_bits_offset,
  input  [4:0] input_6_bits_readLane,
  input  [1:0] input_6_bits_dataOffset,
  output       input_7_ready,
  input        input_7_valid,
  input  [4:0] input_7_bits_vs,
  input        input_7_bits_offset,
  input  [4:0] input_7_bits_readLane,
  input  [1:0] input_7_bits_dataOffset,
  output       input_8_ready,
  input        input_8_valid,
  input  [4:0] input_8_bits_vs,
  input        input_8_bits_offset,
  input  [4:0] input_8_bits_readLane,
  input  [1:0] input_8_bits_dataOffset,
  output       input_9_ready,
  input        input_9_valid,
  input  [4:0] input_9_bits_vs,
  input        input_9_bits_offset,
  input  [4:0] input_9_bits_readLane,
  input  [1:0] input_9_bits_dataOffset,
  output       input_10_ready,
  input        input_10_valid,
  input  [4:0] input_10_bits_vs,
  input        input_10_bits_offset,
  input  [4:0] input_10_bits_readLane,
  input  [1:0] input_10_bits_dataOffset,
  output       input_11_ready,
  input        input_11_valid,
  input  [4:0] input_11_bits_vs,
  input        input_11_bits_offset,
  input  [4:0] input_11_bits_readLane,
  input  [1:0] input_11_bits_dataOffset,
  output       input_12_ready,
  input        input_12_valid,
  input  [4:0] input_12_bits_vs,
  input        input_12_bits_offset,
  input  [4:0] input_12_bits_readLane,
  input  [1:0] input_12_bits_dataOffset,
  output       input_13_ready,
  input        input_13_valid,
  input  [4:0] input_13_bits_vs,
  input        input_13_bits_offset,
  input  [4:0] input_13_bits_readLane,
  input  [1:0] input_13_bits_dataOffset,
  output       input_14_ready,
  input        input_14_valid,
  input  [4:0] input_14_bits_vs,
  input        input_14_bits_offset,
  input  [4:0] input_14_bits_readLane,
  input  [1:0] input_14_bits_dataOffset,
  output       input_15_ready,
  input        input_15_valid,
  input  [4:0] input_15_bits_vs,
  input        input_15_bits_offset,
  input  [4:0] input_15_bits_readLane,
  input  [1:0] input_15_bits_dataOffset,
  output       input_16_ready,
  input        input_16_valid,
  input  [4:0] input_16_bits_vs,
  input        input_16_bits_offset,
  input  [4:0] input_16_bits_readLane,
  input  [1:0] input_16_bits_dataOffset,
  output       input_17_ready,
  input        input_17_valid,
  input  [4:0] input_17_bits_vs,
  input        input_17_bits_offset,
  input  [4:0] input_17_bits_readLane,
  input  [1:0] input_17_bits_dataOffset,
  output       input_18_ready,
  input        input_18_valid,
  input  [4:0] input_18_bits_vs,
  input        input_18_bits_offset,
  input  [4:0] input_18_bits_readLane,
  input  [1:0] input_18_bits_dataOffset,
  output       input_19_ready,
  input        input_19_valid,
  input  [4:0] input_19_bits_vs,
  input        input_19_bits_offset,
  input  [4:0] input_19_bits_readLane,
  input  [1:0] input_19_bits_dataOffset,
  output       input_20_ready,
  input        input_20_valid,
  input  [4:0] input_20_bits_vs,
  input        input_20_bits_offset,
  input  [4:0] input_20_bits_readLane,
  input  [1:0] input_20_bits_dataOffset,
  output       input_21_ready,
  input        input_21_valid,
  input  [4:0] input_21_bits_vs,
  input        input_21_bits_offset,
  input  [4:0] input_21_bits_readLane,
  input  [1:0] input_21_bits_dataOffset,
  output       input_22_ready,
  input        input_22_valid,
  input  [4:0] input_22_bits_vs,
  input        input_22_bits_offset,
  input  [4:0] input_22_bits_readLane,
  input  [1:0] input_22_bits_dataOffset,
  output       input_23_ready,
  input        input_23_valid,
  input  [4:0] input_23_bits_vs,
  input        input_23_bits_offset,
  input  [4:0] input_23_bits_readLane,
  input  [1:0] input_23_bits_dataOffset,
  output       input_24_ready,
  input        input_24_valid,
  input  [4:0] input_24_bits_vs,
  input        input_24_bits_offset,
  input  [4:0] input_24_bits_readLane,
  input  [1:0] input_24_bits_dataOffset,
  output       input_25_ready,
  input        input_25_valid,
  input  [4:0] input_25_bits_vs,
  input        input_25_bits_offset,
  input  [4:0] input_25_bits_readLane,
  input  [1:0] input_25_bits_dataOffset,
  output       input_26_ready,
  input        input_26_valid,
  input  [4:0] input_26_bits_vs,
  input        input_26_bits_offset,
  input  [4:0] input_26_bits_readLane,
  input  [1:0] input_26_bits_dataOffset,
  output       input_27_ready,
  input        input_27_valid,
  input  [4:0] input_27_bits_vs,
  input        input_27_bits_offset,
  input  [4:0] input_27_bits_readLane,
  input  [1:0] input_27_bits_dataOffset,
  output       input_28_ready,
  input        input_28_valid,
  input  [4:0] input_28_bits_vs,
  input        input_28_bits_offset,
  input  [4:0] input_28_bits_readLane,
  input  [1:0] input_28_bits_dataOffset,
  output       input_29_ready,
  input        input_29_valid,
  input  [4:0] input_29_bits_vs,
  input        input_29_bits_offset,
  input  [4:0] input_29_bits_readLane,
  input  [1:0] input_29_bits_dataOffset,
  output       input_30_ready,
  input        input_30_valid,
  input  [4:0] input_30_bits_vs,
  input        input_30_bits_offset,
  input  [4:0] input_30_bits_readLane,
  input  [1:0] input_30_bits_dataOffset,
  output       input_31_ready,
  input        input_31_valid,
  input  [4:0] input_31_bits_vs,
  input        input_31_bits_offset,
  input  [4:0] input_31_bits_readLane,
  input  [1:0] input_31_bits_dataOffset,
  input        output_0_ready,
  output       output_0_valid,
  output [4:0] output_0_bits_vs,
  output       output_0_bits_offset,
  output [4:0] output_0_bits_writeIndex,
  output [1:0] output_0_bits_dataOffset,
  input        output_1_ready,
  output       output_1_valid,
  output [4:0] output_1_bits_vs,
  output       output_1_bits_offset,
  output [4:0] output_1_bits_writeIndex,
  output [1:0] output_1_bits_dataOffset,
  input        output_2_ready,
  output       output_2_valid,
  output [4:0] output_2_bits_vs,
  output       output_2_bits_offset,
  output [4:0] output_2_bits_writeIndex,
  output [1:0] output_2_bits_dataOffset,
  input        output_3_ready,
  output       output_3_valid,
  output [4:0] output_3_bits_vs,
  output       output_3_bits_offset,
  output [4:0] output_3_bits_writeIndex,
  output [1:0] output_3_bits_dataOffset,
  input        output_4_ready,
  output       output_4_valid,
  output [4:0] output_4_bits_vs,
  output       output_4_bits_offset,
  output [4:0] output_4_bits_writeIndex,
  output [1:0] output_4_bits_dataOffset,
  input        output_5_ready,
  output       output_5_valid,
  output [4:0] output_5_bits_vs,
  output       output_5_bits_offset,
  output [4:0] output_5_bits_writeIndex,
  output [1:0] output_5_bits_dataOffset,
  input        output_6_ready,
  output       output_6_valid,
  output [4:0] output_6_bits_vs,
  output       output_6_bits_offset,
  output [4:0] output_6_bits_writeIndex,
  output [1:0] output_6_bits_dataOffset,
  input        output_7_ready,
  output       output_7_valid,
  output [4:0] output_7_bits_vs,
  output       output_7_bits_offset,
  output [4:0] output_7_bits_writeIndex,
  output [1:0] output_7_bits_dataOffset,
  input        output_8_ready,
  output       output_8_valid,
  output [4:0] output_8_bits_vs,
  output       output_8_bits_offset,
  output [4:0] output_8_bits_writeIndex,
  output [1:0] output_8_bits_dataOffset,
  input        output_9_ready,
  output       output_9_valid,
  output [4:0] output_9_bits_vs,
  output       output_9_bits_offset,
  output [4:0] output_9_bits_writeIndex,
  output [1:0] output_9_bits_dataOffset,
  input        output_10_ready,
  output       output_10_valid,
  output [4:0] output_10_bits_vs,
  output       output_10_bits_offset,
  output [4:0] output_10_bits_writeIndex,
  output [1:0] output_10_bits_dataOffset,
  input        output_11_ready,
  output       output_11_valid,
  output [4:0] output_11_bits_vs,
  output       output_11_bits_offset,
  output [4:0] output_11_bits_writeIndex,
  output [1:0] output_11_bits_dataOffset,
  input        output_12_ready,
  output       output_12_valid,
  output [4:0] output_12_bits_vs,
  output       output_12_bits_offset,
  output [4:0] output_12_bits_writeIndex,
  output [1:0] output_12_bits_dataOffset,
  input        output_13_ready,
  output       output_13_valid,
  output [4:0] output_13_bits_vs,
  output       output_13_bits_offset,
  output [4:0] output_13_bits_writeIndex,
  output [1:0] output_13_bits_dataOffset,
  input        output_14_ready,
  output       output_14_valid,
  output [4:0] output_14_bits_vs,
  output       output_14_bits_offset,
  output [4:0] output_14_bits_writeIndex,
  output [1:0] output_14_bits_dataOffset,
  input        output_15_ready,
  output       output_15_valid,
  output [4:0] output_15_bits_vs,
  output       output_15_bits_offset,
  output [4:0] output_15_bits_writeIndex,
  output [1:0] output_15_bits_dataOffset,
  input        output_16_ready,
  output       output_16_valid,
  output [4:0] output_16_bits_vs,
  output       output_16_bits_offset,
  output [4:0] output_16_bits_writeIndex,
  output [1:0] output_16_bits_dataOffset,
  input        output_17_ready,
  output       output_17_valid,
  output [4:0] output_17_bits_vs,
  output       output_17_bits_offset,
  output [4:0] output_17_bits_writeIndex,
  output [1:0] output_17_bits_dataOffset,
  input        output_18_ready,
  output       output_18_valid,
  output [4:0] output_18_bits_vs,
  output       output_18_bits_offset,
  output [4:0] output_18_bits_writeIndex,
  output [1:0] output_18_bits_dataOffset,
  input        output_19_ready,
  output       output_19_valid,
  output [4:0] output_19_bits_vs,
  output       output_19_bits_offset,
  output [4:0] output_19_bits_writeIndex,
  output [1:0] output_19_bits_dataOffset,
  input        output_20_ready,
  output       output_20_valid,
  output [4:0] output_20_bits_vs,
  output       output_20_bits_offset,
  output [4:0] output_20_bits_writeIndex,
  output [1:0] output_20_bits_dataOffset,
  input        output_21_ready,
  output       output_21_valid,
  output [4:0] output_21_bits_vs,
  output       output_21_bits_offset,
  output [4:0] output_21_bits_writeIndex,
  output [1:0] output_21_bits_dataOffset,
  input        output_22_ready,
  output       output_22_valid,
  output [4:0] output_22_bits_vs,
  output       output_22_bits_offset,
  output [4:0] output_22_bits_writeIndex,
  output [1:0] output_22_bits_dataOffset,
  input        output_23_ready,
  output       output_23_valid,
  output [4:0] output_23_bits_vs,
  output       output_23_bits_offset,
  output [4:0] output_23_bits_writeIndex,
  output [1:0] output_23_bits_dataOffset,
  input        output_24_ready,
  output       output_24_valid,
  output [4:0] output_24_bits_vs,
  output       output_24_bits_offset,
  output [4:0] output_24_bits_writeIndex,
  output [1:0] output_24_bits_dataOffset,
  input        output_25_ready,
  output       output_25_valid,
  output [4:0] output_25_bits_vs,
  output       output_25_bits_offset,
  output [4:0] output_25_bits_writeIndex,
  output [1:0] output_25_bits_dataOffset,
  input        output_26_ready,
  output       output_26_valid,
  output [4:0] output_26_bits_vs,
  output       output_26_bits_offset,
  output [4:0] output_26_bits_writeIndex,
  output [1:0] output_26_bits_dataOffset,
  input        output_27_ready,
  output       output_27_valid,
  output [4:0] output_27_bits_vs,
  output       output_27_bits_offset,
  output [4:0] output_27_bits_writeIndex,
  output [1:0] output_27_bits_dataOffset,
  input        output_28_ready,
  output       output_28_valid,
  output [4:0] output_28_bits_vs,
  output       output_28_bits_offset,
  output [4:0] output_28_bits_writeIndex,
  output [1:0] output_28_bits_dataOffset,
  input        output_29_ready,
  output       output_29_valid,
  output [4:0] output_29_bits_vs,
  output       output_29_bits_offset,
  output [4:0] output_29_bits_writeIndex,
  output [1:0] output_29_bits_dataOffset,
  input        output_30_ready,
  output       output_30_valid,
  output [4:0] output_30_bits_vs,
  output       output_30_bits_offset,
  output [4:0] output_30_bits_writeIndex,
  output [1:0] output_30_bits_dataOffset,
  input        output_31_ready,
  output       output_31_valid,
  output [4:0] output_31_bits_vs,
  output       output_31_bits_offset,
  output [4:0] output_31_bits_writeIndex,
  output [1:0] output_31_bits_dataOffset
);

  wire        input_0_valid_0 = input_0_valid;
  wire [4:0]  input_0_bits_vs_0 = input_0_bits_vs;
  wire        input_0_bits_offset_0 = input_0_bits_offset;
  wire [4:0]  input_0_bits_readLane_0 = input_0_bits_readLane;
  wire [1:0]  input_0_bits_dataOffset_0 = input_0_bits_dataOffset;
  wire        input_1_valid_0 = input_1_valid;
  wire [4:0]  input_1_bits_vs_0 = input_1_bits_vs;
  wire        input_1_bits_offset_0 = input_1_bits_offset;
  wire [4:0]  input_1_bits_readLane_0 = input_1_bits_readLane;
  wire [1:0]  input_1_bits_dataOffset_0 = input_1_bits_dataOffset;
  wire        input_2_valid_0 = input_2_valid;
  wire [4:0]  input_2_bits_vs_0 = input_2_bits_vs;
  wire        input_2_bits_offset_0 = input_2_bits_offset;
  wire [4:0]  input_2_bits_readLane_0 = input_2_bits_readLane;
  wire [1:0]  input_2_bits_dataOffset_0 = input_2_bits_dataOffset;
  wire        input_3_valid_0 = input_3_valid;
  wire [4:0]  input_3_bits_vs_0 = input_3_bits_vs;
  wire        input_3_bits_offset_0 = input_3_bits_offset;
  wire [4:0]  input_3_bits_readLane_0 = input_3_bits_readLane;
  wire [1:0]  input_3_bits_dataOffset_0 = input_3_bits_dataOffset;
  wire        input_4_valid_0 = input_4_valid;
  wire [4:0]  input_4_bits_vs_0 = input_4_bits_vs;
  wire        input_4_bits_offset_0 = input_4_bits_offset;
  wire [4:0]  input_4_bits_readLane_0 = input_4_bits_readLane;
  wire [1:0]  input_4_bits_dataOffset_0 = input_4_bits_dataOffset;
  wire        input_5_valid_0 = input_5_valid;
  wire [4:0]  input_5_bits_vs_0 = input_5_bits_vs;
  wire        input_5_bits_offset_0 = input_5_bits_offset;
  wire [4:0]  input_5_bits_readLane_0 = input_5_bits_readLane;
  wire [1:0]  input_5_bits_dataOffset_0 = input_5_bits_dataOffset;
  wire        input_6_valid_0 = input_6_valid;
  wire [4:0]  input_6_bits_vs_0 = input_6_bits_vs;
  wire        input_6_bits_offset_0 = input_6_bits_offset;
  wire [4:0]  input_6_bits_readLane_0 = input_6_bits_readLane;
  wire [1:0]  input_6_bits_dataOffset_0 = input_6_bits_dataOffset;
  wire        input_7_valid_0 = input_7_valid;
  wire [4:0]  input_7_bits_vs_0 = input_7_bits_vs;
  wire        input_7_bits_offset_0 = input_7_bits_offset;
  wire [4:0]  input_7_bits_readLane_0 = input_7_bits_readLane;
  wire [1:0]  input_7_bits_dataOffset_0 = input_7_bits_dataOffset;
  wire        input_8_valid_0 = input_8_valid;
  wire [4:0]  input_8_bits_vs_0 = input_8_bits_vs;
  wire        input_8_bits_offset_0 = input_8_bits_offset;
  wire [4:0]  input_8_bits_readLane_0 = input_8_bits_readLane;
  wire [1:0]  input_8_bits_dataOffset_0 = input_8_bits_dataOffset;
  wire        input_9_valid_0 = input_9_valid;
  wire [4:0]  input_9_bits_vs_0 = input_9_bits_vs;
  wire        input_9_bits_offset_0 = input_9_bits_offset;
  wire [4:0]  input_9_bits_readLane_0 = input_9_bits_readLane;
  wire [1:0]  input_9_bits_dataOffset_0 = input_9_bits_dataOffset;
  wire        input_10_valid_0 = input_10_valid;
  wire [4:0]  input_10_bits_vs_0 = input_10_bits_vs;
  wire        input_10_bits_offset_0 = input_10_bits_offset;
  wire [4:0]  input_10_bits_readLane_0 = input_10_bits_readLane;
  wire [1:0]  input_10_bits_dataOffset_0 = input_10_bits_dataOffset;
  wire        input_11_valid_0 = input_11_valid;
  wire [4:0]  input_11_bits_vs_0 = input_11_bits_vs;
  wire        input_11_bits_offset_0 = input_11_bits_offset;
  wire [4:0]  input_11_bits_readLane_0 = input_11_bits_readLane;
  wire [1:0]  input_11_bits_dataOffset_0 = input_11_bits_dataOffset;
  wire        input_12_valid_0 = input_12_valid;
  wire [4:0]  input_12_bits_vs_0 = input_12_bits_vs;
  wire        input_12_bits_offset_0 = input_12_bits_offset;
  wire [4:0]  input_12_bits_readLane_0 = input_12_bits_readLane;
  wire [1:0]  input_12_bits_dataOffset_0 = input_12_bits_dataOffset;
  wire        input_13_valid_0 = input_13_valid;
  wire [4:0]  input_13_bits_vs_0 = input_13_bits_vs;
  wire        input_13_bits_offset_0 = input_13_bits_offset;
  wire [4:0]  input_13_bits_readLane_0 = input_13_bits_readLane;
  wire [1:0]  input_13_bits_dataOffset_0 = input_13_bits_dataOffset;
  wire        input_14_valid_0 = input_14_valid;
  wire [4:0]  input_14_bits_vs_0 = input_14_bits_vs;
  wire        input_14_bits_offset_0 = input_14_bits_offset;
  wire [4:0]  input_14_bits_readLane_0 = input_14_bits_readLane;
  wire [1:0]  input_14_bits_dataOffset_0 = input_14_bits_dataOffset;
  wire        input_15_valid_0 = input_15_valid;
  wire [4:0]  input_15_bits_vs_0 = input_15_bits_vs;
  wire        input_15_bits_offset_0 = input_15_bits_offset;
  wire [4:0]  input_15_bits_readLane_0 = input_15_bits_readLane;
  wire [1:0]  input_15_bits_dataOffset_0 = input_15_bits_dataOffset;
  wire        input_16_valid_0 = input_16_valid;
  wire [4:0]  input_16_bits_vs_0 = input_16_bits_vs;
  wire        input_16_bits_offset_0 = input_16_bits_offset;
  wire [4:0]  input_16_bits_readLane_0 = input_16_bits_readLane;
  wire [1:0]  input_16_bits_dataOffset_0 = input_16_bits_dataOffset;
  wire        input_17_valid_0 = input_17_valid;
  wire [4:0]  input_17_bits_vs_0 = input_17_bits_vs;
  wire        input_17_bits_offset_0 = input_17_bits_offset;
  wire [4:0]  input_17_bits_readLane_0 = input_17_bits_readLane;
  wire [1:0]  input_17_bits_dataOffset_0 = input_17_bits_dataOffset;
  wire        input_18_valid_0 = input_18_valid;
  wire [4:0]  input_18_bits_vs_0 = input_18_bits_vs;
  wire        input_18_bits_offset_0 = input_18_bits_offset;
  wire [4:0]  input_18_bits_readLane_0 = input_18_bits_readLane;
  wire [1:0]  input_18_bits_dataOffset_0 = input_18_bits_dataOffset;
  wire        input_19_valid_0 = input_19_valid;
  wire [4:0]  input_19_bits_vs_0 = input_19_bits_vs;
  wire        input_19_bits_offset_0 = input_19_bits_offset;
  wire [4:0]  input_19_bits_readLane_0 = input_19_bits_readLane;
  wire [1:0]  input_19_bits_dataOffset_0 = input_19_bits_dataOffset;
  wire        input_20_valid_0 = input_20_valid;
  wire [4:0]  input_20_bits_vs_0 = input_20_bits_vs;
  wire        input_20_bits_offset_0 = input_20_bits_offset;
  wire [4:0]  input_20_bits_readLane_0 = input_20_bits_readLane;
  wire [1:0]  input_20_bits_dataOffset_0 = input_20_bits_dataOffset;
  wire        input_21_valid_0 = input_21_valid;
  wire [4:0]  input_21_bits_vs_0 = input_21_bits_vs;
  wire        input_21_bits_offset_0 = input_21_bits_offset;
  wire [4:0]  input_21_bits_readLane_0 = input_21_bits_readLane;
  wire [1:0]  input_21_bits_dataOffset_0 = input_21_bits_dataOffset;
  wire        input_22_valid_0 = input_22_valid;
  wire [4:0]  input_22_bits_vs_0 = input_22_bits_vs;
  wire        input_22_bits_offset_0 = input_22_bits_offset;
  wire [4:0]  input_22_bits_readLane_0 = input_22_bits_readLane;
  wire [1:0]  input_22_bits_dataOffset_0 = input_22_bits_dataOffset;
  wire        input_23_valid_0 = input_23_valid;
  wire [4:0]  input_23_bits_vs_0 = input_23_bits_vs;
  wire        input_23_bits_offset_0 = input_23_bits_offset;
  wire [4:0]  input_23_bits_readLane_0 = input_23_bits_readLane;
  wire [1:0]  input_23_bits_dataOffset_0 = input_23_bits_dataOffset;
  wire        input_24_valid_0 = input_24_valid;
  wire [4:0]  input_24_bits_vs_0 = input_24_bits_vs;
  wire        input_24_bits_offset_0 = input_24_bits_offset;
  wire [4:0]  input_24_bits_readLane_0 = input_24_bits_readLane;
  wire [1:0]  input_24_bits_dataOffset_0 = input_24_bits_dataOffset;
  wire        input_25_valid_0 = input_25_valid;
  wire [4:0]  input_25_bits_vs_0 = input_25_bits_vs;
  wire        input_25_bits_offset_0 = input_25_bits_offset;
  wire [4:0]  input_25_bits_readLane_0 = input_25_bits_readLane;
  wire [1:0]  input_25_bits_dataOffset_0 = input_25_bits_dataOffset;
  wire        input_26_valid_0 = input_26_valid;
  wire [4:0]  input_26_bits_vs_0 = input_26_bits_vs;
  wire        input_26_bits_offset_0 = input_26_bits_offset;
  wire [4:0]  input_26_bits_readLane_0 = input_26_bits_readLane;
  wire [1:0]  input_26_bits_dataOffset_0 = input_26_bits_dataOffset;
  wire        input_27_valid_0 = input_27_valid;
  wire [4:0]  input_27_bits_vs_0 = input_27_bits_vs;
  wire        input_27_bits_offset_0 = input_27_bits_offset;
  wire [4:0]  input_27_bits_readLane_0 = input_27_bits_readLane;
  wire [1:0]  input_27_bits_dataOffset_0 = input_27_bits_dataOffset;
  wire        input_28_valid_0 = input_28_valid;
  wire [4:0]  input_28_bits_vs_0 = input_28_bits_vs;
  wire        input_28_bits_offset_0 = input_28_bits_offset;
  wire [4:0]  input_28_bits_readLane_0 = input_28_bits_readLane;
  wire [1:0]  input_28_bits_dataOffset_0 = input_28_bits_dataOffset;
  wire        input_29_valid_0 = input_29_valid;
  wire [4:0]  input_29_bits_vs_0 = input_29_bits_vs;
  wire        input_29_bits_offset_0 = input_29_bits_offset;
  wire [4:0]  input_29_bits_readLane_0 = input_29_bits_readLane;
  wire [1:0]  input_29_bits_dataOffset_0 = input_29_bits_dataOffset;
  wire        input_30_valid_0 = input_30_valid;
  wire [4:0]  input_30_bits_vs_0 = input_30_bits_vs;
  wire        input_30_bits_offset_0 = input_30_bits_offset;
  wire [4:0]  input_30_bits_readLane_0 = input_30_bits_readLane;
  wire [1:0]  input_30_bits_dataOffset_0 = input_30_bits_dataOffset;
  wire        input_31_valid_0 = input_31_valid;
  wire [4:0]  input_31_bits_vs_0 = input_31_bits_vs;
  wire        input_31_bits_offset_0 = input_31_bits_offset;
  wire [4:0]  input_31_bits_readLane_0 = input_31_bits_readLane;
  wire [1:0]  input_31_bits_dataOffset_0 = input_31_bits_dataOffset;
  wire        output_0_ready_0 = output_0_ready;
  wire        output_1_ready_0 = output_1_ready;
  wire        output_2_ready_0 = output_2_ready;
  wire        output_3_ready_0 = output_3_ready;
  wire        output_4_ready_0 = output_4_ready;
  wire        output_5_ready_0 = output_5_ready;
  wire        output_6_ready_0 = output_6_ready;
  wire        output_7_ready_0 = output_7_ready;
  wire        output_8_ready_0 = output_8_ready;
  wire        output_9_ready_0 = output_9_ready;
  wire        output_10_ready_0 = output_10_ready;
  wire        output_11_ready_0 = output_11_ready;
  wire        output_12_ready_0 = output_12_ready;
  wire        output_13_ready_0 = output_13_ready;
  wire        output_14_ready_0 = output_14_ready;
  wire        output_15_ready_0 = output_15_ready;
  wire        output_16_ready_0 = output_16_ready;
  wire        output_17_ready_0 = output_17_ready;
  wire        output_18_ready_0 = output_18_ready;
  wire        output_19_ready_0 = output_19_ready;
  wire        output_20_ready_0 = output_20_ready;
  wire        output_21_ready_0 = output_21_ready;
  wire        output_22_ready_0 = output_22_ready;
  wire        output_23_ready_0 = output_23_ready;
  wire        output_24_ready_0 = output_24_ready;
  wire        output_25_ready_0 = output_25_ready;
  wire        output_26_ready_0 = output_26_ready;
  wire        output_27_ready_0 = output_27_ready;
  wire        output_28_ready_0 = output_28_ready;
  wire        output_29_ready_0 = output_29_ready;
  wire        output_30_ready_0 = output_30_ready;
  wire        output_31_ready_0 = output_31_ready;
  wire [4:0]  input_31_bits_requestIndex = 5'h1F;
  wire [4:0]  input_30_bits_requestIndex = 5'h1E;
  wire [4:0]  input_29_bits_requestIndex = 5'h1D;
  wire [4:0]  input_28_bits_requestIndex = 5'h1C;
  wire [4:0]  input_27_bits_requestIndex = 5'h1B;
  wire [4:0]  input_26_bits_requestIndex = 5'h1A;
  wire [4:0]  input_25_bits_requestIndex = 5'h19;
  wire [4:0]  input_24_bits_requestIndex = 5'h18;
  wire [4:0]  input_23_bits_requestIndex = 5'h17;
  wire [4:0]  input_22_bits_requestIndex = 5'h16;
  wire [4:0]  input_21_bits_requestIndex = 5'h15;
  wire [4:0]  input_20_bits_requestIndex = 5'h14;
  wire [4:0]  input_19_bits_requestIndex = 5'h13;
  wire [4:0]  input_18_bits_requestIndex = 5'h12;
  wire [4:0]  input_17_bits_requestIndex = 5'h11;
  wire [4:0]  input_16_bits_requestIndex = 5'h10;
  wire [4:0]  input_15_bits_requestIndex = 5'hF;
  wire [4:0]  input_14_bits_requestIndex = 5'hE;
  wire [4:0]  input_13_bits_requestIndex = 5'hD;
  wire [4:0]  input_12_bits_requestIndex = 5'hC;
  wire [4:0]  input_11_bits_requestIndex = 5'hB;
  wire [4:0]  input_10_bits_requestIndex = 5'hA;
  wire [4:0]  input_9_bits_requestIndex = 5'h9;
  wire [4:0]  input_8_bits_requestIndex = 5'h8;
  wire [4:0]  input_7_bits_requestIndex = 5'h7;
  wire [4:0]  input_6_bits_requestIndex = 5'h6;
  wire [4:0]  input_5_bits_requestIndex = 5'h5;
  wire [4:0]  input_4_bits_requestIndex = 5'h4;
  wire [4:0]  input_3_bits_requestIndex = 5'h3;
  wire [4:0]  input_2_bits_requestIndex = 5'h2;
  wire [4:0]  input_1_bits_requestIndex = 5'h1;
  wire [4:0]  input_0_bits_requestIndex = 5'h0;
  wire [4:0]  selectReq_bits_vs;
  wire        selectReq_bits_offset;
  wire [4:0]  selectReq_bits_requestIndex;
  wire [1:0]  selectReq_bits_dataOffset;
  wire [4:0]  selectReq_1_bits_vs;
  wire        selectReq_1_bits_offset;
  wire [4:0]  selectReq_1_bits_requestIndex;
  wire [1:0]  selectReq_1_bits_dataOffset;
  wire [4:0]  selectReq_2_bits_vs;
  wire        selectReq_2_bits_offset;
  wire [4:0]  selectReq_2_bits_requestIndex;
  wire [1:0]  selectReq_2_bits_dataOffset;
  wire [4:0]  selectReq_3_bits_vs;
  wire        selectReq_3_bits_offset;
  wire [4:0]  selectReq_3_bits_requestIndex;
  wire [1:0]  selectReq_3_bits_dataOffset;
  wire [4:0]  selectReq_4_bits_vs;
  wire        selectReq_4_bits_offset;
  wire [4:0]  selectReq_4_bits_requestIndex;
  wire [1:0]  selectReq_4_bits_dataOffset;
  wire [4:0]  selectReq_5_bits_vs;
  wire        selectReq_5_bits_offset;
  wire [4:0]  selectReq_5_bits_requestIndex;
  wire [1:0]  selectReq_5_bits_dataOffset;
  wire [4:0]  selectReq_6_bits_vs;
  wire        selectReq_6_bits_offset;
  wire [4:0]  selectReq_6_bits_requestIndex;
  wire [1:0]  selectReq_6_bits_dataOffset;
  wire [4:0]  selectReq_7_bits_vs;
  wire        selectReq_7_bits_offset;
  wire [4:0]  selectReq_7_bits_requestIndex;
  wire [1:0]  selectReq_7_bits_dataOffset;
  wire [4:0]  selectReq_8_bits_vs;
  wire        selectReq_8_bits_offset;
  wire [4:0]  selectReq_8_bits_requestIndex;
  wire [1:0]  selectReq_8_bits_dataOffset;
  wire [4:0]  selectReq_9_bits_vs;
  wire        selectReq_9_bits_offset;
  wire [4:0]  selectReq_9_bits_requestIndex;
  wire [1:0]  selectReq_9_bits_dataOffset;
  wire [4:0]  selectReq_10_bits_vs;
  wire        selectReq_10_bits_offset;
  wire [4:0]  selectReq_10_bits_requestIndex;
  wire [1:0]  selectReq_10_bits_dataOffset;
  wire [4:0]  selectReq_11_bits_vs;
  wire        selectReq_11_bits_offset;
  wire [4:0]  selectReq_11_bits_requestIndex;
  wire [1:0]  selectReq_11_bits_dataOffset;
  wire [4:0]  selectReq_12_bits_vs;
  wire        selectReq_12_bits_offset;
  wire [4:0]  selectReq_12_bits_requestIndex;
  wire [1:0]  selectReq_12_bits_dataOffset;
  wire [4:0]  selectReq_13_bits_vs;
  wire        selectReq_13_bits_offset;
  wire [4:0]  selectReq_13_bits_requestIndex;
  wire [1:0]  selectReq_13_bits_dataOffset;
  wire [4:0]  selectReq_14_bits_vs;
  wire        selectReq_14_bits_offset;
  wire [4:0]  selectReq_14_bits_requestIndex;
  wire [1:0]  selectReq_14_bits_dataOffset;
  wire [4:0]  selectReq_15_bits_vs;
  wire        selectReq_15_bits_offset;
  wire [4:0]  selectReq_15_bits_requestIndex;
  wire [1:0]  selectReq_15_bits_dataOffset;
  wire [4:0]  selectReq_16_bits_vs;
  wire        selectReq_16_bits_offset;
  wire [4:0]  selectReq_16_bits_requestIndex;
  wire [1:0]  selectReq_16_bits_dataOffset;
  wire [4:0]  selectReq_17_bits_vs;
  wire        selectReq_17_bits_offset;
  wire [4:0]  selectReq_17_bits_requestIndex;
  wire [1:0]  selectReq_17_bits_dataOffset;
  wire [4:0]  selectReq_18_bits_vs;
  wire        selectReq_18_bits_offset;
  wire [4:0]  selectReq_18_bits_requestIndex;
  wire [1:0]  selectReq_18_bits_dataOffset;
  wire [4:0]  selectReq_19_bits_vs;
  wire        selectReq_19_bits_offset;
  wire [4:0]  selectReq_19_bits_requestIndex;
  wire [1:0]  selectReq_19_bits_dataOffset;
  wire [4:0]  selectReq_20_bits_vs;
  wire        selectReq_20_bits_offset;
  wire [4:0]  selectReq_20_bits_requestIndex;
  wire [1:0]  selectReq_20_bits_dataOffset;
  wire [4:0]  selectReq_21_bits_vs;
  wire        selectReq_21_bits_offset;
  wire [4:0]  selectReq_21_bits_requestIndex;
  wire [1:0]  selectReq_21_bits_dataOffset;
  wire [4:0]  selectReq_22_bits_vs;
  wire        selectReq_22_bits_offset;
  wire [4:0]  selectReq_22_bits_requestIndex;
  wire [1:0]  selectReq_22_bits_dataOffset;
  wire [4:0]  selectReq_23_bits_vs;
  wire        selectReq_23_bits_offset;
  wire [4:0]  selectReq_23_bits_requestIndex;
  wire [1:0]  selectReq_23_bits_dataOffset;
  wire [4:0]  selectReq_24_bits_vs;
  wire        selectReq_24_bits_offset;
  wire [4:0]  selectReq_24_bits_requestIndex;
  wire [1:0]  selectReq_24_bits_dataOffset;
  wire [4:0]  selectReq_25_bits_vs;
  wire        selectReq_25_bits_offset;
  wire [4:0]  selectReq_25_bits_requestIndex;
  wire [1:0]  selectReq_25_bits_dataOffset;
  wire [4:0]  selectReq_26_bits_vs;
  wire        selectReq_26_bits_offset;
  wire [4:0]  selectReq_26_bits_requestIndex;
  wire [1:0]  selectReq_26_bits_dataOffset;
  wire [4:0]  selectReq_27_bits_vs;
  wire        selectReq_27_bits_offset;
  wire [4:0]  selectReq_27_bits_requestIndex;
  wire [1:0]  selectReq_27_bits_dataOffset;
  wire [4:0]  selectReq_28_bits_vs;
  wire        selectReq_28_bits_offset;
  wire [4:0]  selectReq_28_bits_requestIndex;
  wire [1:0]  selectReq_28_bits_dataOffset;
  wire [4:0]  selectReq_29_bits_vs;
  wire        selectReq_29_bits_offset;
  wire [4:0]  selectReq_29_bits_requestIndex;
  wire [1:0]  selectReq_29_bits_dataOffset;
  wire [4:0]  selectReq_30_bits_vs;
  wire        selectReq_30_bits_offset;
  wire [4:0]  selectReq_30_bits_requestIndex;
  wire [1:0]  selectReq_30_bits_dataOffset;
  wire [4:0]  selectReq_31_bits_vs;
  wire        selectReq_31_bits_offset;
  wire [4:0]  selectReq_31_bits_requestIndex;
  wire [1:0]  selectReq_31_bits_dataOffset;
  wire [31:0] requestReadLane = 32'h1 << input_0_bits_readLane_0;
  wire        free = |requestReadLane;
  wire        outReady =
    requestReadLane[0] & output_0_ready_0 | requestReadLane[1] & output_1_ready_0 | requestReadLane[2] & output_2_ready_0 | requestReadLane[3] & output_3_ready_0 | requestReadLane[4] & output_4_ready_0 | requestReadLane[5]
    & output_5_ready_0 | requestReadLane[6] & output_6_ready_0 | requestReadLane[7] & output_7_ready_0 | requestReadLane[8] & output_8_ready_0 | requestReadLane[9] & output_9_ready_0 | requestReadLane[10] & output_10_ready_0
    | requestReadLane[11] & output_11_ready_0 | requestReadLane[12] & output_12_ready_0 | requestReadLane[13] & output_13_ready_0 | requestReadLane[14] & output_14_ready_0 | requestReadLane[15] & output_15_ready_0 | requestReadLane[16]
    & output_16_ready_0 | requestReadLane[17] & output_17_ready_0 | requestReadLane[18] & output_18_ready_0 | requestReadLane[19] & output_19_ready_0 | requestReadLane[20] & output_20_ready_0 | requestReadLane[21] & output_21_ready_0
    | requestReadLane[22] & output_22_ready_0 | requestReadLane[23] & output_23_ready_0 | requestReadLane[24] & output_24_ready_0 | requestReadLane[25] & output_25_ready_0 | requestReadLane[26] & output_26_ready_0 | requestReadLane[27]
    & output_27_ready_0 | requestReadLane[28] & output_28_ready_0 | requestReadLane[29] & output_29_ready_0 | requestReadLane[30] & output_30_ready_0 | requestReadLane[31] & output_31_ready_0;
  wire        input_0_ready_0 = free & outReady;
  wire [31:0] inputSelect1H_0 = input_0_valid_0 & free ? requestReadLane : 32'h0;
  wire [31:0] requestReadLane_1 = 32'h1 << input_1_bits_readLane_0;
  wire        free_1 = |(requestReadLane_1 & ~inputSelect1H_0);
  wire        outReady_1 =
    requestReadLane_1[0] & output_0_ready_0 | requestReadLane_1[1] & output_1_ready_0 | requestReadLane_1[2] & output_2_ready_0 | requestReadLane_1[3] & output_3_ready_0 | requestReadLane_1[4] & output_4_ready_0 | requestReadLane_1[5]
    & output_5_ready_0 | requestReadLane_1[6] & output_6_ready_0 | requestReadLane_1[7] & output_7_ready_0 | requestReadLane_1[8] & output_8_ready_0 | requestReadLane_1[9] & output_9_ready_0 | requestReadLane_1[10] & output_10_ready_0
    | requestReadLane_1[11] & output_11_ready_0 | requestReadLane_1[12] & output_12_ready_0 | requestReadLane_1[13] & output_13_ready_0 | requestReadLane_1[14] & output_14_ready_0 | requestReadLane_1[15] & output_15_ready_0
    | requestReadLane_1[16] & output_16_ready_0 | requestReadLane_1[17] & output_17_ready_0 | requestReadLane_1[18] & output_18_ready_0 | requestReadLane_1[19] & output_19_ready_0 | requestReadLane_1[20] & output_20_ready_0
    | requestReadLane_1[21] & output_21_ready_0 | requestReadLane_1[22] & output_22_ready_0 | requestReadLane_1[23] & output_23_ready_0 | requestReadLane_1[24] & output_24_ready_0 | requestReadLane_1[25] & output_25_ready_0
    | requestReadLane_1[26] & output_26_ready_0 | requestReadLane_1[27] & output_27_ready_0 | requestReadLane_1[28] & output_28_ready_0 | requestReadLane_1[29] & output_29_ready_0 | requestReadLane_1[30] & output_30_ready_0
    | requestReadLane_1[31] & output_31_ready_0;
  wire        input_1_ready_0 = free_1 & outReady_1;
  wire [31:0] inputSelect1H_1 = input_1_valid_0 & free_1 ? requestReadLane_1 : 32'h0;
  wire [31:0] _GEN = inputSelect1H_0 | inputSelect1H_1;
  wire [31:0] requestReadLane_2 = 32'h1 << input_2_bits_readLane_0;
  wire        free_2 = |(requestReadLane_2 & ~_GEN);
  wire        outReady_2 =
    requestReadLane_2[0] & output_0_ready_0 | requestReadLane_2[1] & output_1_ready_0 | requestReadLane_2[2] & output_2_ready_0 | requestReadLane_2[3] & output_3_ready_0 | requestReadLane_2[4] & output_4_ready_0 | requestReadLane_2[5]
    & output_5_ready_0 | requestReadLane_2[6] & output_6_ready_0 | requestReadLane_2[7] & output_7_ready_0 | requestReadLane_2[8] & output_8_ready_0 | requestReadLane_2[9] & output_9_ready_0 | requestReadLane_2[10] & output_10_ready_0
    | requestReadLane_2[11] & output_11_ready_0 | requestReadLane_2[12] & output_12_ready_0 | requestReadLane_2[13] & output_13_ready_0 | requestReadLane_2[14] & output_14_ready_0 | requestReadLane_2[15] & output_15_ready_0
    | requestReadLane_2[16] & output_16_ready_0 | requestReadLane_2[17] & output_17_ready_0 | requestReadLane_2[18] & output_18_ready_0 | requestReadLane_2[19] & output_19_ready_0 | requestReadLane_2[20] & output_20_ready_0
    | requestReadLane_2[21] & output_21_ready_0 | requestReadLane_2[22] & output_22_ready_0 | requestReadLane_2[23] & output_23_ready_0 | requestReadLane_2[24] & output_24_ready_0 | requestReadLane_2[25] & output_25_ready_0
    | requestReadLane_2[26] & output_26_ready_0 | requestReadLane_2[27] & output_27_ready_0 | requestReadLane_2[28] & output_28_ready_0 | requestReadLane_2[29] & output_29_ready_0 | requestReadLane_2[30] & output_30_ready_0
    | requestReadLane_2[31] & output_31_ready_0;
  wire        input_2_ready_0 = free_2 & outReady_2;
  wire [31:0] inputSelect1H_2 = input_2_valid_0 & free_2 ? requestReadLane_2 : 32'h0;
  wire [31:0] _GEN_0 = _GEN | inputSelect1H_2;
  wire [31:0] requestReadLane_3 = 32'h1 << input_3_bits_readLane_0;
  wire        free_3 = |(requestReadLane_3 & ~_GEN_0);
  wire        outReady_3 =
    requestReadLane_3[0] & output_0_ready_0 | requestReadLane_3[1] & output_1_ready_0 | requestReadLane_3[2] & output_2_ready_0 | requestReadLane_3[3] & output_3_ready_0 | requestReadLane_3[4] & output_4_ready_0 | requestReadLane_3[5]
    & output_5_ready_0 | requestReadLane_3[6] & output_6_ready_0 | requestReadLane_3[7] & output_7_ready_0 | requestReadLane_3[8] & output_8_ready_0 | requestReadLane_3[9] & output_9_ready_0 | requestReadLane_3[10] & output_10_ready_0
    | requestReadLane_3[11] & output_11_ready_0 | requestReadLane_3[12] & output_12_ready_0 | requestReadLane_3[13] & output_13_ready_0 | requestReadLane_3[14] & output_14_ready_0 | requestReadLane_3[15] & output_15_ready_0
    | requestReadLane_3[16] & output_16_ready_0 | requestReadLane_3[17] & output_17_ready_0 | requestReadLane_3[18] & output_18_ready_0 | requestReadLane_3[19] & output_19_ready_0 | requestReadLane_3[20] & output_20_ready_0
    | requestReadLane_3[21] & output_21_ready_0 | requestReadLane_3[22] & output_22_ready_0 | requestReadLane_3[23] & output_23_ready_0 | requestReadLane_3[24] & output_24_ready_0 | requestReadLane_3[25] & output_25_ready_0
    | requestReadLane_3[26] & output_26_ready_0 | requestReadLane_3[27] & output_27_ready_0 | requestReadLane_3[28] & output_28_ready_0 | requestReadLane_3[29] & output_29_ready_0 | requestReadLane_3[30] & output_30_ready_0
    | requestReadLane_3[31] & output_31_ready_0;
  wire        input_3_ready_0 = free_3 & outReady_3;
  wire [31:0] inputSelect1H_3 = input_3_valid_0 & free_3 ? requestReadLane_3 : 32'h0;
  wire [31:0] _GEN_1 = _GEN_0 | inputSelect1H_3;
  wire [31:0] requestReadLane_4 = 32'h1 << input_4_bits_readLane_0;
  wire        free_4 = |(requestReadLane_4 & ~_GEN_1);
  wire        outReady_4 =
    requestReadLane_4[0] & output_0_ready_0 | requestReadLane_4[1] & output_1_ready_0 | requestReadLane_4[2] & output_2_ready_0 | requestReadLane_4[3] & output_3_ready_0 | requestReadLane_4[4] & output_4_ready_0 | requestReadLane_4[5]
    & output_5_ready_0 | requestReadLane_4[6] & output_6_ready_0 | requestReadLane_4[7] & output_7_ready_0 | requestReadLane_4[8] & output_8_ready_0 | requestReadLane_4[9] & output_9_ready_0 | requestReadLane_4[10] & output_10_ready_0
    | requestReadLane_4[11] & output_11_ready_0 | requestReadLane_4[12] & output_12_ready_0 | requestReadLane_4[13] & output_13_ready_0 | requestReadLane_4[14] & output_14_ready_0 | requestReadLane_4[15] & output_15_ready_0
    | requestReadLane_4[16] & output_16_ready_0 | requestReadLane_4[17] & output_17_ready_0 | requestReadLane_4[18] & output_18_ready_0 | requestReadLane_4[19] & output_19_ready_0 | requestReadLane_4[20] & output_20_ready_0
    | requestReadLane_4[21] & output_21_ready_0 | requestReadLane_4[22] & output_22_ready_0 | requestReadLane_4[23] & output_23_ready_0 | requestReadLane_4[24] & output_24_ready_0 | requestReadLane_4[25] & output_25_ready_0
    | requestReadLane_4[26] & output_26_ready_0 | requestReadLane_4[27] & output_27_ready_0 | requestReadLane_4[28] & output_28_ready_0 | requestReadLane_4[29] & output_29_ready_0 | requestReadLane_4[30] & output_30_ready_0
    | requestReadLane_4[31] & output_31_ready_0;
  wire        input_4_ready_0 = free_4 & outReady_4;
  wire [31:0] inputSelect1H_4 = input_4_valid_0 & free_4 ? requestReadLane_4 : 32'h0;
  wire [31:0] _GEN_2 = _GEN_1 | inputSelect1H_4;
  wire [31:0] requestReadLane_5 = 32'h1 << input_5_bits_readLane_0;
  wire        free_5 = |(requestReadLane_5 & ~_GEN_2);
  wire        outReady_5 =
    requestReadLane_5[0] & output_0_ready_0 | requestReadLane_5[1] & output_1_ready_0 | requestReadLane_5[2] & output_2_ready_0 | requestReadLane_5[3] & output_3_ready_0 | requestReadLane_5[4] & output_4_ready_0 | requestReadLane_5[5]
    & output_5_ready_0 | requestReadLane_5[6] & output_6_ready_0 | requestReadLane_5[7] & output_7_ready_0 | requestReadLane_5[8] & output_8_ready_0 | requestReadLane_5[9] & output_9_ready_0 | requestReadLane_5[10] & output_10_ready_0
    | requestReadLane_5[11] & output_11_ready_0 | requestReadLane_5[12] & output_12_ready_0 | requestReadLane_5[13] & output_13_ready_0 | requestReadLane_5[14] & output_14_ready_0 | requestReadLane_5[15] & output_15_ready_0
    | requestReadLane_5[16] & output_16_ready_0 | requestReadLane_5[17] & output_17_ready_0 | requestReadLane_5[18] & output_18_ready_0 | requestReadLane_5[19] & output_19_ready_0 | requestReadLane_5[20] & output_20_ready_0
    | requestReadLane_5[21] & output_21_ready_0 | requestReadLane_5[22] & output_22_ready_0 | requestReadLane_5[23] & output_23_ready_0 | requestReadLane_5[24] & output_24_ready_0 | requestReadLane_5[25] & output_25_ready_0
    | requestReadLane_5[26] & output_26_ready_0 | requestReadLane_5[27] & output_27_ready_0 | requestReadLane_5[28] & output_28_ready_0 | requestReadLane_5[29] & output_29_ready_0 | requestReadLane_5[30] & output_30_ready_0
    | requestReadLane_5[31] & output_31_ready_0;
  wire        input_5_ready_0 = free_5 & outReady_5;
  wire [31:0] inputSelect1H_5 = input_5_valid_0 & free_5 ? requestReadLane_5 : 32'h0;
  wire [31:0] _GEN_3 = _GEN_2 | inputSelect1H_5;
  wire [31:0] requestReadLane_6 = 32'h1 << input_6_bits_readLane_0;
  wire        free_6 = |(requestReadLane_6 & ~_GEN_3);
  wire        outReady_6 =
    requestReadLane_6[0] & output_0_ready_0 | requestReadLane_6[1] & output_1_ready_0 | requestReadLane_6[2] & output_2_ready_0 | requestReadLane_6[3] & output_3_ready_0 | requestReadLane_6[4] & output_4_ready_0 | requestReadLane_6[5]
    & output_5_ready_0 | requestReadLane_6[6] & output_6_ready_0 | requestReadLane_6[7] & output_7_ready_0 | requestReadLane_6[8] & output_8_ready_0 | requestReadLane_6[9] & output_9_ready_0 | requestReadLane_6[10] & output_10_ready_0
    | requestReadLane_6[11] & output_11_ready_0 | requestReadLane_6[12] & output_12_ready_0 | requestReadLane_6[13] & output_13_ready_0 | requestReadLane_6[14] & output_14_ready_0 | requestReadLane_6[15] & output_15_ready_0
    | requestReadLane_6[16] & output_16_ready_0 | requestReadLane_6[17] & output_17_ready_0 | requestReadLane_6[18] & output_18_ready_0 | requestReadLane_6[19] & output_19_ready_0 | requestReadLane_6[20] & output_20_ready_0
    | requestReadLane_6[21] & output_21_ready_0 | requestReadLane_6[22] & output_22_ready_0 | requestReadLane_6[23] & output_23_ready_0 | requestReadLane_6[24] & output_24_ready_0 | requestReadLane_6[25] & output_25_ready_0
    | requestReadLane_6[26] & output_26_ready_0 | requestReadLane_6[27] & output_27_ready_0 | requestReadLane_6[28] & output_28_ready_0 | requestReadLane_6[29] & output_29_ready_0 | requestReadLane_6[30] & output_30_ready_0
    | requestReadLane_6[31] & output_31_ready_0;
  wire        input_6_ready_0 = free_6 & outReady_6;
  wire [31:0] inputSelect1H_6 = input_6_valid_0 & free_6 ? requestReadLane_6 : 32'h0;
  wire [31:0] _GEN_4 = _GEN_3 | inputSelect1H_6;
  wire [31:0] requestReadLane_7 = 32'h1 << input_7_bits_readLane_0;
  wire        free_7 = |(requestReadLane_7 & ~_GEN_4);
  wire        outReady_7 =
    requestReadLane_7[0] & output_0_ready_0 | requestReadLane_7[1] & output_1_ready_0 | requestReadLane_7[2] & output_2_ready_0 | requestReadLane_7[3] & output_3_ready_0 | requestReadLane_7[4] & output_4_ready_0 | requestReadLane_7[5]
    & output_5_ready_0 | requestReadLane_7[6] & output_6_ready_0 | requestReadLane_7[7] & output_7_ready_0 | requestReadLane_7[8] & output_8_ready_0 | requestReadLane_7[9] & output_9_ready_0 | requestReadLane_7[10] & output_10_ready_0
    | requestReadLane_7[11] & output_11_ready_0 | requestReadLane_7[12] & output_12_ready_0 | requestReadLane_7[13] & output_13_ready_0 | requestReadLane_7[14] & output_14_ready_0 | requestReadLane_7[15] & output_15_ready_0
    | requestReadLane_7[16] & output_16_ready_0 | requestReadLane_7[17] & output_17_ready_0 | requestReadLane_7[18] & output_18_ready_0 | requestReadLane_7[19] & output_19_ready_0 | requestReadLane_7[20] & output_20_ready_0
    | requestReadLane_7[21] & output_21_ready_0 | requestReadLane_7[22] & output_22_ready_0 | requestReadLane_7[23] & output_23_ready_0 | requestReadLane_7[24] & output_24_ready_0 | requestReadLane_7[25] & output_25_ready_0
    | requestReadLane_7[26] & output_26_ready_0 | requestReadLane_7[27] & output_27_ready_0 | requestReadLane_7[28] & output_28_ready_0 | requestReadLane_7[29] & output_29_ready_0 | requestReadLane_7[30] & output_30_ready_0
    | requestReadLane_7[31] & output_31_ready_0;
  wire        input_7_ready_0 = free_7 & outReady_7;
  wire [31:0] inputSelect1H_7 = input_7_valid_0 & free_7 ? requestReadLane_7 : 32'h0;
  wire [31:0] _GEN_5 = _GEN_4 | inputSelect1H_7;
  wire [31:0] requestReadLane_8 = 32'h1 << input_8_bits_readLane_0;
  wire        free_8 = |(requestReadLane_8 & ~_GEN_5);
  wire        outReady_8 =
    requestReadLane_8[0] & output_0_ready_0 | requestReadLane_8[1] & output_1_ready_0 | requestReadLane_8[2] & output_2_ready_0 | requestReadLane_8[3] & output_3_ready_0 | requestReadLane_8[4] & output_4_ready_0 | requestReadLane_8[5]
    & output_5_ready_0 | requestReadLane_8[6] & output_6_ready_0 | requestReadLane_8[7] & output_7_ready_0 | requestReadLane_8[8] & output_8_ready_0 | requestReadLane_8[9] & output_9_ready_0 | requestReadLane_8[10] & output_10_ready_0
    | requestReadLane_8[11] & output_11_ready_0 | requestReadLane_8[12] & output_12_ready_0 | requestReadLane_8[13] & output_13_ready_0 | requestReadLane_8[14] & output_14_ready_0 | requestReadLane_8[15] & output_15_ready_0
    | requestReadLane_8[16] & output_16_ready_0 | requestReadLane_8[17] & output_17_ready_0 | requestReadLane_8[18] & output_18_ready_0 | requestReadLane_8[19] & output_19_ready_0 | requestReadLane_8[20] & output_20_ready_0
    | requestReadLane_8[21] & output_21_ready_0 | requestReadLane_8[22] & output_22_ready_0 | requestReadLane_8[23] & output_23_ready_0 | requestReadLane_8[24] & output_24_ready_0 | requestReadLane_8[25] & output_25_ready_0
    | requestReadLane_8[26] & output_26_ready_0 | requestReadLane_8[27] & output_27_ready_0 | requestReadLane_8[28] & output_28_ready_0 | requestReadLane_8[29] & output_29_ready_0 | requestReadLane_8[30] & output_30_ready_0
    | requestReadLane_8[31] & output_31_ready_0;
  wire        input_8_ready_0 = free_8 & outReady_8;
  wire [31:0] inputSelect1H_8 = input_8_valid_0 & free_8 ? requestReadLane_8 : 32'h0;
  wire [31:0] _GEN_6 = _GEN_5 | inputSelect1H_8;
  wire [31:0] requestReadLane_9 = 32'h1 << input_9_bits_readLane_0;
  wire        free_9 = |(requestReadLane_9 & ~_GEN_6);
  wire        outReady_9 =
    requestReadLane_9[0] & output_0_ready_0 | requestReadLane_9[1] & output_1_ready_0 | requestReadLane_9[2] & output_2_ready_0 | requestReadLane_9[3] & output_3_ready_0 | requestReadLane_9[4] & output_4_ready_0 | requestReadLane_9[5]
    & output_5_ready_0 | requestReadLane_9[6] & output_6_ready_0 | requestReadLane_9[7] & output_7_ready_0 | requestReadLane_9[8] & output_8_ready_0 | requestReadLane_9[9] & output_9_ready_0 | requestReadLane_9[10] & output_10_ready_0
    | requestReadLane_9[11] & output_11_ready_0 | requestReadLane_9[12] & output_12_ready_0 | requestReadLane_9[13] & output_13_ready_0 | requestReadLane_9[14] & output_14_ready_0 | requestReadLane_9[15] & output_15_ready_0
    | requestReadLane_9[16] & output_16_ready_0 | requestReadLane_9[17] & output_17_ready_0 | requestReadLane_9[18] & output_18_ready_0 | requestReadLane_9[19] & output_19_ready_0 | requestReadLane_9[20] & output_20_ready_0
    | requestReadLane_9[21] & output_21_ready_0 | requestReadLane_9[22] & output_22_ready_0 | requestReadLane_9[23] & output_23_ready_0 | requestReadLane_9[24] & output_24_ready_0 | requestReadLane_9[25] & output_25_ready_0
    | requestReadLane_9[26] & output_26_ready_0 | requestReadLane_9[27] & output_27_ready_0 | requestReadLane_9[28] & output_28_ready_0 | requestReadLane_9[29] & output_29_ready_0 | requestReadLane_9[30] & output_30_ready_0
    | requestReadLane_9[31] & output_31_ready_0;
  wire        input_9_ready_0 = free_9 & outReady_9;
  wire [31:0] inputSelect1H_9 = input_9_valid_0 & free_9 ? requestReadLane_9 : 32'h0;
  wire [31:0] _GEN_7 = _GEN_6 | inputSelect1H_9;
  wire [31:0] requestReadLane_10 = 32'h1 << input_10_bits_readLane_0;
  wire        free_10 = |(requestReadLane_10 & ~_GEN_7);
  wire        outReady_10 =
    requestReadLane_10[0] & output_0_ready_0 | requestReadLane_10[1] & output_1_ready_0 | requestReadLane_10[2] & output_2_ready_0 | requestReadLane_10[3] & output_3_ready_0 | requestReadLane_10[4] & output_4_ready_0 | requestReadLane_10[5]
    & output_5_ready_0 | requestReadLane_10[6] & output_6_ready_0 | requestReadLane_10[7] & output_7_ready_0 | requestReadLane_10[8] & output_8_ready_0 | requestReadLane_10[9] & output_9_ready_0 | requestReadLane_10[10] & output_10_ready_0
    | requestReadLane_10[11] & output_11_ready_0 | requestReadLane_10[12] & output_12_ready_0 | requestReadLane_10[13] & output_13_ready_0 | requestReadLane_10[14] & output_14_ready_0 | requestReadLane_10[15] & output_15_ready_0
    | requestReadLane_10[16] & output_16_ready_0 | requestReadLane_10[17] & output_17_ready_0 | requestReadLane_10[18] & output_18_ready_0 | requestReadLane_10[19] & output_19_ready_0 | requestReadLane_10[20] & output_20_ready_0
    | requestReadLane_10[21] & output_21_ready_0 | requestReadLane_10[22] & output_22_ready_0 | requestReadLane_10[23] & output_23_ready_0 | requestReadLane_10[24] & output_24_ready_0 | requestReadLane_10[25] & output_25_ready_0
    | requestReadLane_10[26] & output_26_ready_0 | requestReadLane_10[27] & output_27_ready_0 | requestReadLane_10[28] & output_28_ready_0 | requestReadLane_10[29] & output_29_ready_0 | requestReadLane_10[30] & output_30_ready_0
    | requestReadLane_10[31] & output_31_ready_0;
  wire        input_10_ready_0 = free_10 & outReady_10;
  wire [31:0] inputSelect1H_10 = input_10_valid_0 & free_10 ? requestReadLane_10 : 32'h0;
  wire [31:0] _GEN_8 = _GEN_7 | inputSelect1H_10;
  wire [31:0] requestReadLane_11 = 32'h1 << input_11_bits_readLane_0;
  wire        free_11 = |(requestReadLane_11 & ~_GEN_8);
  wire        outReady_11 =
    requestReadLane_11[0] & output_0_ready_0 | requestReadLane_11[1] & output_1_ready_0 | requestReadLane_11[2] & output_2_ready_0 | requestReadLane_11[3] & output_3_ready_0 | requestReadLane_11[4] & output_4_ready_0 | requestReadLane_11[5]
    & output_5_ready_0 | requestReadLane_11[6] & output_6_ready_0 | requestReadLane_11[7] & output_7_ready_0 | requestReadLane_11[8] & output_8_ready_0 | requestReadLane_11[9] & output_9_ready_0 | requestReadLane_11[10] & output_10_ready_0
    | requestReadLane_11[11] & output_11_ready_0 | requestReadLane_11[12] & output_12_ready_0 | requestReadLane_11[13] & output_13_ready_0 | requestReadLane_11[14] & output_14_ready_0 | requestReadLane_11[15] & output_15_ready_0
    | requestReadLane_11[16] & output_16_ready_0 | requestReadLane_11[17] & output_17_ready_0 | requestReadLane_11[18] & output_18_ready_0 | requestReadLane_11[19] & output_19_ready_0 | requestReadLane_11[20] & output_20_ready_0
    | requestReadLane_11[21] & output_21_ready_0 | requestReadLane_11[22] & output_22_ready_0 | requestReadLane_11[23] & output_23_ready_0 | requestReadLane_11[24] & output_24_ready_0 | requestReadLane_11[25] & output_25_ready_0
    | requestReadLane_11[26] & output_26_ready_0 | requestReadLane_11[27] & output_27_ready_0 | requestReadLane_11[28] & output_28_ready_0 | requestReadLane_11[29] & output_29_ready_0 | requestReadLane_11[30] & output_30_ready_0
    | requestReadLane_11[31] & output_31_ready_0;
  wire        input_11_ready_0 = free_11 & outReady_11;
  wire [31:0] inputSelect1H_11 = input_11_valid_0 & free_11 ? requestReadLane_11 : 32'h0;
  wire [31:0] _GEN_9 = _GEN_8 | inputSelect1H_11;
  wire [31:0] requestReadLane_12 = 32'h1 << input_12_bits_readLane_0;
  wire        free_12 = |(requestReadLane_12 & ~_GEN_9);
  wire        outReady_12 =
    requestReadLane_12[0] & output_0_ready_0 | requestReadLane_12[1] & output_1_ready_0 | requestReadLane_12[2] & output_2_ready_0 | requestReadLane_12[3] & output_3_ready_0 | requestReadLane_12[4] & output_4_ready_0 | requestReadLane_12[5]
    & output_5_ready_0 | requestReadLane_12[6] & output_6_ready_0 | requestReadLane_12[7] & output_7_ready_0 | requestReadLane_12[8] & output_8_ready_0 | requestReadLane_12[9] & output_9_ready_0 | requestReadLane_12[10] & output_10_ready_0
    | requestReadLane_12[11] & output_11_ready_0 | requestReadLane_12[12] & output_12_ready_0 | requestReadLane_12[13] & output_13_ready_0 | requestReadLane_12[14] & output_14_ready_0 | requestReadLane_12[15] & output_15_ready_0
    | requestReadLane_12[16] & output_16_ready_0 | requestReadLane_12[17] & output_17_ready_0 | requestReadLane_12[18] & output_18_ready_0 | requestReadLane_12[19] & output_19_ready_0 | requestReadLane_12[20] & output_20_ready_0
    | requestReadLane_12[21] & output_21_ready_0 | requestReadLane_12[22] & output_22_ready_0 | requestReadLane_12[23] & output_23_ready_0 | requestReadLane_12[24] & output_24_ready_0 | requestReadLane_12[25] & output_25_ready_0
    | requestReadLane_12[26] & output_26_ready_0 | requestReadLane_12[27] & output_27_ready_0 | requestReadLane_12[28] & output_28_ready_0 | requestReadLane_12[29] & output_29_ready_0 | requestReadLane_12[30] & output_30_ready_0
    | requestReadLane_12[31] & output_31_ready_0;
  wire        input_12_ready_0 = free_12 & outReady_12;
  wire [31:0] inputSelect1H_12 = input_12_valid_0 & free_12 ? requestReadLane_12 : 32'h0;
  wire [31:0] _GEN_10 = _GEN_9 | inputSelect1H_12;
  wire [31:0] requestReadLane_13 = 32'h1 << input_13_bits_readLane_0;
  wire        free_13 = |(requestReadLane_13 & ~_GEN_10);
  wire        outReady_13 =
    requestReadLane_13[0] & output_0_ready_0 | requestReadLane_13[1] & output_1_ready_0 | requestReadLane_13[2] & output_2_ready_0 | requestReadLane_13[3] & output_3_ready_0 | requestReadLane_13[4] & output_4_ready_0 | requestReadLane_13[5]
    & output_5_ready_0 | requestReadLane_13[6] & output_6_ready_0 | requestReadLane_13[7] & output_7_ready_0 | requestReadLane_13[8] & output_8_ready_0 | requestReadLane_13[9] & output_9_ready_0 | requestReadLane_13[10] & output_10_ready_0
    | requestReadLane_13[11] & output_11_ready_0 | requestReadLane_13[12] & output_12_ready_0 | requestReadLane_13[13] & output_13_ready_0 | requestReadLane_13[14] & output_14_ready_0 | requestReadLane_13[15] & output_15_ready_0
    | requestReadLane_13[16] & output_16_ready_0 | requestReadLane_13[17] & output_17_ready_0 | requestReadLane_13[18] & output_18_ready_0 | requestReadLane_13[19] & output_19_ready_0 | requestReadLane_13[20] & output_20_ready_0
    | requestReadLane_13[21] & output_21_ready_0 | requestReadLane_13[22] & output_22_ready_0 | requestReadLane_13[23] & output_23_ready_0 | requestReadLane_13[24] & output_24_ready_0 | requestReadLane_13[25] & output_25_ready_0
    | requestReadLane_13[26] & output_26_ready_0 | requestReadLane_13[27] & output_27_ready_0 | requestReadLane_13[28] & output_28_ready_0 | requestReadLane_13[29] & output_29_ready_0 | requestReadLane_13[30] & output_30_ready_0
    | requestReadLane_13[31] & output_31_ready_0;
  wire        input_13_ready_0 = free_13 & outReady_13;
  wire [31:0] inputSelect1H_13 = input_13_valid_0 & free_13 ? requestReadLane_13 : 32'h0;
  wire [31:0] _GEN_11 = _GEN_10 | inputSelect1H_13;
  wire [31:0] requestReadLane_14 = 32'h1 << input_14_bits_readLane_0;
  wire        free_14 = |(requestReadLane_14 & ~_GEN_11);
  wire        outReady_14 =
    requestReadLane_14[0] & output_0_ready_0 | requestReadLane_14[1] & output_1_ready_0 | requestReadLane_14[2] & output_2_ready_0 | requestReadLane_14[3] & output_3_ready_0 | requestReadLane_14[4] & output_4_ready_0 | requestReadLane_14[5]
    & output_5_ready_0 | requestReadLane_14[6] & output_6_ready_0 | requestReadLane_14[7] & output_7_ready_0 | requestReadLane_14[8] & output_8_ready_0 | requestReadLane_14[9] & output_9_ready_0 | requestReadLane_14[10] & output_10_ready_0
    | requestReadLane_14[11] & output_11_ready_0 | requestReadLane_14[12] & output_12_ready_0 | requestReadLane_14[13] & output_13_ready_0 | requestReadLane_14[14] & output_14_ready_0 | requestReadLane_14[15] & output_15_ready_0
    | requestReadLane_14[16] & output_16_ready_0 | requestReadLane_14[17] & output_17_ready_0 | requestReadLane_14[18] & output_18_ready_0 | requestReadLane_14[19] & output_19_ready_0 | requestReadLane_14[20] & output_20_ready_0
    | requestReadLane_14[21] & output_21_ready_0 | requestReadLane_14[22] & output_22_ready_0 | requestReadLane_14[23] & output_23_ready_0 | requestReadLane_14[24] & output_24_ready_0 | requestReadLane_14[25] & output_25_ready_0
    | requestReadLane_14[26] & output_26_ready_0 | requestReadLane_14[27] & output_27_ready_0 | requestReadLane_14[28] & output_28_ready_0 | requestReadLane_14[29] & output_29_ready_0 | requestReadLane_14[30] & output_30_ready_0
    | requestReadLane_14[31] & output_31_ready_0;
  wire        input_14_ready_0 = free_14 & outReady_14;
  wire [31:0] inputSelect1H_14 = input_14_valid_0 & free_14 ? requestReadLane_14 : 32'h0;
  wire [31:0] _GEN_12 = _GEN_11 | inputSelect1H_14;
  wire [31:0] requestReadLane_15 = 32'h1 << input_15_bits_readLane_0;
  wire        free_15 = |(requestReadLane_15 & ~_GEN_12);
  wire        outReady_15 =
    requestReadLane_15[0] & output_0_ready_0 | requestReadLane_15[1] & output_1_ready_0 | requestReadLane_15[2] & output_2_ready_0 | requestReadLane_15[3] & output_3_ready_0 | requestReadLane_15[4] & output_4_ready_0 | requestReadLane_15[5]
    & output_5_ready_0 | requestReadLane_15[6] & output_6_ready_0 | requestReadLane_15[7] & output_7_ready_0 | requestReadLane_15[8] & output_8_ready_0 | requestReadLane_15[9] & output_9_ready_0 | requestReadLane_15[10] & output_10_ready_0
    | requestReadLane_15[11] & output_11_ready_0 | requestReadLane_15[12] & output_12_ready_0 | requestReadLane_15[13] & output_13_ready_0 | requestReadLane_15[14] & output_14_ready_0 | requestReadLane_15[15] & output_15_ready_0
    | requestReadLane_15[16] & output_16_ready_0 | requestReadLane_15[17] & output_17_ready_0 | requestReadLane_15[18] & output_18_ready_0 | requestReadLane_15[19] & output_19_ready_0 | requestReadLane_15[20] & output_20_ready_0
    | requestReadLane_15[21] & output_21_ready_0 | requestReadLane_15[22] & output_22_ready_0 | requestReadLane_15[23] & output_23_ready_0 | requestReadLane_15[24] & output_24_ready_0 | requestReadLane_15[25] & output_25_ready_0
    | requestReadLane_15[26] & output_26_ready_0 | requestReadLane_15[27] & output_27_ready_0 | requestReadLane_15[28] & output_28_ready_0 | requestReadLane_15[29] & output_29_ready_0 | requestReadLane_15[30] & output_30_ready_0
    | requestReadLane_15[31] & output_31_ready_0;
  wire        input_15_ready_0 = free_15 & outReady_15;
  wire [31:0] inputSelect1H_15 = input_15_valid_0 & free_15 ? requestReadLane_15 : 32'h0;
  wire [31:0] _GEN_13 = _GEN_12 | inputSelect1H_15;
  wire [31:0] requestReadLane_16 = 32'h1 << input_16_bits_readLane_0;
  wire        free_16 = |(requestReadLane_16 & ~_GEN_13);
  wire        outReady_16 =
    requestReadLane_16[0] & output_0_ready_0 | requestReadLane_16[1] & output_1_ready_0 | requestReadLane_16[2] & output_2_ready_0 | requestReadLane_16[3] & output_3_ready_0 | requestReadLane_16[4] & output_4_ready_0 | requestReadLane_16[5]
    & output_5_ready_0 | requestReadLane_16[6] & output_6_ready_0 | requestReadLane_16[7] & output_7_ready_0 | requestReadLane_16[8] & output_8_ready_0 | requestReadLane_16[9] & output_9_ready_0 | requestReadLane_16[10] & output_10_ready_0
    | requestReadLane_16[11] & output_11_ready_0 | requestReadLane_16[12] & output_12_ready_0 | requestReadLane_16[13] & output_13_ready_0 | requestReadLane_16[14] & output_14_ready_0 | requestReadLane_16[15] & output_15_ready_0
    | requestReadLane_16[16] & output_16_ready_0 | requestReadLane_16[17] & output_17_ready_0 | requestReadLane_16[18] & output_18_ready_0 | requestReadLane_16[19] & output_19_ready_0 | requestReadLane_16[20] & output_20_ready_0
    | requestReadLane_16[21] & output_21_ready_0 | requestReadLane_16[22] & output_22_ready_0 | requestReadLane_16[23] & output_23_ready_0 | requestReadLane_16[24] & output_24_ready_0 | requestReadLane_16[25] & output_25_ready_0
    | requestReadLane_16[26] & output_26_ready_0 | requestReadLane_16[27] & output_27_ready_0 | requestReadLane_16[28] & output_28_ready_0 | requestReadLane_16[29] & output_29_ready_0 | requestReadLane_16[30] & output_30_ready_0
    | requestReadLane_16[31] & output_31_ready_0;
  wire        input_16_ready_0 = free_16 & outReady_16;
  wire [31:0] inputSelect1H_16 = input_16_valid_0 & free_16 ? requestReadLane_16 : 32'h0;
  wire [31:0] _GEN_14 = _GEN_13 | inputSelect1H_16;
  wire [31:0] requestReadLane_17 = 32'h1 << input_17_bits_readLane_0;
  wire        free_17 = |(requestReadLane_17 & ~_GEN_14);
  wire        outReady_17 =
    requestReadLane_17[0] & output_0_ready_0 | requestReadLane_17[1] & output_1_ready_0 | requestReadLane_17[2] & output_2_ready_0 | requestReadLane_17[3] & output_3_ready_0 | requestReadLane_17[4] & output_4_ready_0 | requestReadLane_17[5]
    & output_5_ready_0 | requestReadLane_17[6] & output_6_ready_0 | requestReadLane_17[7] & output_7_ready_0 | requestReadLane_17[8] & output_8_ready_0 | requestReadLane_17[9] & output_9_ready_0 | requestReadLane_17[10] & output_10_ready_0
    | requestReadLane_17[11] & output_11_ready_0 | requestReadLane_17[12] & output_12_ready_0 | requestReadLane_17[13] & output_13_ready_0 | requestReadLane_17[14] & output_14_ready_0 | requestReadLane_17[15] & output_15_ready_0
    | requestReadLane_17[16] & output_16_ready_0 | requestReadLane_17[17] & output_17_ready_0 | requestReadLane_17[18] & output_18_ready_0 | requestReadLane_17[19] & output_19_ready_0 | requestReadLane_17[20] & output_20_ready_0
    | requestReadLane_17[21] & output_21_ready_0 | requestReadLane_17[22] & output_22_ready_0 | requestReadLane_17[23] & output_23_ready_0 | requestReadLane_17[24] & output_24_ready_0 | requestReadLane_17[25] & output_25_ready_0
    | requestReadLane_17[26] & output_26_ready_0 | requestReadLane_17[27] & output_27_ready_0 | requestReadLane_17[28] & output_28_ready_0 | requestReadLane_17[29] & output_29_ready_0 | requestReadLane_17[30] & output_30_ready_0
    | requestReadLane_17[31] & output_31_ready_0;
  wire        input_17_ready_0 = free_17 & outReady_17;
  wire [31:0] inputSelect1H_17 = input_17_valid_0 & free_17 ? requestReadLane_17 : 32'h0;
  wire [31:0] _GEN_15 = _GEN_14 | inputSelect1H_17;
  wire [31:0] requestReadLane_18 = 32'h1 << input_18_bits_readLane_0;
  wire        free_18 = |(requestReadLane_18 & ~_GEN_15);
  wire        outReady_18 =
    requestReadLane_18[0] & output_0_ready_0 | requestReadLane_18[1] & output_1_ready_0 | requestReadLane_18[2] & output_2_ready_0 | requestReadLane_18[3] & output_3_ready_0 | requestReadLane_18[4] & output_4_ready_0 | requestReadLane_18[5]
    & output_5_ready_0 | requestReadLane_18[6] & output_6_ready_0 | requestReadLane_18[7] & output_7_ready_0 | requestReadLane_18[8] & output_8_ready_0 | requestReadLane_18[9] & output_9_ready_0 | requestReadLane_18[10] & output_10_ready_0
    | requestReadLane_18[11] & output_11_ready_0 | requestReadLane_18[12] & output_12_ready_0 | requestReadLane_18[13] & output_13_ready_0 | requestReadLane_18[14] & output_14_ready_0 | requestReadLane_18[15] & output_15_ready_0
    | requestReadLane_18[16] & output_16_ready_0 | requestReadLane_18[17] & output_17_ready_0 | requestReadLane_18[18] & output_18_ready_0 | requestReadLane_18[19] & output_19_ready_0 | requestReadLane_18[20] & output_20_ready_0
    | requestReadLane_18[21] & output_21_ready_0 | requestReadLane_18[22] & output_22_ready_0 | requestReadLane_18[23] & output_23_ready_0 | requestReadLane_18[24] & output_24_ready_0 | requestReadLane_18[25] & output_25_ready_0
    | requestReadLane_18[26] & output_26_ready_0 | requestReadLane_18[27] & output_27_ready_0 | requestReadLane_18[28] & output_28_ready_0 | requestReadLane_18[29] & output_29_ready_0 | requestReadLane_18[30] & output_30_ready_0
    | requestReadLane_18[31] & output_31_ready_0;
  wire        input_18_ready_0 = free_18 & outReady_18;
  wire [31:0] inputSelect1H_18 = input_18_valid_0 & free_18 ? requestReadLane_18 : 32'h0;
  wire [31:0] _GEN_16 = _GEN_15 | inputSelect1H_18;
  wire [31:0] requestReadLane_19 = 32'h1 << input_19_bits_readLane_0;
  wire        free_19 = |(requestReadLane_19 & ~_GEN_16);
  wire        outReady_19 =
    requestReadLane_19[0] & output_0_ready_0 | requestReadLane_19[1] & output_1_ready_0 | requestReadLane_19[2] & output_2_ready_0 | requestReadLane_19[3] & output_3_ready_0 | requestReadLane_19[4] & output_4_ready_0 | requestReadLane_19[5]
    & output_5_ready_0 | requestReadLane_19[6] & output_6_ready_0 | requestReadLane_19[7] & output_7_ready_0 | requestReadLane_19[8] & output_8_ready_0 | requestReadLane_19[9] & output_9_ready_0 | requestReadLane_19[10] & output_10_ready_0
    | requestReadLane_19[11] & output_11_ready_0 | requestReadLane_19[12] & output_12_ready_0 | requestReadLane_19[13] & output_13_ready_0 | requestReadLane_19[14] & output_14_ready_0 | requestReadLane_19[15] & output_15_ready_0
    | requestReadLane_19[16] & output_16_ready_0 | requestReadLane_19[17] & output_17_ready_0 | requestReadLane_19[18] & output_18_ready_0 | requestReadLane_19[19] & output_19_ready_0 | requestReadLane_19[20] & output_20_ready_0
    | requestReadLane_19[21] & output_21_ready_0 | requestReadLane_19[22] & output_22_ready_0 | requestReadLane_19[23] & output_23_ready_0 | requestReadLane_19[24] & output_24_ready_0 | requestReadLane_19[25] & output_25_ready_0
    | requestReadLane_19[26] & output_26_ready_0 | requestReadLane_19[27] & output_27_ready_0 | requestReadLane_19[28] & output_28_ready_0 | requestReadLane_19[29] & output_29_ready_0 | requestReadLane_19[30] & output_30_ready_0
    | requestReadLane_19[31] & output_31_ready_0;
  wire        input_19_ready_0 = free_19 & outReady_19;
  wire [31:0] inputSelect1H_19 = input_19_valid_0 & free_19 ? requestReadLane_19 : 32'h0;
  wire [31:0] _GEN_17 = _GEN_16 | inputSelect1H_19;
  wire [31:0] requestReadLane_20 = 32'h1 << input_20_bits_readLane_0;
  wire        free_20 = |(requestReadLane_20 & ~_GEN_17);
  wire        outReady_20 =
    requestReadLane_20[0] & output_0_ready_0 | requestReadLane_20[1] & output_1_ready_0 | requestReadLane_20[2] & output_2_ready_0 | requestReadLane_20[3] & output_3_ready_0 | requestReadLane_20[4] & output_4_ready_0 | requestReadLane_20[5]
    & output_5_ready_0 | requestReadLane_20[6] & output_6_ready_0 | requestReadLane_20[7] & output_7_ready_0 | requestReadLane_20[8] & output_8_ready_0 | requestReadLane_20[9] & output_9_ready_0 | requestReadLane_20[10] & output_10_ready_0
    | requestReadLane_20[11] & output_11_ready_0 | requestReadLane_20[12] & output_12_ready_0 | requestReadLane_20[13] & output_13_ready_0 | requestReadLane_20[14] & output_14_ready_0 | requestReadLane_20[15] & output_15_ready_0
    | requestReadLane_20[16] & output_16_ready_0 | requestReadLane_20[17] & output_17_ready_0 | requestReadLane_20[18] & output_18_ready_0 | requestReadLane_20[19] & output_19_ready_0 | requestReadLane_20[20] & output_20_ready_0
    | requestReadLane_20[21] & output_21_ready_0 | requestReadLane_20[22] & output_22_ready_0 | requestReadLane_20[23] & output_23_ready_0 | requestReadLane_20[24] & output_24_ready_0 | requestReadLane_20[25] & output_25_ready_0
    | requestReadLane_20[26] & output_26_ready_0 | requestReadLane_20[27] & output_27_ready_0 | requestReadLane_20[28] & output_28_ready_0 | requestReadLane_20[29] & output_29_ready_0 | requestReadLane_20[30] & output_30_ready_0
    | requestReadLane_20[31] & output_31_ready_0;
  wire        input_20_ready_0 = free_20 & outReady_20;
  wire [31:0] inputSelect1H_20 = input_20_valid_0 & free_20 ? requestReadLane_20 : 32'h0;
  wire [31:0] _GEN_18 = _GEN_17 | inputSelect1H_20;
  wire [31:0] requestReadLane_21 = 32'h1 << input_21_bits_readLane_0;
  wire        free_21 = |(requestReadLane_21 & ~_GEN_18);
  wire        outReady_21 =
    requestReadLane_21[0] & output_0_ready_0 | requestReadLane_21[1] & output_1_ready_0 | requestReadLane_21[2] & output_2_ready_0 | requestReadLane_21[3] & output_3_ready_0 | requestReadLane_21[4] & output_4_ready_0 | requestReadLane_21[5]
    & output_5_ready_0 | requestReadLane_21[6] & output_6_ready_0 | requestReadLane_21[7] & output_7_ready_0 | requestReadLane_21[8] & output_8_ready_0 | requestReadLane_21[9] & output_9_ready_0 | requestReadLane_21[10] & output_10_ready_0
    | requestReadLane_21[11] & output_11_ready_0 | requestReadLane_21[12] & output_12_ready_0 | requestReadLane_21[13] & output_13_ready_0 | requestReadLane_21[14] & output_14_ready_0 | requestReadLane_21[15] & output_15_ready_0
    | requestReadLane_21[16] & output_16_ready_0 | requestReadLane_21[17] & output_17_ready_0 | requestReadLane_21[18] & output_18_ready_0 | requestReadLane_21[19] & output_19_ready_0 | requestReadLane_21[20] & output_20_ready_0
    | requestReadLane_21[21] & output_21_ready_0 | requestReadLane_21[22] & output_22_ready_0 | requestReadLane_21[23] & output_23_ready_0 | requestReadLane_21[24] & output_24_ready_0 | requestReadLane_21[25] & output_25_ready_0
    | requestReadLane_21[26] & output_26_ready_0 | requestReadLane_21[27] & output_27_ready_0 | requestReadLane_21[28] & output_28_ready_0 | requestReadLane_21[29] & output_29_ready_0 | requestReadLane_21[30] & output_30_ready_0
    | requestReadLane_21[31] & output_31_ready_0;
  wire        input_21_ready_0 = free_21 & outReady_21;
  wire [31:0] inputSelect1H_21 = input_21_valid_0 & free_21 ? requestReadLane_21 : 32'h0;
  wire [31:0] _GEN_19 = _GEN_18 | inputSelect1H_21;
  wire [31:0] requestReadLane_22 = 32'h1 << input_22_bits_readLane_0;
  wire        free_22 = |(requestReadLane_22 & ~_GEN_19);
  wire        outReady_22 =
    requestReadLane_22[0] & output_0_ready_0 | requestReadLane_22[1] & output_1_ready_0 | requestReadLane_22[2] & output_2_ready_0 | requestReadLane_22[3] & output_3_ready_0 | requestReadLane_22[4] & output_4_ready_0 | requestReadLane_22[5]
    & output_5_ready_0 | requestReadLane_22[6] & output_6_ready_0 | requestReadLane_22[7] & output_7_ready_0 | requestReadLane_22[8] & output_8_ready_0 | requestReadLane_22[9] & output_9_ready_0 | requestReadLane_22[10] & output_10_ready_0
    | requestReadLane_22[11] & output_11_ready_0 | requestReadLane_22[12] & output_12_ready_0 | requestReadLane_22[13] & output_13_ready_0 | requestReadLane_22[14] & output_14_ready_0 | requestReadLane_22[15] & output_15_ready_0
    | requestReadLane_22[16] & output_16_ready_0 | requestReadLane_22[17] & output_17_ready_0 | requestReadLane_22[18] & output_18_ready_0 | requestReadLane_22[19] & output_19_ready_0 | requestReadLane_22[20] & output_20_ready_0
    | requestReadLane_22[21] & output_21_ready_0 | requestReadLane_22[22] & output_22_ready_0 | requestReadLane_22[23] & output_23_ready_0 | requestReadLane_22[24] & output_24_ready_0 | requestReadLane_22[25] & output_25_ready_0
    | requestReadLane_22[26] & output_26_ready_0 | requestReadLane_22[27] & output_27_ready_0 | requestReadLane_22[28] & output_28_ready_0 | requestReadLane_22[29] & output_29_ready_0 | requestReadLane_22[30] & output_30_ready_0
    | requestReadLane_22[31] & output_31_ready_0;
  wire        input_22_ready_0 = free_22 & outReady_22;
  wire [31:0] inputSelect1H_22 = input_22_valid_0 & free_22 ? requestReadLane_22 : 32'h0;
  wire [31:0] _GEN_20 = _GEN_19 | inputSelect1H_22;
  wire [31:0] requestReadLane_23 = 32'h1 << input_23_bits_readLane_0;
  wire        free_23 = |(requestReadLane_23 & ~_GEN_20);
  wire        outReady_23 =
    requestReadLane_23[0] & output_0_ready_0 | requestReadLane_23[1] & output_1_ready_0 | requestReadLane_23[2] & output_2_ready_0 | requestReadLane_23[3] & output_3_ready_0 | requestReadLane_23[4] & output_4_ready_0 | requestReadLane_23[5]
    & output_5_ready_0 | requestReadLane_23[6] & output_6_ready_0 | requestReadLane_23[7] & output_7_ready_0 | requestReadLane_23[8] & output_8_ready_0 | requestReadLane_23[9] & output_9_ready_0 | requestReadLane_23[10] & output_10_ready_0
    | requestReadLane_23[11] & output_11_ready_0 | requestReadLane_23[12] & output_12_ready_0 | requestReadLane_23[13] & output_13_ready_0 | requestReadLane_23[14] & output_14_ready_0 | requestReadLane_23[15] & output_15_ready_0
    | requestReadLane_23[16] & output_16_ready_0 | requestReadLane_23[17] & output_17_ready_0 | requestReadLane_23[18] & output_18_ready_0 | requestReadLane_23[19] & output_19_ready_0 | requestReadLane_23[20] & output_20_ready_0
    | requestReadLane_23[21] & output_21_ready_0 | requestReadLane_23[22] & output_22_ready_0 | requestReadLane_23[23] & output_23_ready_0 | requestReadLane_23[24] & output_24_ready_0 | requestReadLane_23[25] & output_25_ready_0
    | requestReadLane_23[26] & output_26_ready_0 | requestReadLane_23[27] & output_27_ready_0 | requestReadLane_23[28] & output_28_ready_0 | requestReadLane_23[29] & output_29_ready_0 | requestReadLane_23[30] & output_30_ready_0
    | requestReadLane_23[31] & output_31_ready_0;
  wire        input_23_ready_0 = free_23 & outReady_23;
  wire [31:0] inputSelect1H_23 = input_23_valid_0 & free_23 ? requestReadLane_23 : 32'h0;
  wire [31:0] _GEN_21 = _GEN_20 | inputSelect1H_23;
  wire [31:0] requestReadLane_24 = 32'h1 << input_24_bits_readLane_0;
  wire        free_24 = |(requestReadLane_24 & ~_GEN_21);
  wire        outReady_24 =
    requestReadLane_24[0] & output_0_ready_0 | requestReadLane_24[1] & output_1_ready_0 | requestReadLane_24[2] & output_2_ready_0 | requestReadLane_24[3] & output_3_ready_0 | requestReadLane_24[4] & output_4_ready_0 | requestReadLane_24[5]
    & output_5_ready_0 | requestReadLane_24[6] & output_6_ready_0 | requestReadLane_24[7] & output_7_ready_0 | requestReadLane_24[8] & output_8_ready_0 | requestReadLane_24[9] & output_9_ready_0 | requestReadLane_24[10] & output_10_ready_0
    | requestReadLane_24[11] & output_11_ready_0 | requestReadLane_24[12] & output_12_ready_0 | requestReadLane_24[13] & output_13_ready_0 | requestReadLane_24[14] & output_14_ready_0 | requestReadLane_24[15] & output_15_ready_0
    | requestReadLane_24[16] & output_16_ready_0 | requestReadLane_24[17] & output_17_ready_0 | requestReadLane_24[18] & output_18_ready_0 | requestReadLane_24[19] & output_19_ready_0 | requestReadLane_24[20] & output_20_ready_0
    | requestReadLane_24[21] & output_21_ready_0 | requestReadLane_24[22] & output_22_ready_0 | requestReadLane_24[23] & output_23_ready_0 | requestReadLane_24[24] & output_24_ready_0 | requestReadLane_24[25] & output_25_ready_0
    | requestReadLane_24[26] & output_26_ready_0 | requestReadLane_24[27] & output_27_ready_0 | requestReadLane_24[28] & output_28_ready_0 | requestReadLane_24[29] & output_29_ready_0 | requestReadLane_24[30] & output_30_ready_0
    | requestReadLane_24[31] & output_31_ready_0;
  wire        input_24_ready_0 = free_24 & outReady_24;
  wire [31:0] inputSelect1H_24 = input_24_valid_0 & free_24 ? requestReadLane_24 : 32'h0;
  wire [31:0] _GEN_22 = _GEN_21 | inputSelect1H_24;
  wire [31:0] requestReadLane_25 = 32'h1 << input_25_bits_readLane_0;
  wire        free_25 = |(requestReadLane_25 & ~_GEN_22);
  wire        outReady_25 =
    requestReadLane_25[0] & output_0_ready_0 | requestReadLane_25[1] & output_1_ready_0 | requestReadLane_25[2] & output_2_ready_0 | requestReadLane_25[3] & output_3_ready_0 | requestReadLane_25[4] & output_4_ready_0 | requestReadLane_25[5]
    & output_5_ready_0 | requestReadLane_25[6] & output_6_ready_0 | requestReadLane_25[7] & output_7_ready_0 | requestReadLane_25[8] & output_8_ready_0 | requestReadLane_25[9] & output_9_ready_0 | requestReadLane_25[10] & output_10_ready_0
    | requestReadLane_25[11] & output_11_ready_0 | requestReadLane_25[12] & output_12_ready_0 | requestReadLane_25[13] & output_13_ready_0 | requestReadLane_25[14] & output_14_ready_0 | requestReadLane_25[15] & output_15_ready_0
    | requestReadLane_25[16] & output_16_ready_0 | requestReadLane_25[17] & output_17_ready_0 | requestReadLane_25[18] & output_18_ready_0 | requestReadLane_25[19] & output_19_ready_0 | requestReadLane_25[20] & output_20_ready_0
    | requestReadLane_25[21] & output_21_ready_0 | requestReadLane_25[22] & output_22_ready_0 | requestReadLane_25[23] & output_23_ready_0 | requestReadLane_25[24] & output_24_ready_0 | requestReadLane_25[25] & output_25_ready_0
    | requestReadLane_25[26] & output_26_ready_0 | requestReadLane_25[27] & output_27_ready_0 | requestReadLane_25[28] & output_28_ready_0 | requestReadLane_25[29] & output_29_ready_0 | requestReadLane_25[30] & output_30_ready_0
    | requestReadLane_25[31] & output_31_ready_0;
  wire        input_25_ready_0 = free_25 & outReady_25;
  wire [31:0] inputSelect1H_25 = input_25_valid_0 & free_25 ? requestReadLane_25 : 32'h0;
  wire [31:0] _GEN_23 = _GEN_22 | inputSelect1H_25;
  wire [31:0] requestReadLane_26 = 32'h1 << input_26_bits_readLane_0;
  wire        free_26 = |(requestReadLane_26 & ~_GEN_23);
  wire        outReady_26 =
    requestReadLane_26[0] & output_0_ready_0 | requestReadLane_26[1] & output_1_ready_0 | requestReadLane_26[2] & output_2_ready_0 | requestReadLane_26[3] & output_3_ready_0 | requestReadLane_26[4] & output_4_ready_0 | requestReadLane_26[5]
    & output_5_ready_0 | requestReadLane_26[6] & output_6_ready_0 | requestReadLane_26[7] & output_7_ready_0 | requestReadLane_26[8] & output_8_ready_0 | requestReadLane_26[9] & output_9_ready_0 | requestReadLane_26[10] & output_10_ready_0
    | requestReadLane_26[11] & output_11_ready_0 | requestReadLane_26[12] & output_12_ready_0 | requestReadLane_26[13] & output_13_ready_0 | requestReadLane_26[14] & output_14_ready_0 | requestReadLane_26[15] & output_15_ready_0
    | requestReadLane_26[16] & output_16_ready_0 | requestReadLane_26[17] & output_17_ready_0 | requestReadLane_26[18] & output_18_ready_0 | requestReadLane_26[19] & output_19_ready_0 | requestReadLane_26[20] & output_20_ready_0
    | requestReadLane_26[21] & output_21_ready_0 | requestReadLane_26[22] & output_22_ready_0 | requestReadLane_26[23] & output_23_ready_0 | requestReadLane_26[24] & output_24_ready_0 | requestReadLane_26[25] & output_25_ready_0
    | requestReadLane_26[26] & output_26_ready_0 | requestReadLane_26[27] & output_27_ready_0 | requestReadLane_26[28] & output_28_ready_0 | requestReadLane_26[29] & output_29_ready_0 | requestReadLane_26[30] & output_30_ready_0
    | requestReadLane_26[31] & output_31_ready_0;
  wire        input_26_ready_0 = free_26 & outReady_26;
  wire [31:0] inputSelect1H_26 = input_26_valid_0 & free_26 ? requestReadLane_26 : 32'h0;
  wire [31:0] _GEN_24 = _GEN_23 | inputSelect1H_26;
  wire [31:0] requestReadLane_27 = 32'h1 << input_27_bits_readLane_0;
  wire        free_27 = |(requestReadLane_27 & ~_GEN_24);
  wire        outReady_27 =
    requestReadLane_27[0] & output_0_ready_0 | requestReadLane_27[1] & output_1_ready_0 | requestReadLane_27[2] & output_2_ready_0 | requestReadLane_27[3] & output_3_ready_0 | requestReadLane_27[4] & output_4_ready_0 | requestReadLane_27[5]
    & output_5_ready_0 | requestReadLane_27[6] & output_6_ready_0 | requestReadLane_27[7] & output_7_ready_0 | requestReadLane_27[8] & output_8_ready_0 | requestReadLane_27[9] & output_9_ready_0 | requestReadLane_27[10] & output_10_ready_0
    | requestReadLane_27[11] & output_11_ready_0 | requestReadLane_27[12] & output_12_ready_0 | requestReadLane_27[13] & output_13_ready_0 | requestReadLane_27[14] & output_14_ready_0 | requestReadLane_27[15] & output_15_ready_0
    | requestReadLane_27[16] & output_16_ready_0 | requestReadLane_27[17] & output_17_ready_0 | requestReadLane_27[18] & output_18_ready_0 | requestReadLane_27[19] & output_19_ready_0 | requestReadLane_27[20] & output_20_ready_0
    | requestReadLane_27[21] & output_21_ready_0 | requestReadLane_27[22] & output_22_ready_0 | requestReadLane_27[23] & output_23_ready_0 | requestReadLane_27[24] & output_24_ready_0 | requestReadLane_27[25] & output_25_ready_0
    | requestReadLane_27[26] & output_26_ready_0 | requestReadLane_27[27] & output_27_ready_0 | requestReadLane_27[28] & output_28_ready_0 | requestReadLane_27[29] & output_29_ready_0 | requestReadLane_27[30] & output_30_ready_0
    | requestReadLane_27[31] & output_31_ready_0;
  wire        input_27_ready_0 = free_27 & outReady_27;
  wire [31:0] inputSelect1H_27 = input_27_valid_0 & free_27 ? requestReadLane_27 : 32'h0;
  wire [31:0] _GEN_25 = _GEN_24 | inputSelect1H_27;
  wire [31:0] requestReadLane_28 = 32'h1 << input_28_bits_readLane_0;
  wire        free_28 = |(requestReadLane_28 & ~_GEN_25);
  wire        outReady_28 =
    requestReadLane_28[0] & output_0_ready_0 | requestReadLane_28[1] & output_1_ready_0 | requestReadLane_28[2] & output_2_ready_0 | requestReadLane_28[3] & output_3_ready_0 | requestReadLane_28[4] & output_4_ready_0 | requestReadLane_28[5]
    & output_5_ready_0 | requestReadLane_28[6] & output_6_ready_0 | requestReadLane_28[7] & output_7_ready_0 | requestReadLane_28[8] & output_8_ready_0 | requestReadLane_28[9] & output_9_ready_0 | requestReadLane_28[10] & output_10_ready_0
    | requestReadLane_28[11] & output_11_ready_0 | requestReadLane_28[12] & output_12_ready_0 | requestReadLane_28[13] & output_13_ready_0 | requestReadLane_28[14] & output_14_ready_0 | requestReadLane_28[15] & output_15_ready_0
    | requestReadLane_28[16] & output_16_ready_0 | requestReadLane_28[17] & output_17_ready_0 | requestReadLane_28[18] & output_18_ready_0 | requestReadLane_28[19] & output_19_ready_0 | requestReadLane_28[20] & output_20_ready_0
    | requestReadLane_28[21] & output_21_ready_0 | requestReadLane_28[22] & output_22_ready_0 | requestReadLane_28[23] & output_23_ready_0 | requestReadLane_28[24] & output_24_ready_0 | requestReadLane_28[25] & output_25_ready_0
    | requestReadLane_28[26] & output_26_ready_0 | requestReadLane_28[27] & output_27_ready_0 | requestReadLane_28[28] & output_28_ready_0 | requestReadLane_28[29] & output_29_ready_0 | requestReadLane_28[30] & output_30_ready_0
    | requestReadLane_28[31] & output_31_ready_0;
  wire        input_28_ready_0 = free_28 & outReady_28;
  wire [31:0] inputSelect1H_28 = input_28_valid_0 & free_28 ? requestReadLane_28 : 32'h0;
  wire [31:0] _GEN_26 = _GEN_25 | inputSelect1H_28;
  wire [31:0] requestReadLane_29 = 32'h1 << input_29_bits_readLane_0;
  wire        free_29 = |(requestReadLane_29 & ~_GEN_26);
  wire        outReady_29 =
    requestReadLane_29[0] & output_0_ready_0 | requestReadLane_29[1] & output_1_ready_0 | requestReadLane_29[2] & output_2_ready_0 | requestReadLane_29[3] & output_3_ready_0 | requestReadLane_29[4] & output_4_ready_0 | requestReadLane_29[5]
    & output_5_ready_0 | requestReadLane_29[6] & output_6_ready_0 | requestReadLane_29[7] & output_7_ready_0 | requestReadLane_29[8] & output_8_ready_0 | requestReadLane_29[9] & output_9_ready_0 | requestReadLane_29[10] & output_10_ready_0
    | requestReadLane_29[11] & output_11_ready_0 | requestReadLane_29[12] & output_12_ready_0 | requestReadLane_29[13] & output_13_ready_0 | requestReadLane_29[14] & output_14_ready_0 | requestReadLane_29[15] & output_15_ready_0
    | requestReadLane_29[16] & output_16_ready_0 | requestReadLane_29[17] & output_17_ready_0 | requestReadLane_29[18] & output_18_ready_0 | requestReadLane_29[19] & output_19_ready_0 | requestReadLane_29[20] & output_20_ready_0
    | requestReadLane_29[21] & output_21_ready_0 | requestReadLane_29[22] & output_22_ready_0 | requestReadLane_29[23] & output_23_ready_0 | requestReadLane_29[24] & output_24_ready_0 | requestReadLane_29[25] & output_25_ready_0
    | requestReadLane_29[26] & output_26_ready_0 | requestReadLane_29[27] & output_27_ready_0 | requestReadLane_29[28] & output_28_ready_0 | requestReadLane_29[29] & output_29_ready_0 | requestReadLane_29[30] & output_30_ready_0
    | requestReadLane_29[31] & output_31_ready_0;
  wire        input_29_ready_0 = free_29 & outReady_29;
  wire [31:0] inputSelect1H_29 = input_29_valid_0 & free_29 ? requestReadLane_29 : 32'h0;
  wire [31:0] _GEN_27 = _GEN_26 | inputSelect1H_29;
  wire [31:0] requestReadLane_30 = 32'h1 << input_30_bits_readLane_0;
  wire        free_30 = |(requestReadLane_30 & ~_GEN_27);
  wire        outReady_30 =
    requestReadLane_30[0] & output_0_ready_0 | requestReadLane_30[1] & output_1_ready_0 | requestReadLane_30[2] & output_2_ready_0 | requestReadLane_30[3] & output_3_ready_0 | requestReadLane_30[4] & output_4_ready_0 | requestReadLane_30[5]
    & output_5_ready_0 | requestReadLane_30[6] & output_6_ready_0 | requestReadLane_30[7] & output_7_ready_0 | requestReadLane_30[8] & output_8_ready_0 | requestReadLane_30[9] & output_9_ready_0 | requestReadLane_30[10] & output_10_ready_0
    | requestReadLane_30[11] & output_11_ready_0 | requestReadLane_30[12] & output_12_ready_0 | requestReadLane_30[13] & output_13_ready_0 | requestReadLane_30[14] & output_14_ready_0 | requestReadLane_30[15] & output_15_ready_0
    | requestReadLane_30[16] & output_16_ready_0 | requestReadLane_30[17] & output_17_ready_0 | requestReadLane_30[18] & output_18_ready_0 | requestReadLane_30[19] & output_19_ready_0 | requestReadLane_30[20] & output_20_ready_0
    | requestReadLane_30[21] & output_21_ready_0 | requestReadLane_30[22] & output_22_ready_0 | requestReadLane_30[23] & output_23_ready_0 | requestReadLane_30[24] & output_24_ready_0 | requestReadLane_30[25] & output_25_ready_0
    | requestReadLane_30[26] & output_26_ready_0 | requestReadLane_30[27] & output_27_ready_0 | requestReadLane_30[28] & output_28_ready_0 | requestReadLane_30[29] & output_29_ready_0 | requestReadLane_30[30] & output_30_ready_0
    | requestReadLane_30[31] & output_31_ready_0;
  wire        input_30_ready_0 = free_30 & outReady_30;
  wire [31:0] inputSelect1H_30 = input_30_valid_0 & free_30 ? requestReadLane_30 : 32'h0;
  wire [31:0] requestReadLane_31 = 32'h1 << input_31_bits_readLane_0;
  wire        free_31 = |(requestReadLane_31 & ~(_GEN_27 | inputSelect1H_30));
  wire        outReady_31 =
    requestReadLane_31[0] & output_0_ready_0 | requestReadLane_31[1] & output_1_ready_0 | requestReadLane_31[2] & output_2_ready_0 | requestReadLane_31[3] & output_3_ready_0 | requestReadLane_31[4] & output_4_ready_0 | requestReadLane_31[5]
    & output_5_ready_0 | requestReadLane_31[6] & output_6_ready_0 | requestReadLane_31[7] & output_7_ready_0 | requestReadLane_31[8] & output_8_ready_0 | requestReadLane_31[9] & output_9_ready_0 | requestReadLane_31[10] & output_10_ready_0
    | requestReadLane_31[11] & output_11_ready_0 | requestReadLane_31[12] & output_12_ready_0 | requestReadLane_31[13] & output_13_ready_0 | requestReadLane_31[14] & output_14_ready_0 | requestReadLane_31[15] & output_15_ready_0
    | requestReadLane_31[16] & output_16_ready_0 | requestReadLane_31[17] & output_17_ready_0 | requestReadLane_31[18] & output_18_ready_0 | requestReadLane_31[19] & output_19_ready_0 | requestReadLane_31[20] & output_20_ready_0
    | requestReadLane_31[21] & output_21_ready_0 | requestReadLane_31[22] & output_22_ready_0 | requestReadLane_31[23] & output_23_ready_0 | requestReadLane_31[24] & output_24_ready_0 | requestReadLane_31[25] & output_25_ready_0
    | requestReadLane_31[26] & output_26_ready_0 | requestReadLane_31[27] & output_27_ready_0 | requestReadLane_31[28] & output_28_ready_0 | requestReadLane_31[29] & output_29_ready_0 | requestReadLane_31[30] & output_30_ready_0
    | requestReadLane_31[31] & output_31_ready_0;
  wire        input_31_ready_0 = free_31 & outReady_31;
  wire [31:0] inputSelect1H_31 = input_31_valid_0 & free_31 ? requestReadLane_31 : 32'h0;
  wire [1:0]  tryToRead_lo_lo_lo_lo = {inputSelect1H_1[0], inputSelect1H_0[0]};
  wire [1:0]  tryToRead_lo_lo_lo_hi = {inputSelect1H_3[0], inputSelect1H_2[0]};
  wire [3:0]  tryToRead_lo_lo_lo = {tryToRead_lo_lo_lo_hi, tryToRead_lo_lo_lo_lo};
  wire [1:0]  tryToRead_lo_lo_hi_lo = {inputSelect1H_5[0], inputSelect1H_4[0]};
  wire [1:0]  tryToRead_lo_lo_hi_hi = {inputSelect1H_7[0], inputSelect1H_6[0]};
  wire [3:0]  tryToRead_lo_lo_hi = {tryToRead_lo_lo_hi_hi, tryToRead_lo_lo_hi_lo};
  wire [7:0]  tryToRead_lo_lo = {tryToRead_lo_lo_hi, tryToRead_lo_lo_lo};
  wire [1:0]  tryToRead_lo_hi_lo_lo = {inputSelect1H_9[0], inputSelect1H_8[0]};
  wire [1:0]  tryToRead_lo_hi_lo_hi = {inputSelect1H_11[0], inputSelect1H_10[0]};
  wire [3:0]  tryToRead_lo_hi_lo = {tryToRead_lo_hi_lo_hi, tryToRead_lo_hi_lo_lo};
  wire [1:0]  tryToRead_lo_hi_hi_lo = {inputSelect1H_13[0], inputSelect1H_12[0]};
  wire [1:0]  tryToRead_lo_hi_hi_hi = {inputSelect1H_15[0], inputSelect1H_14[0]};
  wire [3:0]  tryToRead_lo_hi_hi = {tryToRead_lo_hi_hi_hi, tryToRead_lo_hi_hi_lo};
  wire [7:0]  tryToRead_lo_hi = {tryToRead_lo_hi_hi, tryToRead_lo_hi_lo};
  wire [15:0] tryToRead_lo = {tryToRead_lo_hi, tryToRead_lo_lo};
  wire [1:0]  tryToRead_hi_lo_lo_lo = {inputSelect1H_17[0], inputSelect1H_16[0]};
  wire [1:0]  tryToRead_hi_lo_lo_hi = {inputSelect1H_19[0], inputSelect1H_18[0]};
  wire [3:0]  tryToRead_hi_lo_lo = {tryToRead_hi_lo_lo_hi, tryToRead_hi_lo_lo_lo};
  wire [1:0]  tryToRead_hi_lo_hi_lo = {inputSelect1H_21[0], inputSelect1H_20[0]};
  wire [1:0]  tryToRead_hi_lo_hi_hi = {inputSelect1H_23[0], inputSelect1H_22[0]};
  wire [3:0]  tryToRead_hi_lo_hi = {tryToRead_hi_lo_hi_hi, tryToRead_hi_lo_hi_lo};
  wire [7:0]  tryToRead_hi_lo = {tryToRead_hi_lo_hi, tryToRead_hi_lo_lo};
  wire [1:0]  tryToRead_hi_hi_lo_lo = {inputSelect1H_25[0], inputSelect1H_24[0]};
  wire [1:0]  tryToRead_hi_hi_lo_hi = {inputSelect1H_27[0], inputSelect1H_26[0]};
  wire [3:0]  tryToRead_hi_hi_lo = {tryToRead_hi_hi_lo_hi, tryToRead_hi_hi_lo_lo};
  wire [1:0]  tryToRead_hi_hi_hi_lo = {inputSelect1H_29[0], inputSelect1H_28[0]};
  wire [1:0]  tryToRead_hi_hi_hi_hi = {inputSelect1H_31[0], inputSelect1H_30[0]};
  wire [3:0]  tryToRead_hi_hi_hi = {tryToRead_hi_hi_hi_hi, tryToRead_hi_hi_hi_lo};
  wire [7:0]  tryToRead_hi_hi = {tryToRead_hi_hi_hi, tryToRead_hi_hi_lo};
  wire [15:0] tryToRead_hi = {tryToRead_hi_hi, tryToRead_hi_lo};
  wire [31:0] tryToRead = {tryToRead_hi, tryToRead_lo};
  wire        output_0_valid_0 = |tryToRead;
  wire [4:0]  output_0_bits_vs_0 = selectReq_bits_vs;
  wire        output_0_bits_offset_0 = selectReq_bits_offset;
  wire [4:0]  output_0_bits_writeIndex_0 = selectReq_bits_requestIndex;
  wire [1:0]  output_0_bits_dataOffset_0 = selectReq_bits_dataOffset;
  assign selectReq_bits_dataOffset =
    (tryToRead[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_bits_requestIndex =
    {4'h0, tryToRead[1]} | {3'h0, tryToRead[2], 1'h0} | (tryToRead[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead[4], 2'h0} | (tryToRead[5] ? 5'h5 : 5'h0) | (tryToRead[6] ? 5'h6 : 5'h0) | (tryToRead[7] ? 5'h7 : 5'h0) | {1'h0, tryToRead[8], 3'h0}
    | (tryToRead[9] ? 5'h9 : 5'h0) | (tryToRead[10] ? 5'hA : 5'h0) | (tryToRead[11] ? 5'hB : 5'h0) | (tryToRead[12] ? 5'hC : 5'h0) | (tryToRead[13] ? 5'hD : 5'h0) | (tryToRead[14] ? 5'hE : 5'h0) | (tryToRead[15] ? 5'hF : 5'h0)
    | {tryToRead[16], 4'h0} | (tryToRead[17] ? 5'h11 : 5'h0) | (tryToRead[18] ? 5'h12 : 5'h0) | (tryToRead[19] ? 5'h13 : 5'h0) | (tryToRead[20] ? 5'h14 : 5'h0) | (tryToRead[21] ? 5'h15 : 5'h0) | (tryToRead[22] ? 5'h16 : 5'h0)
    | (tryToRead[23] ? 5'h17 : 5'h0) | (tryToRead[24] ? 5'h18 : 5'h0) | (tryToRead[25] ? 5'h19 : 5'h0) | (tryToRead[26] ? 5'h1A : 5'h0) | (tryToRead[27] ? 5'h1B : 5'h0) | (tryToRead[28] ? 5'h1C : 5'h0) | (tryToRead[29] ? 5'h1D : 5'h0)
    | (tryToRead[30] ? 5'h1E : 5'h0) | {5{tryToRead[31]}};
  wire [4:0]  selectReq_bits_readLane =
    (tryToRead[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_bits_offset =
    tryToRead[0] & input_0_bits_offset_0 | tryToRead[1] & input_1_bits_offset_0 | tryToRead[2] & input_2_bits_offset_0 | tryToRead[3] & input_3_bits_offset_0 | tryToRead[4] & input_4_bits_offset_0 | tryToRead[5] & input_5_bits_offset_0
    | tryToRead[6] & input_6_bits_offset_0 | tryToRead[7] & input_7_bits_offset_0 | tryToRead[8] & input_8_bits_offset_0 | tryToRead[9] & input_9_bits_offset_0 | tryToRead[10] & input_10_bits_offset_0 | tryToRead[11]
    & input_11_bits_offset_0 | tryToRead[12] & input_12_bits_offset_0 | tryToRead[13] & input_13_bits_offset_0 | tryToRead[14] & input_14_bits_offset_0 | tryToRead[15] & input_15_bits_offset_0 | tryToRead[16] & input_16_bits_offset_0
    | tryToRead[17] & input_17_bits_offset_0 | tryToRead[18] & input_18_bits_offset_0 | tryToRead[19] & input_19_bits_offset_0 | tryToRead[20] & input_20_bits_offset_0 | tryToRead[21] & input_21_bits_offset_0 | tryToRead[22]
    & input_22_bits_offset_0 | tryToRead[23] & input_23_bits_offset_0 | tryToRead[24] & input_24_bits_offset_0 | tryToRead[25] & input_25_bits_offset_0 | tryToRead[26] & input_26_bits_offset_0 | tryToRead[27] & input_27_bits_offset_0
    | tryToRead[28] & input_28_bits_offset_0 | tryToRead[29] & input_29_bits_offset_0 | tryToRead[30] & input_30_bits_offset_0 | tryToRead[31] & input_31_bits_offset_0;
  assign selectReq_bits_vs =
    (tryToRead[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead[13] ? input_13_bits_vs_0 : 5'h0) | (tryToRead[14] ? input_14_bits_vs_0 : 5'h0)
    | (tryToRead[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead[17] ? input_17_bits_vs_0 : 5'h0) | (tryToRead[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead[19] ? input_19_bits_vs_0 : 5'h0)
    | (tryToRead[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead[21] ? input_21_bits_vs_0 : 5'h0) | (tryToRead[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead[24] ? input_24_bits_vs_0 : 5'h0)
    | (tryToRead[25] ? input_25_bits_vs_0 : 5'h0) | (tryToRead[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_valid =
    tryToRead[0] & input_0_valid_0 | tryToRead[1] & input_1_valid_0 | tryToRead[2] & input_2_valid_0 | tryToRead[3] & input_3_valid_0 | tryToRead[4] & input_4_valid_0 | tryToRead[5] & input_5_valid_0 | tryToRead[6] & input_6_valid_0
    | tryToRead[7] & input_7_valid_0 | tryToRead[8] & input_8_valid_0 | tryToRead[9] & input_9_valid_0 | tryToRead[10] & input_10_valid_0 | tryToRead[11] & input_11_valid_0 | tryToRead[12] & input_12_valid_0 | tryToRead[13]
    & input_13_valid_0 | tryToRead[14] & input_14_valid_0 | tryToRead[15] & input_15_valid_0 | tryToRead[16] & input_16_valid_0 | tryToRead[17] & input_17_valid_0 | tryToRead[18] & input_18_valid_0 | tryToRead[19] & input_19_valid_0
    | tryToRead[20] & input_20_valid_0 | tryToRead[21] & input_21_valid_0 | tryToRead[22] & input_22_valid_0 | tryToRead[23] & input_23_valid_0 | tryToRead[24] & input_24_valid_0 | tryToRead[25] & input_25_valid_0 | tryToRead[26]
    & input_26_valid_0 | tryToRead[27] & input_27_valid_0 | tryToRead[28] & input_28_valid_0 | tryToRead[29] & input_29_valid_0 | tryToRead[30] & input_30_valid_0 | tryToRead[31] & input_31_valid_0;
  wire        selectReq_ready =
    tryToRead[0] & input_0_ready_0 | tryToRead[1] & input_1_ready_0 | tryToRead[2] & input_2_ready_0 | tryToRead[3] & input_3_ready_0 | tryToRead[4] & input_4_ready_0 | tryToRead[5] & input_5_ready_0 | tryToRead[6] & input_6_ready_0
    | tryToRead[7] & input_7_ready_0 | tryToRead[8] & input_8_ready_0 | tryToRead[9] & input_9_ready_0 | tryToRead[10] & input_10_ready_0 | tryToRead[11] & input_11_ready_0 | tryToRead[12] & input_12_ready_0 | tryToRead[13]
    & input_13_ready_0 | tryToRead[14] & input_14_ready_0 | tryToRead[15] & input_15_ready_0 | tryToRead[16] & input_16_ready_0 | tryToRead[17] & input_17_ready_0 | tryToRead[18] & input_18_ready_0 | tryToRead[19] & input_19_ready_0
    | tryToRead[20] & input_20_ready_0 | tryToRead[21] & input_21_ready_0 | tryToRead[22] & input_22_ready_0 | tryToRead[23] & input_23_ready_0 | tryToRead[24] & input_24_ready_0 | tryToRead[25] & input_25_ready_0 | tryToRead[26]
    & input_26_ready_0 | tryToRead[27] & input_27_ready_0 | tryToRead[28] & input_28_ready_0 | tryToRead[29] & input_29_ready_0 | tryToRead[30] & input_30_ready_0 | tryToRead[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_1 = {inputSelect1H_1[1], inputSelect1H_0[1]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_1 = {inputSelect1H_3[1], inputSelect1H_2[1]};
  wire [3:0]  tryToRead_lo_lo_lo_1 = {tryToRead_lo_lo_lo_hi_1, tryToRead_lo_lo_lo_lo_1};
  wire [1:0]  tryToRead_lo_lo_hi_lo_1 = {inputSelect1H_5[1], inputSelect1H_4[1]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_1 = {inputSelect1H_7[1], inputSelect1H_6[1]};
  wire [3:0]  tryToRead_lo_lo_hi_1 = {tryToRead_lo_lo_hi_hi_1, tryToRead_lo_lo_hi_lo_1};
  wire [7:0]  tryToRead_lo_lo_1 = {tryToRead_lo_lo_hi_1, tryToRead_lo_lo_lo_1};
  wire [1:0]  tryToRead_lo_hi_lo_lo_1 = {inputSelect1H_9[1], inputSelect1H_8[1]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_1 = {inputSelect1H_11[1], inputSelect1H_10[1]};
  wire [3:0]  tryToRead_lo_hi_lo_1 = {tryToRead_lo_hi_lo_hi_1, tryToRead_lo_hi_lo_lo_1};
  wire [1:0]  tryToRead_lo_hi_hi_lo_1 = {inputSelect1H_13[1], inputSelect1H_12[1]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_1 = {inputSelect1H_15[1], inputSelect1H_14[1]};
  wire [3:0]  tryToRead_lo_hi_hi_1 = {tryToRead_lo_hi_hi_hi_1, tryToRead_lo_hi_hi_lo_1};
  wire [7:0]  tryToRead_lo_hi_1 = {tryToRead_lo_hi_hi_1, tryToRead_lo_hi_lo_1};
  wire [15:0] tryToRead_lo_1 = {tryToRead_lo_hi_1, tryToRead_lo_lo_1};
  wire [1:0]  tryToRead_hi_lo_lo_lo_1 = {inputSelect1H_17[1], inputSelect1H_16[1]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_1 = {inputSelect1H_19[1], inputSelect1H_18[1]};
  wire [3:0]  tryToRead_hi_lo_lo_1 = {tryToRead_hi_lo_lo_hi_1, tryToRead_hi_lo_lo_lo_1};
  wire [1:0]  tryToRead_hi_lo_hi_lo_1 = {inputSelect1H_21[1], inputSelect1H_20[1]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_1 = {inputSelect1H_23[1], inputSelect1H_22[1]};
  wire [3:0]  tryToRead_hi_lo_hi_1 = {tryToRead_hi_lo_hi_hi_1, tryToRead_hi_lo_hi_lo_1};
  wire [7:0]  tryToRead_hi_lo_1 = {tryToRead_hi_lo_hi_1, tryToRead_hi_lo_lo_1};
  wire [1:0]  tryToRead_hi_hi_lo_lo_1 = {inputSelect1H_25[1], inputSelect1H_24[1]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_1 = {inputSelect1H_27[1], inputSelect1H_26[1]};
  wire [3:0]  tryToRead_hi_hi_lo_1 = {tryToRead_hi_hi_lo_hi_1, tryToRead_hi_hi_lo_lo_1};
  wire [1:0]  tryToRead_hi_hi_hi_lo_1 = {inputSelect1H_29[1], inputSelect1H_28[1]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_1 = {inputSelect1H_31[1], inputSelect1H_30[1]};
  wire [3:0]  tryToRead_hi_hi_hi_1 = {tryToRead_hi_hi_hi_hi_1, tryToRead_hi_hi_hi_lo_1};
  wire [7:0]  tryToRead_hi_hi_1 = {tryToRead_hi_hi_hi_1, tryToRead_hi_hi_lo_1};
  wire [15:0] tryToRead_hi_1 = {tryToRead_hi_hi_1, tryToRead_hi_lo_1};
  wire [31:0] tryToRead_1 = {tryToRead_hi_1, tryToRead_lo_1};
  wire        output_1_valid_0 = |tryToRead_1;
  wire [4:0]  output_1_bits_vs_0 = selectReq_1_bits_vs;
  wire        output_1_bits_offset_0 = selectReq_1_bits_offset;
  wire [4:0]  output_1_bits_writeIndex_0 = selectReq_1_bits_requestIndex;
  wire [1:0]  output_1_bits_dataOffset_0 = selectReq_1_bits_dataOffset;
  assign selectReq_1_bits_dataOffset =
    (tryToRead_1[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_1[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_1[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_1[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_1[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_1[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_1[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_1[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_1[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_1[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_1[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_1[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_1[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_1[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_1[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_1[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_1[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_1[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_1[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_1[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_1[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_1[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_1[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_1[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_1[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_1_bits_requestIndex =
    {4'h0, tryToRead_1[1]} | {3'h0, tryToRead_1[2], 1'h0} | (tryToRead_1[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_1[4], 2'h0} | (tryToRead_1[5] ? 5'h5 : 5'h0) | (tryToRead_1[6] ? 5'h6 : 5'h0) | (tryToRead_1[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_1[8], 3'h0} | (tryToRead_1[9] ? 5'h9 : 5'h0) | (tryToRead_1[10] ? 5'hA : 5'h0) | (tryToRead_1[11] ? 5'hB : 5'h0) | (tryToRead_1[12] ? 5'hC : 5'h0) | (tryToRead_1[13] ? 5'hD : 5'h0) | (tryToRead_1[14] ? 5'hE : 5'h0)
    | (tryToRead_1[15] ? 5'hF : 5'h0) | {tryToRead_1[16], 4'h0} | (tryToRead_1[17] ? 5'h11 : 5'h0) | (tryToRead_1[18] ? 5'h12 : 5'h0) | (tryToRead_1[19] ? 5'h13 : 5'h0) | (tryToRead_1[20] ? 5'h14 : 5'h0) | (tryToRead_1[21] ? 5'h15 : 5'h0)
    | (tryToRead_1[22] ? 5'h16 : 5'h0) | (tryToRead_1[23] ? 5'h17 : 5'h0) | (tryToRead_1[24] ? 5'h18 : 5'h0) | (tryToRead_1[25] ? 5'h19 : 5'h0) | (tryToRead_1[26] ? 5'h1A : 5'h0) | (tryToRead_1[27] ? 5'h1B : 5'h0)
    | (tryToRead_1[28] ? 5'h1C : 5'h0) | (tryToRead_1[29] ? 5'h1D : 5'h0) | (tryToRead_1[30] ? 5'h1E : 5'h0) | {5{tryToRead_1[31]}};
  wire [4:0]  selectReq_1_bits_readLane =
    (tryToRead_1[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_1[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_1[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_1[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_1[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_1[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_1[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_1[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_1[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_1[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_1[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_1[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_1[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_1[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_1[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_1[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_1[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_1[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_1[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_1[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_1[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_1[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_1[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_1[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_1[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_1[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_1[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_1[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_1[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_1[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_1[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_1[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_1_bits_offset =
    tryToRead_1[0] & input_0_bits_offset_0 | tryToRead_1[1] & input_1_bits_offset_0 | tryToRead_1[2] & input_2_bits_offset_0 | tryToRead_1[3] & input_3_bits_offset_0 | tryToRead_1[4] & input_4_bits_offset_0 | tryToRead_1[5]
    & input_5_bits_offset_0 | tryToRead_1[6] & input_6_bits_offset_0 | tryToRead_1[7] & input_7_bits_offset_0 | tryToRead_1[8] & input_8_bits_offset_0 | tryToRead_1[9] & input_9_bits_offset_0 | tryToRead_1[10] & input_10_bits_offset_0
    | tryToRead_1[11] & input_11_bits_offset_0 | tryToRead_1[12] & input_12_bits_offset_0 | tryToRead_1[13] & input_13_bits_offset_0 | tryToRead_1[14] & input_14_bits_offset_0 | tryToRead_1[15] & input_15_bits_offset_0 | tryToRead_1[16]
    & input_16_bits_offset_0 | tryToRead_1[17] & input_17_bits_offset_0 | tryToRead_1[18] & input_18_bits_offset_0 | tryToRead_1[19] & input_19_bits_offset_0 | tryToRead_1[20] & input_20_bits_offset_0 | tryToRead_1[21]
    & input_21_bits_offset_0 | tryToRead_1[22] & input_22_bits_offset_0 | tryToRead_1[23] & input_23_bits_offset_0 | tryToRead_1[24] & input_24_bits_offset_0 | tryToRead_1[25] & input_25_bits_offset_0 | tryToRead_1[26]
    & input_26_bits_offset_0 | tryToRead_1[27] & input_27_bits_offset_0 | tryToRead_1[28] & input_28_bits_offset_0 | tryToRead_1[29] & input_29_bits_offset_0 | tryToRead_1[30] & input_30_bits_offset_0 | tryToRead_1[31]
    & input_31_bits_offset_0;
  assign selectReq_1_bits_vs =
    (tryToRead_1[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_1[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_1[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_1[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_1[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_1[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_1[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_1[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_1[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_1[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_1[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_1[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_1[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_1[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_1[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_1[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_1[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_1[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_1[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_1[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_1[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_1[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_1[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_1[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_1[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_1[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_1[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_1[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_1[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_1[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_1[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_1[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_1_valid =
    tryToRead_1[0] & input_0_valid_0 | tryToRead_1[1] & input_1_valid_0 | tryToRead_1[2] & input_2_valid_0 | tryToRead_1[3] & input_3_valid_0 | tryToRead_1[4] & input_4_valid_0 | tryToRead_1[5] & input_5_valid_0 | tryToRead_1[6]
    & input_6_valid_0 | tryToRead_1[7] & input_7_valid_0 | tryToRead_1[8] & input_8_valid_0 | tryToRead_1[9] & input_9_valid_0 | tryToRead_1[10] & input_10_valid_0 | tryToRead_1[11] & input_11_valid_0 | tryToRead_1[12] & input_12_valid_0
    | tryToRead_1[13] & input_13_valid_0 | tryToRead_1[14] & input_14_valid_0 | tryToRead_1[15] & input_15_valid_0 | tryToRead_1[16] & input_16_valid_0 | tryToRead_1[17] & input_17_valid_0 | tryToRead_1[18] & input_18_valid_0
    | tryToRead_1[19] & input_19_valid_0 | tryToRead_1[20] & input_20_valid_0 | tryToRead_1[21] & input_21_valid_0 | tryToRead_1[22] & input_22_valid_0 | tryToRead_1[23] & input_23_valid_0 | tryToRead_1[24] & input_24_valid_0
    | tryToRead_1[25] & input_25_valid_0 | tryToRead_1[26] & input_26_valid_0 | tryToRead_1[27] & input_27_valid_0 | tryToRead_1[28] & input_28_valid_0 | tryToRead_1[29] & input_29_valid_0 | tryToRead_1[30] & input_30_valid_0
    | tryToRead_1[31] & input_31_valid_0;
  wire        selectReq_1_ready =
    tryToRead_1[0] & input_0_ready_0 | tryToRead_1[1] & input_1_ready_0 | tryToRead_1[2] & input_2_ready_0 | tryToRead_1[3] & input_3_ready_0 | tryToRead_1[4] & input_4_ready_0 | tryToRead_1[5] & input_5_ready_0 | tryToRead_1[6]
    & input_6_ready_0 | tryToRead_1[7] & input_7_ready_0 | tryToRead_1[8] & input_8_ready_0 | tryToRead_1[9] & input_9_ready_0 | tryToRead_1[10] & input_10_ready_0 | tryToRead_1[11] & input_11_ready_0 | tryToRead_1[12] & input_12_ready_0
    | tryToRead_1[13] & input_13_ready_0 | tryToRead_1[14] & input_14_ready_0 | tryToRead_1[15] & input_15_ready_0 | tryToRead_1[16] & input_16_ready_0 | tryToRead_1[17] & input_17_ready_0 | tryToRead_1[18] & input_18_ready_0
    | tryToRead_1[19] & input_19_ready_0 | tryToRead_1[20] & input_20_ready_0 | tryToRead_1[21] & input_21_ready_0 | tryToRead_1[22] & input_22_ready_0 | tryToRead_1[23] & input_23_ready_0 | tryToRead_1[24] & input_24_ready_0
    | tryToRead_1[25] & input_25_ready_0 | tryToRead_1[26] & input_26_ready_0 | tryToRead_1[27] & input_27_ready_0 | tryToRead_1[28] & input_28_ready_0 | tryToRead_1[29] & input_29_ready_0 | tryToRead_1[30] & input_30_ready_0
    | tryToRead_1[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_2 = {inputSelect1H_1[2], inputSelect1H_0[2]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_2 = {inputSelect1H_3[2], inputSelect1H_2[2]};
  wire [3:0]  tryToRead_lo_lo_lo_2 = {tryToRead_lo_lo_lo_hi_2, tryToRead_lo_lo_lo_lo_2};
  wire [1:0]  tryToRead_lo_lo_hi_lo_2 = {inputSelect1H_5[2], inputSelect1H_4[2]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_2 = {inputSelect1H_7[2], inputSelect1H_6[2]};
  wire [3:0]  tryToRead_lo_lo_hi_2 = {tryToRead_lo_lo_hi_hi_2, tryToRead_lo_lo_hi_lo_2};
  wire [7:0]  tryToRead_lo_lo_2 = {tryToRead_lo_lo_hi_2, tryToRead_lo_lo_lo_2};
  wire [1:0]  tryToRead_lo_hi_lo_lo_2 = {inputSelect1H_9[2], inputSelect1H_8[2]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_2 = {inputSelect1H_11[2], inputSelect1H_10[2]};
  wire [3:0]  tryToRead_lo_hi_lo_2 = {tryToRead_lo_hi_lo_hi_2, tryToRead_lo_hi_lo_lo_2};
  wire [1:0]  tryToRead_lo_hi_hi_lo_2 = {inputSelect1H_13[2], inputSelect1H_12[2]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_2 = {inputSelect1H_15[2], inputSelect1H_14[2]};
  wire [3:0]  tryToRead_lo_hi_hi_2 = {tryToRead_lo_hi_hi_hi_2, tryToRead_lo_hi_hi_lo_2};
  wire [7:0]  tryToRead_lo_hi_2 = {tryToRead_lo_hi_hi_2, tryToRead_lo_hi_lo_2};
  wire [15:0] tryToRead_lo_2 = {tryToRead_lo_hi_2, tryToRead_lo_lo_2};
  wire [1:0]  tryToRead_hi_lo_lo_lo_2 = {inputSelect1H_17[2], inputSelect1H_16[2]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_2 = {inputSelect1H_19[2], inputSelect1H_18[2]};
  wire [3:0]  tryToRead_hi_lo_lo_2 = {tryToRead_hi_lo_lo_hi_2, tryToRead_hi_lo_lo_lo_2};
  wire [1:0]  tryToRead_hi_lo_hi_lo_2 = {inputSelect1H_21[2], inputSelect1H_20[2]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_2 = {inputSelect1H_23[2], inputSelect1H_22[2]};
  wire [3:0]  tryToRead_hi_lo_hi_2 = {tryToRead_hi_lo_hi_hi_2, tryToRead_hi_lo_hi_lo_2};
  wire [7:0]  tryToRead_hi_lo_2 = {tryToRead_hi_lo_hi_2, tryToRead_hi_lo_lo_2};
  wire [1:0]  tryToRead_hi_hi_lo_lo_2 = {inputSelect1H_25[2], inputSelect1H_24[2]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_2 = {inputSelect1H_27[2], inputSelect1H_26[2]};
  wire [3:0]  tryToRead_hi_hi_lo_2 = {tryToRead_hi_hi_lo_hi_2, tryToRead_hi_hi_lo_lo_2};
  wire [1:0]  tryToRead_hi_hi_hi_lo_2 = {inputSelect1H_29[2], inputSelect1H_28[2]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_2 = {inputSelect1H_31[2], inputSelect1H_30[2]};
  wire [3:0]  tryToRead_hi_hi_hi_2 = {tryToRead_hi_hi_hi_hi_2, tryToRead_hi_hi_hi_lo_2};
  wire [7:0]  tryToRead_hi_hi_2 = {tryToRead_hi_hi_hi_2, tryToRead_hi_hi_lo_2};
  wire [15:0] tryToRead_hi_2 = {tryToRead_hi_hi_2, tryToRead_hi_lo_2};
  wire [31:0] tryToRead_2 = {tryToRead_hi_2, tryToRead_lo_2};
  wire        output_2_valid_0 = |tryToRead_2;
  wire [4:0]  output_2_bits_vs_0 = selectReq_2_bits_vs;
  wire        output_2_bits_offset_0 = selectReq_2_bits_offset;
  wire [4:0]  output_2_bits_writeIndex_0 = selectReq_2_bits_requestIndex;
  wire [1:0]  output_2_bits_dataOffset_0 = selectReq_2_bits_dataOffset;
  assign selectReq_2_bits_dataOffset =
    (tryToRead_2[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_2[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_2[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_2[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_2[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_2[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_2[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_2[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_2[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_2[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_2[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_2[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_2[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_2[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_2[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_2[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_2[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_2[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_2[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_2[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_2[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_2[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_2[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_2[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_2[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_2_bits_requestIndex =
    {4'h0, tryToRead_2[1]} | {3'h0, tryToRead_2[2], 1'h0} | (tryToRead_2[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_2[4], 2'h0} | (tryToRead_2[5] ? 5'h5 : 5'h0) | (tryToRead_2[6] ? 5'h6 : 5'h0) | (tryToRead_2[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_2[8], 3'h0} | (tryToRead_2[9] ? 5'h9 : 5'h0) | (tryToRead_2[10] ? 5'hA : 5'h0) | (tryToRead_2[11] ? 5'hB : 5'h0) | (tryToRead_2[12] ? 5'hC : 5'h0) | (tryToRead_2[13] ? 5'hD : 5'h0) | (tryToRead_2[14] ? 5'hE : 5'h0)
    | (tryToRead_2[15] ? 5'hF : 5'h0) | {tryToRead_2[16], 4'h0} | (tryToRead_2[17] ? 5'h11 : 5'h0) | (tryToRead_2[18] ? 5'h12 : 5'h0) | (tryToRead_2[19] ? 5'h13 : 5'h0) | (tryToRead_2[20] ? 5'h14 : 5'h0) | (tryToRead_2[21] ? 5'h15 : 5'h0)
    | (tryToRead_2[22] ? 5'h16 : 5'h0) | (tryToRead_2[23] ? 5'h17 : 5'h0) | (tryToRead_2[24] ? 5'h18 : 5'h0) | (tryToRead_2[25] ? 5'h19 : 5'h0) | (tryToRead_2[26] ? 5'h1A : 5'h0) | (tryToRead_2[27] ? 5'h1B : 5'h0)
    | (tryToRead_2[28] ? 5'h1C : 5'h0) | (tryToRead_2[29] ? 5'h1D : 5'h0) | (tryToRead_2[30] ? 5'h1E : 5'h0) | {5{tryToRead_2[31]}};
  wire [4:0]  selectReq_2_bits_readLane =
    (tryToRead_2[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_2[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_2[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_2[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_2[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_2[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_2[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_2[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_2[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_2[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_2[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_2[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_2[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_2[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_2[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_2[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_2[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_2[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_2[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_2[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_2[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_2[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_2[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_2[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_2[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_2[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_2[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_2[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_2[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_2[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_2[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_2[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_2_bits_offset =
    tryToRead_2[0] & input_0_bits_offset_0 | tryToRead_2[1] & input_1_bits_offset_0 | tryToRead_2[2] & input_2_bits_offset_0 | tryToRead_2[3] & input_3_bits_offset_0 | tryToRead_2[4] & input_4_bits_offset_0 | tryToRead_2[5]
    & input_5_bits_offset_0 | tryToRead_2[6] & input_6_bits_offset_0 | tryToRead_2[7] & input_7_bits_offset_0 | tryToRead_2[8] & input_8_bits_offset_0 | tryToRead_2[9] & input_9_bits_offset_0 | tryToRead_2[10] & input_10_bits_offset_0
    | tryToRead_2[11] & input_11_bits_offset_0 | tryToRead_2[12] & input_12_bits_offset_0 | tryToRead_2[13] & input_13_bits_offset_0 | tryToRead_2[14] & input_14_bits_offset_0 | tryToRead_2[15] & input_15_bits_offset_0 | tryToRead_2[16]
    & input_16_bits_offset_0 | tryToRead_2[17] & input_17_bits_offset_0 | tryToRead_2[18] & input_18_bits_offset_0 | tryToRead_2[19] & input_19_bits_offset_0 | tryToRead_2[20] & input_20_bits_offset_0 | tryToRead_2[21]
    & input_21_bits_offset_0 | tryToRead_2[22] & input_22_bits_offset_0 | tryToRead_2[23] & input_23_bits_offset_0 | tryToRead_2[24] & input_24_bits_offset_0 | tryToRead_2[25] & input_25_bits_offset_0 | tryToRead_2[26]
    & input_26_bits_offset_0 | tryToRead_2[27] & input_27_bits_offset_0 | tryToRead_2[28] & input_28_bits_offset_0 | tryToRead_2[29] & input_29_bits_offset_0 | tryToRead_2[30] & input_30_bits_offset_0 | tryToRead_2[31]
    & input_31_bits_offset_0;
  assign selectReq_2_bits_vs =
    (tryToRead_2[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_2[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_2[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_2[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_2[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_2[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_2[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_2[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_2[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_2[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_2[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_2[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_2[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_2[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_2[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_2[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_2[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_2[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_2[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_2[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_2[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_2[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_2[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_2[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_2[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_2[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_2[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_2[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_2[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_2[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_2[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_2[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_2_valid =
    tryToRead_2[0] & input_0_valid_0 | tryToRead_2[1] & input_1_valid_0 | tryToRead_2[2] & input_2_valid_0 | tryToRead_2[3] & input_3_valid_0 | tryToRead_2[4] & input_4_valid_0 | tryToRead_2[5] & input_5_valid_0 | tryToRead_2[6]
    & input_6_valid_0 | tryToRead_2[7] & input_7_valid_0 | tryToRead_2[8] & input_8_valid_0 | tryToRead_2[9] & input_9_valid_0 | tryToRead_2[10] & input_10_valid_0 | tryToRead_2[11] & input_11_valid_0 | tryToRead_2[12] & input_12_valid_0
    | tryToRead_2[13] & input_13_valid_0 | tryToRead_2[14] & input_14_valid_0 | tryToRead_2[15] & input_15_valid_0 | tryToRead_2[16] & input_16_valid_0 | tryToRead_2[17] & input_17_valid_0 | tryToRead_2[18] & input_18_valid_0
    | tryToRead_2[19] & input_19_valid_0 | tryToRead_2[20] & input_20_valid_0 | tryToRead_2[21] & input_21_valid_0 | tryToRead_2[22] & input_22_valid_0 | tryToRead_2[23] & input_23_valid_0 | tryToRead_2[24] & input_24_valid_0
    | tryToRead_2[25] & input_25_valid_0 | tryToRead_2[26] & input_26_valid_0 | tryToRead_2[27] & input_27_valid_0 | tryToRead_2[28] & input_28_valid_0 | tryToRead_2[29] & input_29_valid_0 | tryToRead_2[30] & input_30_valid_0
    | tryToRead_2[31] & input_31_valid_0;
  wire        selectReq_2_ready =
    tryToRead_2[0] & input_0_ready_0 | tryToRead_2[1] & input_1_ready_0 | tryToRead_2[2] & input_2_ready_0 | tryToRead_2[3] & input_3_ready_0 | tryToRead_2[4] & input_4_ready_0 | tryToRead_2[5] & input_5_ready_0 | tryToRead_2[6]
    & input_6_ready_0 | tryToRead_2[7] & input_7_ready_0 | tryToRead_2[8] & input_8_ready_0 | tryToRead_2[9] & input_9_ready_0 | tryToRead_2[10] & input_10_ready_0 | tryToRead_2[11] & input_11_ready_0 | tryToRead_2[12] & input_12_ready_0
    | tryToRead_2[13] & input_13_ready_0 | tryToRead_2[14] & input_14_ready_0 | tryToRead_2[15] & input_15_ready_0 | tryToRead_2[16] & input_16_ready_0 | tryToRead_2[17] & input_17_ready_0 | tryToRead_2[18] & input_18_ready_0
    | tryToRead_2[19] & input_19_ready_0 | tryToRead_2[20] & input_20_ready_0 | tryToRead_2[21] & input_21_ready_0 | tryToRead_2[22] & input_22_ready_0 | tryToRead_2[23] & input_23_ready_0 | tryToRead_2[24] & input_24_ready_0
    | tryToRead_2[25] & input_25_ready_0 | tryToRead_2[26] & input_26_ready_0 | tryToRead_2[27] & input_27_ready_0 | tryToRead_2[28] & input_28_ready_0 | tryToRead_2[29] & input_29_ready_0 | tryToRead_2[30] & input_30_ready_0
    | tryToRead_2[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_3 = {inputSelect1H_1[3], inputSelect1H_0[3]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_3 = {inputSelect1H_3[3], inputSelect1H_2[3]};
  wire [3:0]  tryToRead_lo_lo_lo_3 = {tryToRead_lo_lo_lo_hi_3, tryToRead_lo_lo_lo_lo_3};
  wire [1:0]  tryToRead_lo_lo_hi_lo_3 = {inputSelect1H_5[3], inputSelect1H_4[3]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_3 = {inputSelect1H_7[3], inputSelect1H_6[3]};
  wire [3:0]  tryToRead_lo_lo_hi_3 = {tryToRead_lo_lo_hi_hi_3, tryToRead_lo_lo_hi_lo_3};
  wire [7:0]  tryToRead_lo_lo_3 = {tryToRead_lo_lo_hi_3, tryToRead_lo_lo_lo_3};
  wire [1:0]  tryToRead_lo_hi_lo_lo_3 = {inputSelect1H_9[3], inputSelect1H_8[3]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_3 = {inputSelect1H_11[3], inputSelect1H_10[3]};
  wire [3:0]  tryToRead_lo_hi_lo_3 = {tryToRead_lo_hi_lo_hi_3, tryToRead_lo_hi_lo_lo_3};
  wire [1:0]  tryToRead_lo_hi_hi_lo_3 = {inputSelect1H_13[3], inputSelect1H_12[3]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_3 = {inputSelect1H_15[3], inputSelect1H_14[3]};
  wire [3:0]  tryToRead_lo_hi_hi_3 = {tryToRead_lo_hi_hi_hi_3, tryToRead_lo_hi_hi_lo_3};
  wire [7:0]  tryToRead_lo_hi_3 = {tryToRead_lo_hi_hi_3, tryToRead_lo_hi_lo_3};
  wire [15:0] tryToRead_lo_3 = {tryToRead_lo_hi_3, tryToRead_lo_lo_3};
  wire [1:0]  tryToRead_hi_lo_lo_lo_3 = {inputSelect1H_17[3], inputSelect1H_16[3]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_3 = {inputSelect1H_19[3], inputSelect1H_18[3]};
  wire [3:0]  tryToRead_hi_lo_lo_3 = {tryToRead_hi_lo_lo_hi_3, tryToRead_hi_lo_lo_lo_3};
  wire [1:0]  tryToRead_hi_lo_hi_lo_3 = {inputSelect1H_21[3], inputSelect1H_20[3]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_3 = {inputSelect1H_23[3], inputSelect1H_22[3]};
  wire [3:0]  tryToRead_hi_lo_hi_3 = {tryToRead_hi_lo_hi_hi_3, tryToRead_hi_lo_hi_lo_3};
  wire [7:0]  tryToRead_hi_lo_3 = {tryToRead_hi_lo_hi_3, tryToRead_hi_lo_lo_3};
  wire [1:0]  tryToRead_hi_hi_lo_lo_3 = {inputSelect1H_25[3], inputSelect1H_24[3]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_3 = {inputSelect1H_27[3], inputSelect1H_26[3]};
  wire [3:0]  tryToRead_hi_hi_lo_3 = {tryToRead_hi_hi_lo_hi_3, tryToRead_hi_hi_lo_lo_3};
  wire [1:0]  tryToRead_hi_hi_hi_lo_3 = {inputSelect1H_29[3], inputSelect1H_28[3]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_3 = {inputSelect1H_31[3], inputSelect1H_30[3]};
  wire [3:0]  tryToRead_hi_hi_hi_3 = {tryToRead_hi_hi_hi_hi_3, tryToRead_hi_hi_hi_lo_3};
  wire [7:0]  tryToRead_hi_hi_3 = {tryToRead_hi_hi_hi_3, tryToRead_hi_hi_lo_3};
  wire [15:0] tryToRead_hi_3 = {tryToRead_hi_hi_3, tryToRead_hi_lo_3};
  wire [31:0] tryToRead_3 = {tryToRead_hi_3, tryToRead_lo_3};
  wire        output_3_valid_0 = |tryToRead_3;
  wire [4:0]  output_3_bits_vs_0 = selectReq_3_bits_vs;
  wire        output_3_bits_offset_0 = selectReq_3_bits_offset;
  wire [4:0]  output_3_bits_writeIndex_0 = selectReq_3_bits_requestIndex;
  wire [1:0]  output_3_bits_dataOffset_0 = selectReq_3_bits_dataOffset;
  assign selectReq_3_bits_dataOffset =
    (tryToRead_3[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_3[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_3[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_3[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_3[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_3[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_3[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_3[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_3[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_3[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_3[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_3[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_3[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_3[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_3[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_3[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_3[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_3[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_3[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_3[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_3[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_3[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_3[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_3[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_3[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_3_bits_requestIndex =
    {4'h0, tryToRead_3[1]} | {3'h0, tryToRead_3[2], 1'h0} | (tryToRead_3[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_3[4], 2'h0} | (tryToRead_3[5] ? 5'h5 : 5'h0) | (tryToRead_3[6] ? 5'h6 : 5'h0) | (tryToRead_3[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_3[8], 3'h0} | (tryToRead_3[9] ? 5'h9 : 5'h0) | (tryToRead_3[10] ? 5'hA : 5'h0) | (tryToRead_3[11] ? 5'hB : 5'h0) | (tryToRead_3[12] ? 5'hC : 5'h0) | (tryToRead_3[13] ? 5'hD : 5'h0) | (tryToRead_3[14] ? 5'hE : 5'h0)
    | (tryToRead_3[15] ? 5'hF : 5'h0) | {tryToRead_3[16], 4'h0} | (tryToRead_3[17] ? 5'h11 : 5'h0) | (tryToRead_3[18] ? 5'h12 : 5'h0) | (tryToRead_3[19] ? 5'h13 : 5'h0) | (tryToRead_3[20] ? 5'h14 : 5'h0) | (tryToRead_3[21] ? 5'h15 : 5'h0)
    | (tryToRead_3[22] ? 5'h16 : 5'h0) | (tryToRead_3[23] ? 5'h17 : 5'h0) | (tryToRead_3[24] ? 5'h18 : 5'h0) | (tryToRead_3[25] ? 5'h19 : 5'h0) | (tryToRead_3[26] ? 5'h1A : 5'h0) | (tryToRead_3[27] ? 5'h1B : 5'h0)
    | (tryToRead_3[28] ? 5'h1C : 5'h0) | (tryToRead_3[29] ? 5'h1D : 5'h0) | (tryToRead_3[30] ? 5'h1E : 5'h0) | {5{tryToRead_3[31]}};
  wire [4:0]  selectReq_3_bits_readLane =
    (tryToRead_3[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_3[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_3[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_3[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_3[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_3[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_3[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_3[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_3[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_3[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_3[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_3[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_3[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_3[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_3[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_3[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_3[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_3[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_3[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_3[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_3[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_3[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_3[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_3[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_3[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_3[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_3[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_3[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_3[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_3[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_3[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_3[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_3_bits_offset =
    tryToRead_3[0] & input_0_bits_offset_0 | tryToRead_3[1] & input_1_bits_offset_0 | tryToRead_3[2] & input_2_bits_offset_0 | tryToRead_3[3] & input_3_bits_offset_0 | tryToRead_3[4] & input_4_bits_offset_0 | tryToRead_3[5]
    & input_5_bits_offset_0 | tryToRead_3[6] & input_6_bits_offset_0 | tryToRead_3[7] & input_7_bits_offset_0 | tryToRead_3[8] & input_8_bits_offset_0 | tryToRead_3[9] & input_9_bits_offset_0 | tryToRead_3[10] & input_10_bits_offset_0
    | tryToRead_3[11] & input_11_bits_offset_0 | tryToRead_3[12] & input_12_bits_offset_0 | tryToRead_3[13] & input_13_bits_offset_0 | tryToRead_3[14] & input_14_bits_offset_0 | tryToRead_3[15] & input_15_bits_offset_0 | tryToRead_3[16]
    & input_16_bits_offset_0 | tryToRead_3[17] & input_17_bits_offset_0 | tryToRead_3[18] & input_18_bits_offset_0 | tryToRead_3[19] & input_19_bits_offset_0 | tryToRead_3[20] & input_20_bits_offset_0 | tryToRead_3[21]
    & input_21_bits_offset_0 | tryToRead_3[22] & input_22_bits_offset_0 | tryToRead_3[23] & input_23_bits_offset_0 | tryToRead_3[24] & input_24_bits_offset_0 | tryToRead_3[25] & input_25_bits_offset_0 | tryToRead_3[26]
    & input_26_bits_offset_0 | tryToRead_3[27] & input_27_bits_offset_0 | tryToRead_3[28] & input_28_bits_offset_0 | tryToRead_3[29] & input_29_bits_offset_0 | tryToRead_3[30] & input_30_bits_offset_0 | tryToRead_3[31]
    & input_31_bits_offset_0;
  assign selectReq_3_bits_vs =
    (tryToRead_3[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_3[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_3[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_3[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_3[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_3[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_3[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_3[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_3[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_3[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_3[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_3[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_3[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_3[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_3[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_3[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_3[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_3[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_3[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_3[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_3[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_3[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_3[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_3[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_3[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_3[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_3[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_3[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_3[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_3[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_3[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_3[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_3_valid =
    tryToRead_3[0] & input_0_valid_0 | tryToRead_3[1] & input_1_valid_0 | tryToRead_3[2] & input_2_valid_0 | tryToRead_3[3] & input_3_valid_0 | tryToRead_3[4] & input_4_valid_0 | tryToRead_3[5] & input_5_valid_0 | tryToRead_3[6]
    & input_6_valid_0 | tryToRead_3[7] & input_7_valid_0 | tryToRead_3[8] & input_8_valid_0 | tryToRead_3[9] & input_9_valid_0 | tryToRead_3[10] & input_10_valid_0 | tryToRead_3[11] & input_11_valid_0 | tryToRead_3[12] & input_12_valid_0
    | tryToRead_3[13] & input_13_valid_0 | tryToRead_3[14] & input_14_valid_0 | tryToRead_3[15] & input_15_valid_0 | tryToRead_3[16] & input_16_valid_0 | tryToRead_3[17] & input_17_valid_0 | tryToRead_3[18] & input_18_valid_0
    | tryToRead_3[19] & input_19_valid_0 | tryToRead_3[20] & input_20_valid_0 | tryToRead_3[21] & input_21_valid_0 | tryToRead_3[22] & input_22_valid_0 | tryToRead_3[23] & input_23_valid_0 | tryToRead_3[24] & input_24_valid_0
    | tryToRead_3[25] & input_25_valid_0 | tryToRead_3[26] & input_26_valid_0 | tryToRead_3[27] & input_27_valid_0 | tryToRead_3[28] & input_28_valid_0 | tryToRead_3[29] & input_29_valid_0 | tryToRead_3[30] & input_30_valid_0
    | tryToRead_3[31] & input_31_valid_0;
  wire        selectReq_3_ready =
    tryToRead_3[0] & input_0_ready_0 | tryToRead_3[1] & input_1_ready_0 | tryToRead_3[2] & input_2_ready_0 | tryToRead_3[3] & input_3_ready_0 | tryToRead_3[4] & input_4_ready_0 | tryToRead_3[5] & input_5_ready_0 | tryToRead_3[6]
    & input_6_ready_0 | tryToRead_3[7] & input_7_ready_0 | tryToRead_3[8] & input_8_ready_0 | tryToRead_3[9] & input_9_ready_0 | tryToRead_3[10] & input_10_ready_0 | tryToRead_3[11] & input_11_ready_0 | tryToRead_3[12] & input_12_ready_0
    | tryToRead_3[13] & input_13_ready_0 | tryToRead_3[14] & input_14_ready_0 | tryToRead_3[15] & input_15_ready_0 | tryToRead_3[16] & input_16_ready_0 | tryToRead_3[17] & input_17_ready_0 | tryToRead_3[18] & input_18_ready_0
    | tryToRead_3[19] & input_19_ready_0 | tryToRead_3[20] & input_20_ready_0 | tryToRead_3[21] & input_21_ready_0 | tryToRead_3[22] & input_22_ready_0 | tryToRead_3[23] & input_23_ready_0 | tryToRead_3[24] & input_24_ready_0
    | tryToRead_3[25] & input_25_ready_0 | tryToRead_3[26] & input_26_ready_0 | tryToRead_3[27] & input_27_ready_0 | tryToRead_3[28] & input_28_ready_0 | tryToRead_3[29] & input_29_ready_0 | tryToRead_3[30] & input_30_ready_0
    | tryToRead_3[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_4 = {inputSelect1H_1[4], inputSelect1H_0[4]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_4 = {inputSelect1H_3[4], inputSelect1H_2[4]};
  wire [3:0]  tryToRead_lo_lo_lo_4 = {tryToRead_lo_lo_lo_hi_4, tryToRead_lo_lo_lo_lo_4};
  wire [1:0]  tryToRead_lo_lo_hi_lo_4 = {inputSelect1H_5[4], inputSelect1H_4[4]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_4 = {inputSelect1H_7[4], inputSelect1H_6[4]};
  wire [3:0]  tryToRead_lo_lo_hi_4 = {tryToRead_lo_lo_hi_hi_4, tryToRead_lo_lo_hi_lo_4};
  wire [7:0]  tryToRead_lo_lo_4 = {tryToRead_lo_lo_hi_4, tryToRead_lo_lo_lo_4};
  wire [1:0]  tryToRead_lo_hi_lo_lo_4 = {inputSelect1H_9[4], inputSelect1H_8[4]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_4 = {inputSelect1H_11[4], inputSelect1H_10[4]};
  wire [3:0]  tryToRead_lo_hi_lo_4 = {tryToRead_lo_hi_lo_hi_4, tryToRead_lo_hi_lo_lo_4};
  wire [1:0]  tryToRead_lo_hi_hi_lo_4 = {inputSelect1H_13[4], inputSelect1H_12[4]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_4 = {inputSelect1H_15[4], inputSelect1H_14[4]};
  wire [3:0]  tryToRead_lo_hi_hi_4 = {tryToRead_lo_hi_hi_hi_4, tryToRead_lo_hi_hi_lo_4};
  wire [7:0]  tryToRead_lo_hi_4 = {tryToRead_lo_hi_hi_4, tryToRead_lo_hi_lo_4};
  wire [15:0] tryToRead_lo_4 = {tryToRead_lo_hi_4, tryToRead_lo_lo_4};
  wire [1:0]  tryToRead_hi_lo_lo_lo_4 = {inputSelect1H_17[4], inputSelect1H_16[4]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_4 = {inputSelect1H_19[4], inputSelect1H_18[4]};
  wire [3:0]  tryToRead_hi_lo_lo_4 = {tryToRead_hi_lo_lo_hi_4, tryToRead_hi_lo_lo_lo_4};
  wire [1:0]  tryToRead_hi_lo_hi_lo_4 = {inputSelect1H_21[4], inputSelect1H_20[4]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_4 = {inputSelect1H_23[4], inputSelect1H_22[4]};
  wire [3:0]  tryToRead_hi_lo_hi_4 = {tryToRead_hi_lo_hi_hi_4, tryToRead_hi_lo_hi_lo_4};
  wire [7:0]  tryToRead_hi_lo_4 = {tryToRead_hi_lo_hi_4, tryToRead_hi_lo_lo_4};
  wire [1:0]  tryToRead_hi_hi_lo_lo_4 = {inputSelect1H_25[4], inputSelect1H_24[4]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_4 = {inputSelect1H_27[4], inputSelect1H_26[4]};
  wire [3:0]  tryToRead_hi_hi_lo_4 = {tryToRead_hi_hi_lo_hi_4, tryToRead_hi_hi_lo_lo_4};
  wire [1:0]  tryToRead_hi_hi_hi_lo_4 = {inputSelect1H_29[4], inputSelect1H_28[4]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_4 = {inputSelect1H_31[4], inputSelect1H_30[4]};
  wire [3:0]  tryToRead_hi_hi_hi_4 = {tryToRead_hi_hi_hi_hi_4, tryToRead_hi_hi_hi_lo_4};
  wire [7:0]  tryToRead_hi_hi_4 = {tryToRead_hi_hi_hi_4, tryToRead_hi_hi_lo_4};
  wire [15:0] tryToRead_hi_4 = {tryToRead_hi_hi_4, tryToRead_hi_lo_4};
  wire [31:0] tryToRead_4 = {tryToRead_hi_4, tryToRead_lo_4};
  wire        output_4_valid_0 = |tryToRead_4;
  wire [4:0]  output_4_bits_vs_0 = selectReq_4_bits_vs;
  wire        output_4_bits_offset_0 = selectReq_4_bits_offset;
  wire [4:0]  output_4_bits_writeIndex_0 = selectReq_4_bits_requestIndex;
  wire [1:0]  output_4_bits_dataOffset_0 = selectReq_4_bits_dataOffset;
  assign selectReq_4_bits_dataOffset =
    (tryToRead_4[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_4[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_4[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_4[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_4[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_4[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_4[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_4[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_4[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_4[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_4[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_4[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_4[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_4[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_4[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_4[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_4[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_4[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_4[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_4[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_4[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_4[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_4[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_4[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_4[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_4_bits_requestIndex =
    {4'h0, tryToRead_4[1]} | {3'h0, tryToRead_4[2], 1'h0} | (tryToRead_4[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_4[4], 2'h0} | (tryToRead_4[5] ? 5'h5 : 5'h0) | (tryToRead_4[6] ? 5'h6 : 5'h0) | (tryToRead_4[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_4[8], 3'h0} | (tryToRead_4[9] ? 5'h9 : 5'h0) | (tryToRead_4[10] ? 5'hA : 5'h0) | (tryToRead_4[11] ? 5'hB : 5'h0) | (tryToRead_4[12] ? 5'hC : 5'h0) | (tryToRead_4[13] ? 5'hD : 5'h0) | (tryToRead_4[14] ? 5'hE : 5'h0)
    | (tryToRead_4[15] ? 5'hF : 5'h0) | {tryToRead_4[16], 4'h0} | (tryToRead_4[17] ? 5'h11 : 5'h0) | (tryToRead_4[18] ? 5'h12 : 5'h0) | (tryToRead_4[19] ? 5'h13 : 5'h0) | (tryToRead_4[20] ? 5'h14 : 5'h0) | (tryToRead_4[21] ? 5'h15 : 5'h0)
    | (tryToRead_4[22] ? 5'h16 : 5'h0) | (tryToRead_4[23] ? 5'h17 : 5'h0) | (tryToRead_4[24] ? 5'h18 : 5'h0) | (tryToRead_4[25] ? 5'h19 : 5'h0) | (tryToRead_4[26] ? 5'h1A : 5'h0) | (tryToRead_4[27] ? 5'h1B : 5'h0)
    | (tryToRead_4[28] ? 5'h1C : 5'h0) | (tryToRead_4[29] ? 5'h1D : 5'h0) | (tryToRead_4[30] ? 5'h1E : 5'h0) | {5{tryToRead_4[31]}};
  wire [4:0]  selectReq_4_bits_readLane =
    (tryToRead_4[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_4[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_4[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_4[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_4[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_4[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_4[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_4[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_4[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_4[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_4[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_4[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_4[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_4[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_4[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_4[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_4[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_4[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_4[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_4[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_4[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_4[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_4[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_4[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_4[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_4[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_4[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_4[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_4[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_4[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_4[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_4[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_4_bits_offset =
    tryToRead_4[0] & input_0_bits_offset_0 | tryToRead_4[1] & input_1_bits_offset_0 | tryToRead_4[2] & input_2_bits_offset_0 | tryToRead_4[3] & input_3_bits_offset_0 | tryToRead_4[4] & input_4_bits_offset_0 | tryToRead_4[5]
    & input_5_bits_offset_0 | tryToRead_4[6] & input_6_bits_offset_0 | tryToRead_4[7] & input_7_bits_offset_0 | tryToRead_4[8] & input_8_bits_offset_0 | tryToRead_4[9] & input_9_bits_offset_0 | tryToRead_4[10] & input_10_bits_offset_0
    | tryToRead_4[11] & input_11_bits_offset_0 | tryToRead_4[12] & input_12_bits_offset_0 | tryToRead_4[13] & input_13_bits_offset_0 | tryToRead_4[14] & input_14_bits_offset_0 | tryToRead_4[15] & input_15_bits_offset_0 | tryToRead_4[16]
    & input_16_bits_offset_0 | tryToRead_4[17] & input_17_bits_offset_0 | tryToRead_4[18] & input_18_bits_offset_0 | tryToRead_4[19] & input_19_bits_offset_0 | tryToRead_4[20] & input_20_bits_offset_0 | tryToRead_4[21]
    & input_21_bits_offset_0 | tryToRead_4[22] & input_22_bits_offset_0 | tryToRead_4[23] & input_23_bits_offset_0 | tryToRead_4[24] & input_24_bits_offset_0 | tryToRead_4[25] & input_25_bits_offset_0 | tryToRead_4[26]
    & input_26_bits_offset_0 | tryToRead_4[27] & input_27_bits_offset_0 | tryToRead_4[28] & input_28_bits_offset_0 | tryToRead_4[29] & input_29_bits_offset_0 | tryToRead_4[30] & input_30_bits_offset_0 | tryToRead_4[31]
    & input_31_bits_offset_0;
  assign selectReq_4_bits_vs =
    (tryToRead_4[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_4[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_4[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_4[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_4[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_4[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_4[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_4[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_4[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_4[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_4[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_4[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_4[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_4[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_4[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_4[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_4[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_4[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_4[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_4[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_4[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_4[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_4[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_4[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_4[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_4[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_4[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_4[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_4[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_4[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_4[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_4[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_4_valid =
    tryToRead_4[0] & input_0_valid_0 | tryToRead_4[1] & input_1_valid_0 | tryToRead_4[2] & input_2_valid_0 | tryToRead_4[3] & input_3_valid_0 | tryToRead_4[4] & input_4_valid_0 | tryToRead_4[5] & input_5_valid_0 | tryToRead_4[6]
    & input_6_valid_0 | tryToRead_4[7] & input_7_valid_0 | tryToRead_4[8] & input_8_valid_0 | tryToRead_4[9] & input_9_valid_0 | tryToRead_4[10] & input_10_valid_0 | tryToRead_4[11] & input_11_valid_0 | tryToRead_4[12] & input_12_valid_0
    | tryToRead_4[13] & input_13_valid_0 | tryToRead_4[14] & input_14_valid_0 | tryToRead_4[15] & input_15_valid_0 | tryToRead_4[16] & input_16_valid_0 | tryToRead_4[17] & input_17_valid_0 | tryToRead_4[18] & input_18_valid_0
    | tryToRead_4[19] & input_19_valid_0 | tryToRead_4[20] & input_20_valid_0 | tryToRead_4[21] & input_21_valid_0 | tryToRead_4[22] & input_22_valid_0 | tryToRead_4[23] & input_23_valid_0 | tryToRead_4[24] & input_24_valid_0
    | tryToRead_4[25] & input_25_valid_0 | tryToRead_4[26] & input_26_valid_0 | tryToRead_4[27] & input_27_valid_0 | tryToRead_4[28] & input_28_valid_0 | tryToRead_4[29] & input_29_valid_0 | tryToRead_4[30] & input_30_valid_0
    | tryToRead_4[31] & input_31_valid_0;
  wire        selectReq_4_ready =
    tryToRead_4[0] & input_0_ready_0 | tryToRead_4[1] & input_1_ready_0 | tryToRead_4[2] & input_2_ready_0 | tryToRead_4[3] & input_3_ready_0 | tryToRead_4[4] & input_4_ready_0 | tryToRead_4[5] & input_5_ready_0 | tryToRead_4[6]
    & input_6_ready_0 | tryToRead_4[7] & input_7_ready_0 | tryToRead_4[8] & input_8_ready_0 | tryToRead_4[9] & input_9_ready_0 | tryToRead_4[10] & input_10_ready_0 | tryToRead_4[11] & input_11_ready_0 | tryToRead_4[12] & input_12_ready_0
    | tryToRead_4[13] & input_13_ready_0 | tryToRead_4[14] & input_14_ready_0 | tryToRead_4[15] & input_15_ready_0 | tryToRead_4[16] & input_16_ready_0 | tryToRead_4[17] & input_17_ready_0 | tryToRead_4[18] & input_18_ready_0
    | tryToRead_4[19] & input_19_ready_0 | tryToRead_4[20] & input_20_ready_0 | tryToRead_4[21] & input_21_ready_0 | tryToRead_4[22] & input_22_ready_0 | tryToRead_4[23] & input_23_ready_0 | tryToRead_4[24] & input_24_ready_0
    | tryToRead_4[25] & input_25_ready_0 | tryToRead_4[26] & input_26_ready_0 | tryToRead_4[27] & input_27_ready_0 | tryToRead_4[28] & input_28_ready_0 | tryToRead_4[29] & input_29_ready_0 | tryToRead_4[30] & input_30_ready_0
    | tryToRead_4[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_5 = {inputSelect1H_1[5], inputSelect1H_0[5]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_5 = {inputSelect1H_3[5], inputSelect1H_2[5]};
  wire [3:0]  tryToRead_lo_lo_lo_5 = {tryToRead_lo_lo_lo_hi_5, tryToRead_lo_lo_lo_lo_5};
  wire [1:0]  tryToRead_lo_lo_hi_lo_5 = {inputSelect1H_5[5], inputSelect1H_4[5]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_5 = {inputSelect1H_7[5], inputSelect1H_6[5]};
  wire [3:0]  tryToRead_lo_lo_hi_5 = {tryToRead_lo_lo_hi_hi_5, tryToRead_lo_lo_hi_lo_5};
  wire [7:0]  tryToRead_lo_lo_5 = {tryToRead_lo_lo_hi_5, tryToRead_lo_lo_lo_5};
  wire [1:0]  tryToRead_lo_hi_lo_lo_5 = {inputSelect1H_9[5], inputSelect1H_8[5]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_5 = {inputSelect1H_11[5], inputSelect1H_10[5]};
  wire [3:0]  tryToRead_lo_hi_lo_5 = {tryToRead_lo_hi_lo_hi_5, tryToRead_lo_hi_lo_lo_5};
  wire [1:0]  tryToRead_lo_hi_hi_lo_5 = {inputSelect1H_13[5], inputSelect1H_12[5]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_5 = {inputSelect1H_15[5], inputSelect1H_14[5]};
  wire [3:0]  tryToRead_lo_hi_hi_5 = {tryToRead_lo_hi_hi_hi_5, tryToRead_lo_hi_hi_lo_5};
  wire [7:0]  tryToRead_lo_hi_5 = {tryToRead_lo_hi_hi_5, tryToRead_lo_hi_lo_5};
  wire [15:0] tryToRead_lo_5 = {tryToRead_lo_hi_5, tryToRead_lo_lo_5};
  wire [1:0]  tryToRead_hi_lo_lo_lo_5 = {inputSelect1H_17[5], inputSelect1H_16[5]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_5 = {inputSelect1H_19[5], inputSelect1H_18[5]};
  wire [3:0]  tryToRead_hi_lo_lo_5 = {tryToRead_hi_lo_lo_hi_5, tryToRead_hi_lo_lo_lo_5};
  wire [1:0]  tryToRead_hi_lo_hi_lo_5 = {inputSelect1H_21[5], inputSelect1H_20[5]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_5 = {inputSelect1H_23[5], inputSelect1H_22[5]};
  wire [3:0]  tryToRead_hi_lo_hi_5 = {tryToRead_hi_lo_hi_hi_5, tryToRead_hi_lo_hi_lo_5};
  wire [7:0]  tryToRead_hi_lo_5 = {tryToRead_hi_lo_hi_5, tryToRead_hi_lo_lo_5};
  wire [1:0]  tryToRead_hi_hi_lo_lo_5 = {inputSelect1H_25[5], inputSelect1H_24[5]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_5 = {inputSelect1H_27[5], inputSelect1H_26[5]};
  wire [3:0]  tryToRead_hi_hi_lo_5 = {tryToRead_hi_hi_lo_hi_5, tryToRead_hi_hi_lo_lo_5};
  wire [1:0]  tryToRead_hi_hi_hi_lo_5 = {inputSelect1H_29[5], inputSelect1H_28[5]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_5 = {inputSelect1H_31[5], inputSelect1H_30[5]};
  wire [3:0]  tryToRead_hi_hi_hi_5 = {tryToRead_hi_hi_hi_hi_5, tryToRead_hi_hi_hi_lo_5};
  wire [7:0]  tryToRead_hi_hi_5 = {tryToRead_hi_hi_hi_5, tryToRead_hi_hi_lo_5};
  wire [15:0] tryToRead_hi_5 = {tryToRead_hi_hi_5, tryToRead_hi_lo_5};
  wire [31:0] tryToRead_5 = {tryToRead_hi_5, tryToRead_lo_5};
  wire        output_5_valid_0 = |tryToRead_5;
  wire [4:0]  output_5_bits_vs_0 = selectReq_5_bits_vs;
  wire        output_5_bits_offset_0 = selectReq_5_bits_offset;
  wire [4:0]  output_5_bits_writeIndex_0 = selectReq_5_bits_requestIndex;
  wire [1:0]  output_5_bits_dataOffset_0 = selectReq_5_bits_dataOffset;
  assign selectReq_5_bits_dataOffset =
    (tryToRead_5[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_5[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_5[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_5[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_5[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_5[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_5[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_5[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_5[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_5[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_5[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_5[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_5[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_5[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_5[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_5[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_5[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_5[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_5[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_5[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_5[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_5[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_5[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_5[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_5[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_5_bits_requestIndex =
    {4'h0, tryToRead_5[1]} | {3'h0, tryToRead_5[2], 1'h0} | (tryToRead_5[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_5[4], 2'h0} | (tryToRead_5[5] ? 5'h5 : 5'h0) | (tryToRead_5[6] ? 5'h6 : 5'h0) | (tryToRead_5[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_5[8], 3'h0} | (tryToRead_5[9] ? 5'h9 : 5'h0) | (tryToRead_5[10] ? 5'hA : 5'h0) | (tryToRead_5[11] ? 5'hB : 5'h0) | (tryToRead_5[12] ? 5'hC : 5'h0) | (tryToRead_5[13] ? 5'hD : 5'h0) | (tryToRead_5[14] ? 5'hE : 5'h0)
    | (tryToRead_5[15] ? 5'hF : 5'h0) | {tryToRead_5[16], 4'h0} | (tryToRead_5[17] ? 5'h11 : 5'h0) | (tryToRead_5[18] ? 5'h12 : 5'h0) | (tryToRead_5[19] ? 5'h13 : 5'h0) | (tryToRead_5[20] ? 5'h14 : 5'h0) | (tryToRead_5[21] ? 5'h15 : 5'h0)
    | (tryToRead_5[22] ? 5'h16 : 5'h0) | (tryToRead_5[23] ? 5'h17 : 5'h0) | (tryToRead_5[24] ? 5'h18 : 5'h0) | (tryToRead_5[25] ? 5'h19 : 5'h0) | (tryToRead_5[26] ? 5'h1A : 5'h0) | (tryToRead_5[27] ? 5'h1B : 5'h0)
    | (tryToRead_5[28] ? 5'h1C : 5'h0) | (tryToRead_5[29] ? 5'h1D : 5'h0) | (tryToRead_5[30] ? 5'h1E : 5'h0) | {5{tryToRead_5[31]}};
  wire [4:0]  selectReq_5_bits_readLane =
    (tryToRead_5[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_5[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_5[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_5[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_5[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_5[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_5[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_5[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_5[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_5[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_5[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_5[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_5[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_5[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_5[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_5[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_5[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_5[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_5[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_5[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_5[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_5[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_5[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_5[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_5[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_5[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_5[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_5[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_5[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_5[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_5[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_5[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_5_bits_offset =
    tryToRead_5[0] & input_0_bits_offset_0 | tryToRead_5[1] & input_1_bits_offset_0 | tryToRead_5[2] & input_2_bits_offset_0 | tryToRead_5[3] & input_3_bits_offset_0 | tryToRead_5[4] & input_4_bits_offset_0 | tryToRead_5[5]
    & input_5_bits_offset_0 | tryToRead_5[6] & input_6_bits_offset_0 | tryToRead_5[7] & input_7_bits_offset_0 | tryToRead_5[8] & input_8_bits_offset_0 | tryToRead_5[9] & input_9_bits_offset_0 | tryToRead_5[10] & input_10_bits_offset_0
    | tryToRead_5[11] & input_11_bits_offset_0 | tryToRead_5[12] & input_12_bits_offset_0 | tryToRead_5[13] & input_13_bits_offset_0 | tryToRead_5[14] & input_14_bits_offset_0 | tryToRead_5[15] & input_15_bits_offset_0 | tryToRead_5[16]
    & input_16_bits_offset_0 | tryToRead_5[17] & input_17_bits_offset_0 | tryToRead_5[18] & input_18_bits_offset_0 | tryToRead_5[19] & input_19_bits_offset_0 | tryToRead_5[20] & input_20_bits_offset_0 | tryToRead_5[21]
    & input_21_bits_offset_0 | tryToRead_5[22] & input_22_bits_offset_0 | tryToRead_5[23] & input_23_bits_offset_0 | tryToRead_5[24] & input_24_bits_offset_0 | tryToRead_5[25] & input_25_bits_offset_0 | tryToRead_5[26]
    & input_26_bits_offset_0 | tryToRead_5[27] & input_27_bits_offset_0 | tryToRead_5[28] & input_28_bits_offset_0 | tryToRead_5[29] & input_29_bits_offset_0 | tryToRead_5[30] & input_30_bits_offset_0 | tryToRead_5[31]
    & input_31_bits_offset_0;
  assign selectReq_5_bits_vs =
    (tryToRead_5[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_5[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_5[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_5[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_5[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_5[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_5[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_5[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_5[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_5[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_5[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_5[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_5[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_5[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_5[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_5[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_5[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_5[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_5[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_5[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_5[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_5[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_5[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_5[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_5[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_5[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_5[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_5[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_5[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_5[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_5[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_5[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_5_valid =
    tryToRead_5[0] & input_0_valid_0 | tryToRead_5[1] & input_1_valid_0 | tryToRead_5[2] & input_2_valid_0 | tryToRead_5[3] & input_3_valid_0 | tryToRead_5[4] & input_4_valid_0 | tryToRead_5[5] & input_5_valid_0 | tryToRead_5[6]
    & input_6_valid_0 | tryToRead_5[7] & input_7_valid_0 | tryToRead_5[8] & input_8_valid_0 | tryToRead_5[9] & input_9_valid_0 | tryToRead_5[10] & input_10_valid_0 | tryToRead_5[11] & input_11_valid_0 | tryToRead_5[12] & input_12_valid_0
    | tryToRead_5[13] & input_13_valid_0 | tryToRead_5[14] & input_14_valid_0 | tryToRead_5[15] & input_15_valid_0 | tryToRead_5[16] & input_16_valid_0 | tryToRead_5[17] & input_17_valid_0 | tryToRead_5[18] & input_18_valid_0
    | tryToRead_5[19] & input_19_valid_0 | tryToRead_5[20] & input_20_valid_0 | tryToRead_5[21] & input_21_valid_0 | tryToRead_5[22] & input_22_valid_0 | tryToRead_5[23] & input_23_valid_0 | tryToRead_5[24] & input_24_valid_0
    | tryToRead_5[25] & input_25_valid_0 | tryToRead_5[26] & input_26_valid_0 | tryToRead_5[27] & input_27_valid_0 | tryToRead_5[28] & input_28_valid_0 | tryToRead_5[29] & input_29_valid_0 | tryToRead_5[30] & input_30_valid_0
    | tryToRead_5[31] & input_31_valid_0;
  wire        selectReq_5_ready =
    tryToRead_5[0] & input_0_ready_0 | tryToRead_5[1] & input_1_ready_0 | tryToRead_5[2] & input_2_ready_0 | tryToRead_5[3] & input_3_ready_0 | tryToRead_5[4] & input_4_ready_0 | tryToRead_5[5] & input_5_ready_0 | tryToRead_5[6]
    & input_6_ready_0 | tryToRead_5[7] & input_7_ready_0 | tryToRead_5[8] & input_8_ready_0 | tryToRead_5[9] & input_9_ready_0 | tryToRead_5[10] & input_10_ready_0 | tryToRead_5[11] & input_11_ready_0 | tryToRead_5[12] & input_12_ready_0
    | tryToRead_5[13] & input_13_ready_0 | tryToRead_5[14] & input_14_ready_0 | tryToRead_5[15] & input_15_ready_0 | tryToRead_5[16] & input_16_ready_0 | tryToRead_5[17] & input_17_ready_0 | tryToRead_5[18] & input_18_ready_0
    | tryToRead_5[19] & input_19_ready_0 | tryToRead_5[20] & input_20_ready_0 | tryToRead_5[21] & input_21_ready_0 | tryToRead_5[22] & input_22_ready_0 | tryToRead_5[23] & input_23_ready_0 | tryToRead_5[24] & input_24_ready_0
    | tryToRead_5[25] & input_25_ready_0 | tryToRead_5[26] & input_26_ready_0 | tryToRead_5[27] & input_27_ready_0 | tryToRead_5[28] & input_28_ready_0 | tryToRead_5[29] & input_29_ready_0 | tryToRead_5[30] & input_30_ready_0
    | tryToRead_5[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_6 = {inputSelect1H_1[6], inputSelect1H_0[6]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_6 = {inputSelect1H_3[6], inputSelect1H_2[6]};
  wire [3:0]  tryToRead_lo_lo_lo_6 = {tryToRead_lo_lo_lo_hi_6, tryToRead_lo_lo_lo_lo_6};
  wire [1:0]  tryToRead_lo_lo_hi_lo_6 = {inputSelect1H_5[6], inputSelect1H_4[6]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_6 = {inputSelect1H_7[6], inputSelect1H_6[6]};
  wire [3:0]  tryToRead_lo_lo_hi_6 = {tryToRead_lo_lo_hi_hi_6, tryToRead_lo_lo_hi_lo_6};
  wire [7:0]  tryToRead_lo_lo_6 = {tryToRead_lo_lo_hi_6, tryToRead_lo_lo_lo_6};
  wire [1:0]  tryToRead_lo_hi_lo_lo_6 = {inputSelect1H_9[6], inputSelect1H_8[6]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_6 = {inputSelect1H_11[6], inputSelect1H_10[6]};
  wire [3:0]  tryToRead_lo_hi_lo_6 = {tryToRead_lo_hi_lo_hi_6, tryToRead_lo_hi_lo_lo_6};
  wire [1:0]  tryToRead_lo_hi_hi_lo_6 = {inputSelect1H_13[6], inputSelect1H_12[6]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_6 = {inputSelect1H_15[6], inputSelect1H_14[6]};
  wire [3:0]  tryToRead_lo_hi_hi_6 = {tryToRead_lo_hi_hi_hi_6, tryToRead_lo_hi_hi_lo_6};
  wire [7:0]  tryToRead_lo_hi_6 = {tryToRead_lo_hi_hi_6, tryToRead_lo_hi_lo_6};
  wire [15:0] tryToRead_lo_6 = {tryToRead_lo_hi_6, tryToRead_lo_lo_6};
  wire [1:0]  tryToRead_hi_lo_lo_lo_6 = {inputSelect1H_17[6], inputSelect1H_16[6]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_6 = {inputSelect1H_19[6], inputSelect1H_18[6]};
  wire [3:0]  tryToRead_hi_lo_lo_6 = {tryToRead_hi_lo_lo_hi_6, tryToRead_hi_lo_lo_lo_6};
  wire [1:0]  tryToRead_hi_lo_hi_lo_6 = {inputSelect1H_21[6], inputSelect1H_20[6]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_6 = {inputSelect1H_23[6], inputSelect1H_22[6]};
  wire [3:0]  tryToRead_hi_lo_hi_6 = {tryToRead_hi_lo_hi_hi_6, tryToRead_hi_lo_hi_lo_6};
  wire [7:0]  tryToRead_hi_lo_6 = {tryToRead_hi_lo_hi_6, tryToRead_hi_lo_lo_6};
  wire [1:0]  tryToRead_hi_hi_lo_lo_6 = {inputSelect1H_25[6], inputSelect1H_24[6]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_6 = {inputSelect1H_27[6], inputSelect1H_26[6]};
  wire [3:0]  tryToRead_hi_hi_lo_6 = {tryToRead_hi_hi_lo_hi_6, tryToRead_hi_hi_lo_lo_6};
  wire [1:0]  tryToRead_hi_hi_hi_lo_6 = {inputSelect1H_29[6], inputSelect1H_28[6]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_6 = {inputSelect1H_31[6], inputSelect1H_30[6]};
  wire [3:0]  tryToRead_hi_hi_hi_6 = {tryToRead_hi_hi_hi_hi_6, tryToRead_hi_hi_hi_lo_6};
  wire [7:0]  tryToRead_hi_hi_6 = {tryToRead_hi_hi_hi_6, tryToRead_hi_hi_lo_6};
  wire [15:0] tryToRead_hi_6 = {tryToRead_hi_hi_6, tryToRead_hi_lo_6};
  wire [31:0] tryToRead_6 = {tryToRead_hi_6, tryToRead_lo_6};
  wire        output_6_valid_0 = |tryToRead_6;
  wire [4:0]  output_6_bits_vs_0 = selectReq_6_bits_vs;
  wire        output_6_bits_offset_0 = selectReq_6_bits_offset;
  wire [4:0]  output_6_bits_writeIndex_0 = selectReq_6_bits_requestIndex;
  wire [1:0]  output_6_bits_dataOffset_0 = selectReq_6_bits_dataOffset;
  assign selectReq_6_bits_dataOffset =
    (tryToRead_6[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_6[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_6[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_6[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_6[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_6[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_6[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_6[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_6[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_6[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_6[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_6[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_6[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_6[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_6[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_6[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_6[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_6[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_6[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_6[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_6[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_6[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_6[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_6[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_6[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_6_bits_requestIndex =
    {4'h0, tryToRead_6[1]} | {3'h0, tryToRead_6[2], 1'h0} | (tryToRead_6[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_6[4], 2'h0} | (tryToRead_6[5] ? 5'h5 : 5'h0) | (tryToRead_6[6] ? 5'h6 : 5'h0) | (tryToRead_6[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_6[8], 3'h0} | (tryToRead_6[9] ? 5'h9 : 5'h0) | (tryToRead_6[10] ? 5'hA : 5'h0) | (tryToRead_6[11] ? 5'hB : 5'h0) | (tryToRead_6[12] ? 5'hC : 5'h0) | (tryToRead_6[13] ? 5'hD : 5'h0) | (tryToRead_6[14] ? 5'hE : 5'h0)
    | (tryToRead_6[15] ? 5'hF : 5'h0) | {tryToRead_6[16], 4'h0} | (tryToRead_6[17] ? 5'h11 : 5'h0) | (tryToRead_6[18] ? 5'h12 : 5'h0) | (tryToRead_6[19] ? 5'h13 : 5'h0) | (tryToRead_6[20] ? 5'h14 : 5'h0) | (tryToRead_6[21] ? 5'h15 : 5'h0)
    | (tryToRead_6[22] ? 5'h16 : 5'h0) | (tryToRead_6[23] ? 5'h17 : 5'h0) | (tryToRead_6[24] ? 5'h18 : 5'h0) | (tryToRead_6[25] ? 5'h19 : 5'h0) | (tryToRead_6[26] ? 5'h1A : 5'h0) | (tryToRead_6[27] ? 5'h1B : 5'h0)
    | (tryToRead_6[28] ? 5'h1C : 5'h0) | (tryToRead_6[29] ? 5'h1D : 5'h0) | (tryToRead_6[30] ? 5'h1E : 5'h0) | {5{tryToRead_6[31]}};
  wire [4:0]  selectReq_6_bits_readLane =
    (tryToRead_6[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_6[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_6[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_6[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_6[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_6[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_6[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_6[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_6[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_6[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_6[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_6[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_6[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_6[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_6[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_6[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_6[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_6[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_6[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_6[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_6[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_6[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_6[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_6[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_6[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_6[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_6[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_6[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_6[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_6[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_6[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_6[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_6_bits_offset =
    tryToRead_6[0] & input_0_bits_offset_0 | tryToRead_6[1] & input_1_bits_offset_0 | tryToRead_6[2] & input_2_bits_offset_0 | tryToRead_6[3] & input_3_bits_offset_0 | tryToRead_6[4] & input_4_bits_offset_0 | tryToRead_6[5]
    & input_5_bits_offset_0 | tryToRead_6[6] & input_6_bits_offset_0 | tryToRead_6[7] & input_7_bits_offset_0 | tryToRead_6[8] & input_8_bits_offset_0 | tryToRead_6[9] & input_9_bits_offset_0 | tryToRead_6[10] & input_10_bits_offset_0
    | tryToRead_6[11] & input_11_bits_offset_0 | tryToRead_6[12] & input_12_bits_offset_0 | tryToRead_6[13] & input_13_bits_offset_0 | tryToRead_6[14] & input_14_bits_offset_0 | tryToRead_6[15] & input_15_bits_offset_0 | tryToRead_6[16]
    & input_16_bits_offset_0 | tryToRead_6[17] & input_17_bits_offset_0 | tryToRead_6[18] & input_18_bits_offset_0 | tryToRead_6[19] & input_19_bits_offset_0 | tryToRead_6[20] & input_20_bits_offset_0 | tryToRead_6[21]
    & input_21_bits_offset_0 | tryToRead_6[22] & input_22_bits_offset_0 | tryToRead_6[23] & input_23_bits_offset_0 | tryToRead_6[24] & input_24_bits_offset_0 | tryToRead_6[25] & input_25_bits_offset_0 | tryToRead_6[26]
    & input_26_bits_offset_0 | tryToRead_6[27] & input_27_bits_offset_0 | tryToRead_6[28] & input_28_bits_offset_0 | tryToRead_6[29] & input_29_bits_offset_0 | tryToRead_6[30] & input_30_bits_offset_0 | tryToRead_6[31]
    & input_31_bits_offset_0;
  assign selectReq_6_bits_vs =
    (tryToRead_6[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_6[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_6[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_6[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_6[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_6[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_6[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_6[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_6[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_6[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_6[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_6[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_6[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_6[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_6[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_6[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_6[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_6[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_6[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_6[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_6[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_6[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_6[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_6[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_6[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_6[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_6[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_6[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_6[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_6[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_6[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_6[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_6_valid =
    tryToRead_6[0] & input_0_valid_0 | tryToRead_6[1] & input_1_valid_0 | tryToRead_6[2] & input_2_valid_0 | tryToRead_6[3] & input_3_valid_0 | tryToRead_6[4] & input_4_valid_0 | tryToRead_6[5] & input_5_valid_0 | tryToRead_6[6]
    & input_6_valid_0 | tryToRead_6[7] & input_7_valid_0 | tryToRead_6[8] & input_8_valid_0 | tryToRead_6[9] & input_9_valid_0 | tryToRead_6[10] & input_10_valid_0 | tryToRead_6[11] & input_11_valid_0 | tryToRead_6[12] & input_12_valid_0
    | tryToRead_6[13] & input_13_valid_0 | tryToRead_6[14] & input_14_valid_0 | tryToRead_6[15] & input_15_valid_0 | tryToRead_6[16] & input_16_valid_0 | tryToRead_6[17] & input_17_valid_0 | tryToRead_6[18] & input_18_valid_0
    | tryToRead_6[19] & input_19_valid_0 | tryToRead_6[20] & input_20_valid_0 | tryToRead_6[21] & input_21_valid_0 | tryToRead_6[22] & input_22_valid_0 | tryToRead_6[23] & input_23_valid_0 | tryToRead_6[24] & input_24_valid_0
    | tryToRead_6[25] & input_25_valid_0 | tryToRead_6[26] & input_26_valid_0 | tryToRead_6[27] & input_27_valid_0 | tryToRead_6[28] & input_28_valid_0 | tryToRead_6[29] & input_29_valid_0 | tryToRead_6[30] & input_30_valid_0
    | tryToRead_6[31] & input_31_valid_0;
  wire        selectReq_6_ready =
    tryToRead_6[0] & input_0_ready_0 | tryToRead_6[1] & input_1_ready_0 | tryToRead_6[2] & input_2_ready_0 | tryToRead_6[3] & input_3_ready_0 | tryToRead_6[4] & input_4_ready_0 | tryToRead_6[5] & input_5_ready_0 | tryToRead_6[6]
    & input_6_ready_0 | tryToRead_6[7] & input_7_ready_0 | tryToRead_6[8] & input_8_ready_0 | tryToRead_6[9] & input_9_ready_0 | tryToRead_6[10] & input_10_ready_0 | tryToRead_6[11] & input_11_ready_0 | tryToRead_6[12] & input_12_ready_0
    | tryToRead_6[13] & input_13_ready_0 | tryToRead_6[14] & input_14_ready_0 | tryToRead_6[15] & input_15_ready_0 | tryToRead_6[16] & input_16_ready_0 | tryToRead_6[17] & input_17_ready_0 | tryToRead_6[18] & input_18_ready_0
    | tryToRead_6[19] & input_19_ready_0 | tryToRead_6[20] & input_20_ready_0 | tryToRead_6[21] & input_21_ready_0 | tryToRead_6[22] & input_22_ready_0 | tryToRead_6[23] & input_23_ready_0 | tryToRead_6[24] & input_24_ready_0
    | tryToRead_6[25] & input_25_ready_0 | tryToRead_6[26] & input_26_ready_0 | tryToRead_6[27] & input_27_ready_0 | tryToRead_6[28] & input_28_ready_0 | tryToRead_6[29] & input_29_ready_0 | tryToRead_6[30] & input_30_ready_0
    | tryToRead_6[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_7 = {inputSelect1H_1[7], inputSelect1H_0[7]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_7 = {inputSelect1H_3[7], inputSelect1H_2[7]};
  wire [3:0]  tryToRead_lo_lo_lo_7 = {tryToRead_lo_lo_lo_hi_7, tryToRead_lo_lo_lo_lo_7};
  wire [1:0]  tryToRead_lo_lo_hi_lo_7 = {inputSelect1H_5[7], inputSelect1H_4[7]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_7 = {inputSelect1H_7[7], inputSelect1H_6[7]};
  wire [3:0]  tryToRead_lo_lo_hi_7 = {tryToRead_lo_lo_hi_hi_7, tryToRead_lo_lo_hi_lo_7};
  wire [7:0]  tryToRead_lo_lo_7 = {tryToRead_lo_lo_hi_7, tryToRead_lo_lo_lo_7};
  wire [1:0]  tryToRead_lo_hi_lo_lo_7 = {inputSelect1H_9[7], inputSelect1H_8[7]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_7 = {inputSelect1H_11[7], inputSelect1H_10[7]};
  wire [3:0]  tryToRead_lo_hi_lo_7 = {tryToRead_lo_hi_lo_hi_7, tryToRead_lo_hi_lo_lo_7};
  wire [1:0]  tryToRead_lo_hi_hi_lo_7 = {inputSelect1H_13[7], inputSelect1H_12[7]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_7 = {inputSelect1H_15[7], inputSelect1H_14[7]};
  wire [3:0]  tryToRead_lo_hi_hi_7 = {tryToRead_lo_hi_hi_hi_7, tryToRead_lo_hi_hi_lo_7};
  wire [7:0]  tryToRead_lo_hi_7 = {tryToRead_lo_hi_hi_7, tryToRead_lo_hi_lo_7};
  wire [15:0] tryToRead_lo_7 = {tryToRead_lo_hi_7, tryToRead_lo_lo_7};
  wire [1:0]  tryToRead_hi_lo_lo_lo_7 = {inputSelect1H_17[7], inputSelect1H_16[7]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_7 = {inputSelect1H_19[7], inputSelect1H_18[7]};
  wire [3:0]  tryToRead_hi_lo_lo_7 = {tryToRead_hi_lo_lo_hi_7, tryToRead_hi_lo_lo_lo_7};
  wire [1:0]  tryToRead_hi_lo_hi_lo_7 = {inputSelect1H_21[7], inputSelect1H_20[7]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_7 = {inputSelect1H_23[7], inputSelect1H_22[7]};
  wire [3:0]  tryToRead_hi_lo_hi_7 = {tryToRead_hi_lo_hi_hi_7, tryToRead_hi_lo_hi_lo_7};
  wire [7:0]  tryToRead_hi_lo_7 = {tryToRead_hi_lo_hi_7, tryToRead_hi_lo_lo_7};
  wire [1:0]  tryToRead_hi_hi_lo_lo_7 = {inputSelect1H_25[7], inputSelect1H_24[7]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_7 = {inputSelect1H_27[7], inputSelect1H_26[7]};
  wire [3:0]  tryToRead_hi_hi_lo_7 = {tryToRead_hi_hi_lo_hi_7, tryToRead_hi_hi_lo_lo_7};
  wire [1:0]  tryToRead_hi_hi_hi_lo_7 = {inputSelect1H_29[7], inputSelect1H_28[7]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_7 = {inputSelect1H_31[7], inputSelect1H_30[7]};
  wire [3:0]  tryToRead_hi_hi_hi_7 = {tryToRead_hi_hi_hi_hi_7, tryToRead_hi_hi_hi_lo_7};
  wire [7:0]  tryToRead_hi_hi_7 = {tryToRead_hi_hi_hi_7, tryToRead_hi_hi_lo_7};
  wire [15:0] tryToRead_hi_7 = {tryToRead_hi_hi_7, tryToRead_hi_lo_7};
  wire [31:0] tryToRead_7 = {tryToRead_hi_7, tryToRead_lo_7};
  wire        output_7_valid_0 = |tryToRead_7;
  wire [4:0]  output_7_bits_vs_0 = selectReq_7_bits_vs;
  wire        output_7_bits_offset_0 = selectReq_7_bits_offset;
  wire [4:0]  output_7_bits_writeIndex_0 = selectReq_7_bits_requestIndex;
  wire [1:0]  output_7_bits_dataOffset_0 = selectReq_7_bits_dataOffset;
  assign selectReq_7_bits_dataOffset =
    (tryToRead_7[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_7[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_7[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_7[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_7[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_7[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_7[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_7[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_7[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_7[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_7[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_7[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_7[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_7[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_7[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_7[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_7[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_7[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_7[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_7[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_7[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_7[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_7[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_7[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_7[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_7_bits_requestIndex =
    {4'h0, tryToRead_7[1]} | {3'h0, tryToRead_7[2], 1'h0} | (tryToRead_7[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_7[4], 2'h0} | (tryToRead_7[5] ? 5'h5 : 5'h0) | (tryToRead_7[6] ? 5'h6 : 5'h0) | (tryToRead_7[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_7[8], 3'h0} | (tryToRead_7[9] ? 5'h9 : 5'h0) | (tryToRead_7[10] ? 5'hA : 5'h0) | (tryToRead_7[11] ? 5'hB : 5'h0) | (tryToRead_7[12] ? 5'hC : 5'h0) | (tryToRead_7[13] ? 5'hD : 5'h0) | (tryToRead_7[14] ? 5'hE : 5'h0)
    | (tryToRead_7[15] ? 5'hF : 5'h0) | {tryToRead_7[16], 4'h0} | (tryToRead_7[17] ? 5'h11 : 5'h0) | (tryToRead_7[18] ? 5'h12 : 5'h0) | (tryToRead_7[19] ? 5'h13 : 5'h0) | (tryToRead_7[20] ? 5'h14 : 5'h0) | (tryToRead_7[21] ? 5'h15 : 5'h0)
    | (tryToRead_7[22] ? 5'h16 : 5'h0) | (tryToRead_7[23] ? 5'h17 : 5'h0) | (tryToRead_7[24] ? 5'h18 : 5'h0) | (tryToRead_7[25] ? 5'h19 : 5'h0) | (tryToRead_7[26] ? 5'h1A : 5'h0) | (tryToRead_7[27] ? 5'h1B : 5'h0)
    | (tryToRead_7[28] ? 5'h1C : 5'h0) | (tryToRead_7[29] ? 5'h1D : 5'h0) | (tryToRead_7[30] ? 5'h1E : 5'h0) | {5{tryToRead_7[31]}};
  wire [4:0]  selectReq_7_bits_readLane =
    (tryToRead_7[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_7[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_7[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_7[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_7[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_7[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_7[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_7[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_7[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_7[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_7[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_7[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_7[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_7[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_7[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_7[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_7[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_7[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_7[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_7[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_7[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_7[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_7[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_7[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_7[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_7[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_7[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_7[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_7[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_7[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_7[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_7[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_7_bits_offset =
    tryToRead_7[0] & input_0_bits_offset_0 | tryToRead_7[1] & input_1_bits_offset_0 | tryToRead_7[2] & input_2_bits_offset_0 | tryToRead_7[3] & input_3_bits_offset_0 | tryToRead_7[4] & input_4_bits_offset_0 | tryToRead_7[5]
    & input_5_bits_offset_0 | tryToRead_7[6] & input_6_bits_offset_0 | tryToRead_7[7] & input_7_bits_offset_0 | tryToRead_7[8] & input_8_bits_offset_0 | tryToRead_7[9] & input_9_bits_offset_0 | tryToRead_7[10] & input_10_bits_offset_0
    | tryToRead_7[11] & input_11_bits_offset_0 | tryToRead_7[12] & input_12_bits_offset_0 | tryToRead_7[13] & input_13_bits_offset_0 | tryToRead_7[14] & input_14_bits_offset_0 | tryToRead_7[15] & input_15_bits_offset_0 | tryToRead_7[16]
    & input_16_bits_offset_0 | tryToRead_7[17] & input_17_bits_offset_0 | tryToRead_7[18] & input_18_bits_offset_0 | tryToRead_7[19] & input_19_bits_offset_0 | tryToRead_7[20] & input_20_bits_offset_0 | tryToRead_7[21]
    & input_21_bits_offset_0 | tryToRead_7[22] & input_22_bits_offset_0 | tryToRead_7[23] & input_23_bits_offset_0 | tryToRead_7[24] & input_24_bits_offset_0 | tryToRead_7[25] & input_25_bits_offset_0 | tryToRead_7[26]
    & input_26_bits_offset_0 | tryToRead_7[27] & input_27_bits_offset_0 | tryToRead_7[28] & input_28_bits_offset_0 | tryToRead_7[29] & input_29_bits_offset_0 | tryToRead_7[30] & input_30_bits_offset_0 | tryToRead_7[31]
    & input_31_bits_offset_0;
  assign selectReq_7_bits_vs =
    (tryToRead_7[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_7[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_7[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_7[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_7[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_7[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_7[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_7[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_7[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_7[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_7[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_7[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_7[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_7[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_7[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_7[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_7[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_7[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_7[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_7[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_7[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_7[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_7[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_7[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_7[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_7[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_7[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_7[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_7[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_7[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_7[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_7[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_7_valid =
    tryToRead_7[0] & input_0_valid_0 | tryToRead_7[1] & input_1_valid_0 | tryToRead_7[2] & input_2_valid_0 | tryToRead_7[3] & input_3_valid_0 | tryToRead_7[4] & input_4_valid_0 | tryToRead_7[5] & input_5_valid_0 | tryToRead_7[6]
    & input_6_valid_0 | tryToRead_7[7] & input_7_valid_0 | tryToRead_7[8] & input_8_valid_0 | tryToRead_7[9] & input_9_valid_0 | tryToRead_7[10] & input_10_valid_0 | tryToRead_7[11] & input_11_valid_0 | tryToRead_7[12] & input_12_valid_0
    | tryToRead_7[13] & input_13_valid_0 | tryToRead_7[14] & input_14_valid_0 | tryToRead_7[15] & input_15_valid_0 | tryToRead_7[16] & input_16_valid_0 | tryToRead_7[17] & input_17_valid_0 | tryToRead_7[18] & input_18_valid_0
    | tryToRead_7[19] & input_19_valid_0 | tryToRead_7[20] & input_20_valid_0 | tryToRead_7[21] & input_21_valid_0 | tryToRead_7[22] & input_22_valid_0 | tryToRead_7[23] & input_23_valid_0 | tryToRead_7[24] & input_24_valid_0
    | tryToRead_7[25] & input_25_valid_0 | tryToRead_7[26] & input_26_valid_0 | tryToRead_7[27] & input_27_valid_0 | tryToRead_7[28] & input_28_valid_0 | tryToRead_7[29] & input_29_valid_0 | tryToRead_7[30] & input_30_valid_0
    | tryToRead_7[31] & input_31_valid_0;
  wire        selectReq_7_ready =
    tryToRead_7[0] & input_0_ready_0 | tryToRead_7[1] & input_1_ready_0 | tryToRead_7[2] & input_2_ready_0 | tryToRead_7[3] & input_3_ready_0 | tryToRead_7[4] & input_4_ready_0 | tryToRead_7[5] & input_5_ready_0 | tryToRead_7[6]
    & input_6_ready_0 | tryToRead_7[7] & input_7_ready_0 | tryToRead_7[8] & input_8_ready_0 | tryToRead_7[9] & input_9_ready_0 | tryToRead_7[10] & input_10_ready_0 | tryToRead_7[11] & input_11_ready_0 | tryToRead_7[12] & input_12_ready_0
    | tryToRead_7[13] & input_13_ready_0 | tryToRead_7[14] & input_14_ready_0 | tryToRead_7[15] & input_15_ready_0 | tryToRead_7[16] & input_16_ready_0 | tryToRead_7[17] & input_17_ready_0 | tryToRead_7[18] & input_18_ready_0
    | tryToRead_7[19] & input_19_ready_0 | tryToRead_7[20] & input_20_ready_0 | tryToRead_7[21] & input_21_ready_0 | tryToRead_7[22] & input_22_ready_0 | tryToRead_7[23] & input_23_ready_0 | tryToRead_7[24] & input_24_ready_0
    | tryToRead_7[25] & input_25_ready_0 | tryToRead_7[26] & input_26_ready_0 | tryToRead_7[27] & input_27_ready_0 | tryToRead_7[28] & input_28_ready_0 | tryToRead_7[29] & input_29_ready_0 | tryToRead_7[30] & input_30_ready_0
    | tryToRead_7[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_8 = {inputSelect1H_1[8], inputSelect1H_0[8]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_8 = {inputSelect1H_3[8], inputSelect1H_2[8]};
  wire [3:0]  tryToRead_lo_lo_lo_8 = {tryToRead_lo_lo_lo_hi_8, tryToRead_lo_lo_lo_lo_8};
  wire [1:0]  tryToRead_lo_lo_hi_lo_8 = {inputSelect1H_5[8], inputSelect1H_4[8]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_8 = {inputSelect1H_7[8], inputSelect1H_6[8]};
  wire [3:0]  tryToRead_lo_lo_hi_8 = {tryToRead_lo_lo_hi_hi_8, tryToRead_lo_lo_hi_lo_8};
  wire [7:0]  tryToRead_lo_lo_8 = {tryToRead_lo_lo_hi_8, tryToRead_lo_lo_lo_8};
  wire [1:0]  tryToRead_lo_hi_lo_lo_8 = {inputSelect1H_9[8], inputSelect1H_8[8]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_8 = {inputSelect1H_11[8], inputSelect1H_10[8]};
  wire [3:0]  tryToRead_lo_hi_lo_8 = {tryToRead_lo_hi_lo_hi_8, tryToRead_lo_hi_lo_lo_8};
  wire [1:0]  tryToRead_lo_hi_hi_lo_8 = {inputSelect1H_13[8], inputSelect1H_12[8]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_8 = {inputSelect1H_15[8], inputSelect1H_14[8]};
  wire [3:0]  tryToRead_lo_hi_hi_8 = {tryToRead_lo_hi_hi_hi_8, tryToRead_lo_hi_hi_lo_8};
  wire [7:0]  tryToRead_lo_hi_8 = {tryToRead_lo_hi_hi_8, tryToRead_lo_hi_lo_8};
  wire [15:0] tryToRead_lo_8 = {tryToRead_lo_hi_8, tryToRead_lo_lo_8};
  wire [1:0]  tryToRead_hi_lo_lo_lo_8 = {inputSelect1H_17[8], inputSelect1H_16[8]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_8 = {inputSelect1H_19[8], inputSelect1H_18[8]};
  wire [3:0]  tryToRead_hi_lo_lo_8 = {tryToRead_hi_lo_lo_hi_8, tryToRead_hi_lo_lo_lo_8};
  wire [1:0]  tryToRead_hi_lo_hi_lo_8 = {inputSelect1H_21[8], inputSelect1H_20[8]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_8 = {inputSelect1H_23[8], inputSelect1H_22[8]};
  wire [3:0]  tryToRead_hi_lo_hi_8 = {tryToRead_hi_lo_hi_hi_8, tryToRead_hi_lo_hi_lo_8};
  wire [7:0]  tryToRead_hi_lo_8 = {tryToRead_hi_lo_hi_8, tryToRead_hi_lo_lo_8};
  wire [1:0]  tryToRead_hi_hi_lo_lo_8 = {inputSelect1H_25[8], inputSelect1H_24[8]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_8 = {inputSelect1H_27[8], inputSelect1H_26[8]};
  wire [3:0]  tryToRead_hi_hi_lo_8 = {tryToRead_hi_hi_lo_hi_8, tryToRead_hi_hi_lo_lo_8};
  wire [1:0]  tryToRead_hi_hi_hi_lo_8 = {inputSelect1H_29[8], inputSelect1H_28[8]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_8 = {inputSelect1H_31[8], inputSelect1H_30[8]};
  wire [3:0]  tryToRead_hi_hi_hi_8 = {tryToRead_hi_hi_hi_hi_8, tryToRead_hi_hi_hi_lo_8};
  wire [7:0]  tryToRead_hi_hi_8 = {tryToRead_hi_hi_hi_8, tryToRead_hi_hi_lo_8};
  wire [15:0] tryToRead_hi_8 = {tryToRead_hi_hi_8, tryToRead_hi_lo_8};
  wire [31:0] tryToRead_8 = {tryToRead_hi_8, tryToRead_lo_8};
  wire        output_8_valid_0 = |tryToRead_8;
  wire [4:0]  output_8_bits_vs_0 = selectReq_8_bits_vs;
  wire        output_8_bits_offset_0 = selectReq_8_bits_offset;
  wire [4:0]  output_8_bits_writeIndex_0 = selectReq_8_bits_requestIndex;
  wire [1:0]  output_8_bits_dataOffset_0 = selectReq_8_bits_dataOffset;
  assign selectReq_8_bits_dataOffset =
    (tryToRead_8[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_8[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_8[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_8[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_8[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_8[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_8[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_8[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_8[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_8[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_8[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_8[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_8[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_8[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_8[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_8[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_8[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_8[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_8[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_8[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_8[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_8[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_8[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_8[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_8[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_8_bits_requestIndex =
    {4'h0, tryToRead_8[1]} | {3'h0, tryToRead_8[2], 1'h0} | (tryToRead_8[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_8[4], 2'h0} | (tryToRead_8[5] ? 5'h5 : 5'h0) | (tryToRead_8[6] ? 5'h6 : 5'h0) | (tryToRead_8[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_8[8], 3'h0} | (tryToRead_8[9] ? 5'h9 : 5'h0) | (tryToRead_8[10] ? 5'hA : 5'h0) | (tryToRead_8[11] ? 5'hB : 5'h0) | (tryToRead_8[12] ? 5'hC : 5'h0) | (tryToRead_8[13] ? 5'hD : 5'h0) | (tryToRead_8[14] ? 5'hE : 5'h0)
    | (tryToRead_8[15] ? 5'hF : 5'h0) | {tryToRead_8[16], 4'h0} | (tryToRead_8[17] ? 5'h11 : 5'h0) | (tryToRead_8[18] ? 5'h12 : 5'h0) | (tryToRead_8[19] ? 5'h13 : 5'h0) | (tryToRead_8[20] ? 5'h14 : 5'h0) | (tryToRead_8[21] ? 5'h15 : 5'h0)
    | (tryToRead_8[22] ? 5'h16 : 5'h0) | (tryToRead_8[23] ? 5'h17 : 5'h0) | (tryToRead_8[24] ? 5'h18 : 5'h0) | (tryToRead_8[25] ? 5'h19 : 5'h0) | (tryToRead_8[26] ? 5'h1A : 5'h0) | (tryToRead_8[27] ? 5'h1B : 5'h0)
    | (tryToRead_8[28] ? 5'h1C : 5'h0) | (tryToRead_8[29] ? 5'h1D : 5'h0) | (tryToRead_8[30] ? 5'h1E : 5'h0) | {5{tryToRead_8[31]}};
  wire [4:0]  selectReq_8_bits_readLane =
    (tryToRead_8[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_8[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_8[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_8[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_8[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_8[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_8[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_8[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_8[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_8[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_8[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_8[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_8[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_8[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_8[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_8[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_8[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_8[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_8[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_8[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_8[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_8[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_8[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_8[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_8[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_8[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_8[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_8[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_8[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_8[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_8[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_8[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_8_bits_offset =
    tryToRead_8[0] & input_0_bits_offset_0 | tryToRead_8[1] & input_1_bits_offset_0 | tryToRead_8[2] & input_2_bits_offset_0 | tryToRead_8[3] & input_3_bits_offset_0 | tryToRead_8[4] & input_4_bits_offset_0 | tryToRead_8[5]
    & input_5_bits_offset_0 | tryToRead_8[6] & input_6_bits_offset_0 | tryToRead_8[7] & input_7_bits_offset_0 | tryToRead_8[8] & input_8_bits_offset_0 | tryToRead_8[9] & input_9_bits_offset_0 | tryToRead_8[10] & input_10_bits_offset_0
    | tryToRead_8[11] & input_11_bits_offset_0 | tryToRead_8[12] & input_12_bits_offset_0 | tryToRead_8[13] & input_13_bits_offset_0 | tryToRead_8[14] & input_14_bits_offset_0 | tryToRead_8[15] & input_15_bits_offset_0 | tryToRead_8[16]
    & input_16_bits_offset_0 | tryToRead_8[17] & input_17_bits_offset_0 | tryToRead_8[18] & input_18_bits_offset_0 | tryToRead_8[19] & input_19_bits_offset_0 | tryToRead_8[20] & input_20_bits_offset_0 | tryToRead_8[21]
    & input_21_bits_offset_0 | tryToRead_8[22] & input_22_bits_offset_0 | tryToRead_8[23] & input_23_bits_offset_0 | tryToRead_8[24] & input_24_bits_offset_0 | tryToRead_8[25] & input_25_bits_offset_0 | tryToRead_8[26]
    & input_26_bits_offset_0 | tryToRead_8[27] & input_27_bits_offset_0 | tryToRead_8[28] & input_28_bits_offset_0 | tryToRead_8[29] & input_29_bits_offset_0 | tryToRead_8[30] & input_30_bits_offset_0 | tryToRead_8[31]
    & input_31_bits_offset_0;
  assign selectReq_8_bits_vs =
    (tryToRead_8[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_8[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_8[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_8[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_8[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_8[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_8[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_8[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_8[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_8[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_8[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_8[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_8[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_8[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_8[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_8[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_8[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_8[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_8[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_8[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_8[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_8[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_8[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_8[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_8[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_8[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_8[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_8[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_8[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_8[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_8[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_8[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_8_valid =
    tryToRead_8[0] & input_0_valid_0 | tryToRead_8[1] & input_1_valid_0 | tryToRead_8[2] & input_2_valid_0 | tryToRead_8[3] & input_3_valid_0 | tryToRead_8[4] & input_4_valid_0 | tryToRead_8[5] & input_5_valid_0 | tryToRead_8[6]
    & input_6_valid_0 | tryToRead_8[7] & input_7_valid_0 | tryToRead_8[8] & input_8_valid_0 | tryToRead_8[9] & input_9_valid_0 | tryToRead_8[10] & input_10_valid_0 | tryToRead_8[11] & input_11_valid_0 | tryToRead_8[12] & input_12_valid_0
    | tryToRead_8[13] & input_13_valid_0 | tryToRead_8[14] & input_14_valid_0 | tryToRead_8[15] & input_15_valid_0 | tryToRead_8[16] & input_16_valid_0 | tryToRead_8[17] & input_17_valid_0 | tryToRead_8[18] & input_18_valid_0
    | tryToRead_8[19] & input_19_valid_0 | tryToRead_8[20] & input_20_valid_0 | tryToRead_8[21] & input_21_valid_0 | tryToRead_8[22] & input_22_valid_0 | tryToRead_8[23] & input_23_valid_0 | tryToRead_8[24] & input_24_valid_0
    | tryToRead_8[25] & input_25_valid_0 | tryToRead_8[26] & input_26_valid_0 | tryToRead_8[27] & input_27_valid_0 | tryToRead_8[28] & input_28_valid_0 | tryToRead_8[29] & input_29_valid_0 | tryToRead_8[30] & input_30_valid_0
    | tryToRead_8[31] & input_31_valid_0;
  wire        selectReq_8_ready =
    tryToRead_8[0] & input_0_ready_0 | tryToRead_8[1] & input_1_ready_0 | tryToRead_8[2] & input_2_ready_0 | tryToRead_8[3] & input_3_ready_0 | tryToRead_8[4] & input_4_ready_0 | tryToRead_8[5] & input_5_ready_0 | tryToRead_8[6]
    & input_6_ready_0 | tryToRead_8[7] & input_7_ready_0 | tryToRead_8[8] & input_8_ready_0 | tryToRead_8[9] & input_9_ready_0 | tryToRead_8[10] & input_10_ready_0 | tryToRead_8[11] & input_11_ready_0 | tryToRead_8[12] & input_12_ready_0
    | tryToRead_8[13] & input_13_ready_0 | tryToRead_8[14] & input_14_ready_0 | tryToRead_8[15] & input_15_ready_0 | tryToRead_8[16] & input_16_ready_0 | tryToRead_8[17] & input_17_ready_0 | tryToRead_8[18] & input_18_ready_0
    | tryToRead_8[19] & input_19_ready_0 | tryToRead_8[20] & input_20_ready_0 | tryToRead_8[21] & input_21_ready_0 | tryToRead_8[22] & input_22_ready_0 | tryToRead_8[23] & input_23_ready_0 | tryToRead_8[24] & input_24_ready_0
    | tryToRead_8[25] & input_25_ready_0 | tryToRead_8[26] & input_26_ready_0 | tryToRead_8[27] & input_27_ready_0 | tryToRead_8[28] & input_28_ready_0 | tryToRead_8[29] & input_29_ready_0 | tryToRead_8[30] & input_30_ready_0
    | tryToRead_8[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_9 = {inputSelect1H_1[9], inputSelect1H_0[9]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_9 = {inputSelect1H_3[9], inputSelect1H_2[9]};
  wire [3:0]  tryToRead_lo_lo_lo_9 = {tryToRead_lo_lo_lo_hi_9, tryToRead_lo_lo_lo_lo_9};
  wire [1:0]  tryToRead_lo_lo_hi_lo_9 = {inputSelect1H_5[9], inputSelect1H_4[9]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_9 = {inputSelect1H_7[9], inputSelect1H_6[9]};
  wire [3:0]  tryToRead_lo_lo_hi_9 = {tryToRead_lo_lo_hi_hi_9, tryToRead_lo_lo_hi_lo_9};
  wire [7:0]  tryToRead_lo_lo_9 = {tryToRead_lo_lo_hi_9, tryToRead_lo_lo_lo_9};
  wire [1:0]  tryToRead_lo_hi_lo_lo_9 = {inputSelect1H_9[9], inputSelect1H_8[9]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_9 = {inputSelect1H_11[9], inputSelect1H_10[9]};
  wire [3:0]  tryToRead_lo_hi_lo_9 = {tryToRead_lo_hi_lo_hi_9, tryToRead_lo_hi_lo_lo_9};
  wire [1:0]  tryToRead_lo_hi_hi_lo_9 = {inputSelect1H_13[9], inputSelect1H_12[9]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_9 = {inputSelect1H_15[9], inputSelect1H_14[9]};
  wire [3:0]  tryToRead_lo_hi_hi_9 = {tryToRead_lo_hi_hi_hi_9, tryToRead_lo_hi_hi_lo_9};
  wire [7:0]  tryToRead_lo_hi_9 = {tryToRead_lo_hi_hi_9, tryToRead_lo_hi_lo_9};
  wire [15:0] tryToRead_lo_9 = {tryToRead_lo_hi_9, tryToRead_lo_lo_9};
  wire [1:0]  tryToRead_hi_lo_lo_lo_9 = {inputSelect1H_17[9], inputSelect1H_16[9]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_9 = {inputSelect1H_19[9], inputSelect1H_18[9]};
  wire [3:0]  tryToRead_hi_lo_lo_9 = {tryToRead_hi_lo_lo_hi_9, tryToRead_hi_lo_lo_lo_9};
  wire [1:0]  tryToRead_hi_lo_hi_lo_9 = {inputSelect1H_21[9], inputSelect1H_20[9]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_9 = {inputSelect1H_23[9], inputSelect1H_22[9]};
  wire [3:0]  tryToRead_hi_lo_hi_9 = {tryToRead_hi_lo_hi_hi_9, tryToRead_hi_lo_hi_lo_9};
  wire [7:0]  tryToRead_hi_lo_9 = {tryToRead_hi_lo_hi_9, tryToRead_hi_lo_lo_9};
  wire [1:0]  tryToRead_hi_hi_lo_lo_9 = {inputSelect1H_25[9], inputSelect1H_24[9]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_9 = {inputSelect1H_27[9], inputSelect1H_26[9]};
  wire [3:0]  tryToRead_hi_hi_lo_9 = {tryToRead_hi_hi_lo_hi_9, tryToRead_hi_hi_lo_lo_9};
  wire [1:0]  tryToRead_hi_hi_hi_lo_9 = {inputSelect1H_29[9], inputSelect1H_28[9]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_9 = {inputSelect1H_31[9], inputSelect1H_30[9]};
  wire [3:0]  tryToRead_hi_hi_hi_9 = {tryToRead_hi_hi_hi_hi_9, tryToRead_hi_hi_hi_lo_9};
  wire [7:0]  tryToRead_hi_hi_9 = {tryToRead_hi_hi_hi_9, tryToRead_hi_hi_lo_9};
  wire [15:0] tryToRead_hi_9 = {tryToRead_hi_hi_9, tryToRead_hi_lo_9};
  wire [31:0] tryToRead_9 = {tryToRead_hi_9, tryToRead_lo_9};
  wire        output_9_valid_0 = |tryToRead_9;
  wire [4:0]  output_9_bits_vs_0 = selectReq_9_bits_vs;
  wire        output_9_bits_offset_0 = selectReq_9_bits_offset;
  wire [4:0]  output_9_bits_writeIndex_0 = selectReq_9_bits_requestIndex;
  wire [1:0]  output_9_bits_dataOffset_0 = selectReq_9_bits_dataOffset;
  assign selectReq_9_bits_dataOffset =
    (tryToRead_9[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_9[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_9[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_9[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_9[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_9[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_9[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_9[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_9[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_9[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_9[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_9[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_9[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_9[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_9[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_9[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_9[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_9[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_9[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_9[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_9[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_9[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_9[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_9[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_9[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_9_bits_requestIndex =
    {4'h0, tryToRead_9[1]} | {3'h0, tryToRead_9[2], 1'h0} | (tryToRead_9[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_9[4], 2'h0} | (tryToRead_9[5] ? 5'h5 : 5'h0) | (tryToRead_9[6] ? 5'h6 : 5'h0) | (tryToRead_9[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_9[8], 3'h0} | (tryToRead_9[9] ? 5'h9 : 5'h0) | (tryToRead_9[10] ? 5'hA : 5'h0) | (tryToRead_9[11] ? 5'hB : 5'h0) | (tryToRead_9[12] ? 5'hC : 5'h0) | (tryToRead_9[13] ? 5'hD : 5'h0) | (tryToRead_9[14] ? 5'hE : 5'h0)
    | (tryToRead_9[15] ? 5'hF : 5'h0) | {tryToRead_9[16], 4'h0} | (tryToRead_9[17] ? 5'h11 : 5'h0) | (tryToRead_9[18] ? 5'h12 : 5'h0) | (tryToRead_9[19] ? 5'h13 : 5'h0) | (tryToRead_9[20] ? 5'h14 : 5'h0) | (tryToRead_9[21] ? 5'h15 : 5'h0)
    | (tryToRead_9[22] ? 5'h16 : 5'h0) | (tryToRead_9[23] ? 5'h17 : 5'h0) | (tryToRead_9[24] ? 5'h18 : 5'h0) | (tryToRead_9[25] ? 5'h19 : 5'h0) | (tryToRead_9[26] ? 5'h1A : 5'h0) | (tryToRead_9[27] ? 5'h1B : 5'h0)
    | (tryToRead_9[28] ? 5'h1C : 5'h0) | (tryToRead_9[29] ? 5'h1D : 5'h0) | (tryToRead_9[30] ? 5'h1E : 5'h0) | {5{tryToRead_9[31]}};
  wire [4:0]  selectReq_9_bits_readLane =
    (tryToRead_9[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_9[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_9[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_9[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_9[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_9[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_9[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_9[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_9[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_9[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_9[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_9[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_9[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_9[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_9[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_9[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_9[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_9[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_9[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_9[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_9[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_9[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_9[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_9[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_9[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_9[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_9[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_9[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_9[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_9[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_9[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_9[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_9_bits_offset =
    tryToRead_9[0] & input_0_bits_offset_0 | tryToRead_9[1] & input_1_bits_offset_0 | tryToRead_9[2] & input_2_bits_offset_0 | tryToRead_9[3] & input_3_bits_offset_0 | tryToRead_9[4] & input_4_bits_offset_0 | tryToRead_9[5]
    & input_5_bits_offset_0 | tryToRead_9[6] & input_6_bits_offset_0 | tryToRead_9[7] & input_7_bits_offset_0 | tryToRead_9[8] & input_8_bits_offset_0 | tryToRead_9[9] & input_9_bits_offset_0 | tryToRead_9[10] & input_10_bits_offset_0
    | tryToRead_9[11] & input_11_bits_offset_0 | tryToRead_9[12] & input_12_bits_offset_0 | tryToRead_9[13] & input_13_bits_offset_0 | tryToRead_9[14] & input_14_bits_offset_0 | tryToRead_9[15] & input_15_bits_offset_0 | tryToRead_9[16]
    & input_16_bits_offset_0 | tryToRead_9[17] & input_17_bits_offset_0 | tryToRead_9[18] & input_18_bits_offset_0 | tryToRead_9[19] & input_19_bits_offset_0 | tryToRead_9[20] & input_20_bits_offset_0 | tryToRead_9[21]
    & input_21_bits_offset_0 | tryToRead_9[22] & input_22_bits_offset_0 | tryToRead_9[23] & input_23_bits_offset_0 | tryToRead_9[24] & input_24_bits_offset_0 | tryToRead_9[25] & input_25_bits_offset_0 | tryToRead_9[26]
    & input_26_bits_offset_0 | tryToRead_9[27] & input_27_bits_offset_0 | tryToRead_9[28] & input_28_bits_offset_0 | tryToRead_9[29] & input_29_bits_offset_0 | tryToRead_9[30] & input_30_bits_offset_0 | tryToRead_9[31]
    & input_31_bits_offset_0;
  assign selectReq_9_bits_vs =
    (tryToRead_9[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_9[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_9[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_9[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_9[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_9[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_9[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_9[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_9[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_9[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_9[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_9[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_9[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_9[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_9[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_9[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_9[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_9[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_9[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_9[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_9[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_9[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_9[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_9[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_9[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_9[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_9[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_9[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_9[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_9[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_9[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_9[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_9_valid =
    tryToRead_9[0] & input_0_valid_0 | tryToRead_9[1] & input_1_valid_0 | tryToRead_9[2] & input_2_valid_0 | tryToRead_9[3] & input_3_valid_0 | tryToRead_9[4] & input_4_valid_0 | tryToRead_9[5] & input_5_valid_0 | tryToRead_9[6]
    & input_6_valid_0 | tryToRead_9[7] & input_7_valid_0 | tryToRead_9[8] & input_8_valid_0 | tryToRead_9[9] & input_9_valid_0 | tryToRead_9[10] & input_10_valid_0 | tryToRead_9[11] & input_11_valid_0 | tryToRead_9[12] & input_12_valid_0
    | tryToRead_9[13] & input_13_valid_0 | tryToRead_9[14] & input_14_valid_0 | tryToRead_9[15] & input_15_valid_0 | tryToRead_9[16] & input_16_valid_0 | tryToRead_9[17] & input_17_valid_0 | tryToRead_9[18] & input_18_valid_0
    | tryToRead_9[19] & input_19_valid_0 | tryToRead_9[20] & input_20_valid_0 | tryToRead_9[21] & input_21_valid_0 | tryToRead_9[22] & input_22_valid_0 | tryToRead_9[23] & input_23_valid_0 | tryToRead_9[24] & input_24_valid_0
    | tryToRead_9[25] & input_25_valid_0 | tryToRead_9[26] & input_26_valid_0 | tryToRead_9[27] & input_27_valid_0 | tryToRead_9[28] & input_28_valid_0 | tryToRead_9[29] & input_29_valid_0 | tryToRead_9[30] & input_30_valid_0
    | tryToRead_9[31] & input_31_valid_0;
  wire        selectReq_9_ready =
    tryToRead_9[0] & input_0_ready_0 | tryToRead_9[1] & input_1_ready_0 | tryToRead_9[2] & input_2_ready_0 | tryToRead_9[3] & input_3_ready_0 | tryToRead_9[4] & input_4_ready_0 | tryToRead_9[5] & input_5_ready_0 | tryToRead_9[6]
    & input_6_ready_0 | tryToRead_9[7] & input_7_ready_0 | tryToRead_9[8] & input_8_ready_0 | tryToRead_9[9] & input_9_ready_0 | tryToRead_9[10] & input_10_ready_0 | tryToRead_9[11] & input_11_ready_0 | tryToRead_9[12] & input_12_ready_0
    | tryToRead_9[13] & input_13_ready_0 | tryToRead_9[14] & input_14_ready_0 | tryToRead_9[15] & input_15_ready_0 | tryToRead_9[16] & input_16_ready_0 | tryToRead_9[17] & input_17_ready_0 | tryToRead_9[18] & input_18_ready_0
    | tryToRead_9[19] & input_19_ready_0 | tryToRead_9[20] & input_20_ready_0 | tryToRead_9[21] & input_21_ready_0 | tryToRead_9[22] & input_22_ready_0 | tryToRead_9[23] & input_23_ready_0 | tryToRead_9[24] & input_24_ready_0
    | tryToRead_9[25] & input_25_ready_0 | tryToRead_9[26] & input_26_ready_0 | tryToRead_9[27] & input_27_ready_0 | tryToRead_9[28] & input_28_ready_0 | tryToRead_9[29] & input_29_ready_0 | tryToRead_9[30] & input_30_ready_0
    | tryToRead_9[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_10 = {inputSelect1H_1[10], inputSelect1H_0[10]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_10 = {inputSelect1H_3[10], inputSelect1H_2[10]};
  wire [3:0]  tryToRead_lo_lo_lo_10 = {tryToRead_lo_lo_lo_hi_10, tryToRead_lo_lo_lo_lo_10};
  wire [1:0]  tryToRead_lo_lo_hi_lo_10 = {inputSelect1H_5[10], inputSelect1H_4[10]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_10 = {inputSelect1H_7[10], inputSelect1H_6[10]};
  wire [3:0]  tryToRead_lo_lo_hi_10 = {tryToRead_lo_lo_hi_hi_10, tryToRead_lo_lo_hi_lo_10};
  wire [7:0]  tryToRead_lo_lo_10 = {tryToRead_lo_lo_hi_10, tryToRead_lo_lo_lo_10};
  wire [1:0]  tryToRead_lo_hi_lo_lo_10 = {inputSelect1H_9[10], inputSelect1H_8[10]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_10 = {inputSelect1H_11[10], inputSelect1H_10[10]};
  wire [3:0]  tryToRead_lo_hi_lo_10 = {tryToRead_lo_hi_lo_hi_10, tryToRead_lo_hi_lo_lo_10};
  wire [1:0]  tryToRead_lo_hi_hi_lo_10 = {inputSelect1H_13[10], inputSelect1H_12[10]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_10 = {inputSelect1H_15[10], inputSelect1H_14[10]};
  wire [3:0]  tryToRead_lo_hi_hi_10 = {tryToRead_lo_hi_hi_hi_10, tryToRead_lo_hi_hi_lo_10};
  wire [7:0]  tryToRead_lo_hi_10 = {tryToRead_lo_hi_hi_10, tryToRead_lo_hi_lo_10};
  wire [15:0] tryToRead_lo_10 = {tryToRead_lo_hi_10, tryToRead_lo_lo_10};
  wire [1:0]  tryToRead_hi_lo_lo_lo_10 = {inputSelect1H_17[10], inputSelect1H_16[10]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_10 = {inputSelect1H_19[10], inputSelect1H_18[10]};
  wire [3:0]  tryToRead_hi_lo_lo_10 = {tryToRead_hi_lo_lo_hi_10, tryToRead_hi_lo_lo_lo_10};
  wire [1:0]  tryToRead_hi_lo_hi_lo_10 = {inputSelect1H_21[10], inputSelect1H_20[10]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_10 = {inputSelect1H_23[10], inputSelect1H_22[10]};
  wire [3:0]  tryToRead_hi_lo_hi_10 = {tryToRead_hi_lo_hi_hi_10, tryToRead_hi_lo_hi_lo_10};
  wire [7:0]  tryToRead_hi_lo_10 = {tryToRead_hi_lo_hi_10, tryToRead_hi_lo_lo_10};
  wire [1:0]  tryToRead_hi_hi_lo_lo_10 = {inputSelect1H_25[10], inputSelect1H_24[10]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_10 = {inputSelect1H_27[10], inputSelect1H_26[10]};
  wire [3:0]  tryToRead_hi_hi_lo_10 = {tryToRead_hi_hi_lo_hi_10, tryToRead_hi_hi_lo_lo_10};
  wire [1:0]  tryToRead_hi_hi_hi_lo_10 = {inputSelect1H_29[10], inputSelect1H_28[10]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_10 = {inputSelect1H_31[10], inputSelect1H_30[10]};
  wire [3:0]  tryToRead_hi_hi_hi_10 = {tryToRead_hi_hi_hi_hi_10, tryToRead_hi_hi_hi_lo_10};
  wire [7:0]  tryToRead_hi_hi_10 = {tryToRead_hi_hi_hi_10, tryToRead_hi_hi_lo_10};
  wire [15:0] tryToRead_hi_10 = {tryToRead_hi_hi_10, tryToRead_hi_lo_10};
  wire [31:0] tryToRead_10 = {tryToRead_hi_10, tryToRead_lo_10};
  wire        output_10_valid_0 = |tryToRead_10;
  wire [4:0]  output_10_bits_vs_0 = selectReq_10_bits_vs;
  wire        output_10_bits_offset_0 = selectReq_10_bits_offset;
  wire [4:0]  output_10_bits_writeIndex_0 = selectReq_10_bits_requestIndex;
  wire [1:0]  output_10_bits_dataOffset_0 = selectReq_10_bits_dataOffset;
  assign selectReq_10_bits_dataOffset =
    (tryToRead_10[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_10[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_10[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_10[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_10[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_10[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_10[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_10[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_10[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_10[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_10[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_10[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_10[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_10[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_10[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_10[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_10[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_10[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_10[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_10[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_10[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_10[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_10[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_10[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_10[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_10_bits_requestIndex =
    {4'h0, tryToRead_10[1]} | {3'h0, tryToRead_10[2], 1'h0} | (tryToRead_10[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_10[4], 2'h0} | (tryToRead_10[5] ? 5'h5 : 5'h0) | (tryToRead_10[6] ? 5'h6 : 5'h0) | (tryToRead_10[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_10[8], 3'h0} | (tryToRead_10[9] ? 5'h9 : 5'h0) | (tryToRead_10[10] ? 5'hA : 5'h0) | (tryToRead_10[11] ? 5'hB : 5'h0) | (tryToRead_10[12] ? 5'hC : 5'h0) | (tryToRead_10[13] ? 5'hD : 5'h0)
    | (tryToRead_10[14] ? 5'hE : 5'h0) | (tryToRead_10[15] ? 5'hF : 5'h0) | {tryToRead_10[16], 4'h0} | (tryToRead_10[17] ? 5'h11 : 5'h0) | (tryToRead_10[18] ? 5'h12 : 5'h0) | (tryToRead_10[19] ? 5'h13 : 5'h0)
    | (tryToRead_10[20] ? 5'h14 : 5'h0) | (tryToRead_10[21] ? 5'h15 : 5'h0) | (tryToRead_10[22] ? 5'h16 : 5'h0) | (tryToRead_10[23] ? 5'h17 : 5'h0) | (tryToRead_10[24] ? 5'h18 : 5'h0) | (tryToRead_10[25] ? 5'h19 : 5'h0)
    | (tryToRead_10[26] ? 5'h1A : 5'h0) | (tryToRead_10[27] ? 5'h1B : 5'h0) | (tryToRead_10[28] ? 5'h1C : 5'h0) | (tryToRead_10[29] ? 5'h1D : 5'h0) | (tryToRead_10[30] ? 5'h1E : 5'h0) | {5{tryToRead_10[31]}};
  wire [4:0]  selectReq_10_bits_readLane =
    (tryToRead_10[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_10[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_10[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_10[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_10[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_10[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_10[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_10[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_10[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_10[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_10[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_10[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_10[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_10[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_10[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_10[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_10[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_10[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_10[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_10[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_10[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_10[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_10[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_10[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_10[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_10[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_10[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_10[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_10[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_10[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_10[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_10[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_10_bits_offset =
    tryToRead_10[0] & input_0_bits_offset_0 | tryToRead_10[1] & input_1_bits_offset_0 | tryToRead_10[2] & input_2_bits_offset_0 | tryToRead_10[3] & input_3_bits_offset_0 | tryToRead_10[4] & input_4_bits_offset_0 | tryToRead_10[5]
    & input_5_bits_offset_0 | tryToRead_10[6] & input_6_bits_offset_0 | tryToRead_10[7] & input_7_bits_offset_0 | tryToRead_10[8] & input_8_bits_offset_0 | tryToRead_10[9] & input_9_bits_offset_0 | tryToRead_10[10] & input_10_bits_offset_0
    | tryToRead_10[11] & input_11_bits_offset_0 | tryToRead_10[12] & input_12_bits_offset_0 | tryToRead_10[13] & input_13_bits_offset_0 | tryToRead_10[14] & input_14_bits_offset_0 | tryToRead_10[15] & input_15_bits_offset_0
    | tryToRead_10[16] & input_16_bits_offset_0 | tryToRead_10[17] & input_17_bits_offset_0 | tryToRead_10[18] & input_18_bits_offset_0 | tryToRead_10[19] & input_19_bits_offset_0 | tryToRead_10[20] & input_20_bits_offset_0
    | tryToRead_10[21] & input_21_bits_offset_0 | tryToRead_10[22] & input_22_bits_offset_0 | tryToRead_10[23] & input_23_bits_offset_0 | tryToRead_10[24] & input_24_bits_offset_0 | tryToRead_10[25] & input_25_bits_offset_0
    | tryToRead_10[26] & input_26_bits_offset_0 | tryToRead_10[27] & input_27_bits_offset_0 | tryToRead_10[28] & input_28_bits_offset_0 | tryToRead_10[29] & input_29_bits_offset_0 | tryToRead_10[30] & input_30_bits_offset_0
    | tryToRead_10[31] & input_31_bits_offset_0;
  assign selectReq_10_bits_vs =
    (tryToRead_10[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_10[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_10[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_10[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_10[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_10[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_10[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_10[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_10[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_10[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_10[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_10[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_10[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_10[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_10[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_10[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_10[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_10[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_10[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_10[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_10[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_10[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_10[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_10[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_10[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_10[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_10[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_10[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_10[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_10[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_10[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_10[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_10_valid =
    tryToRead_10[0] & input_0_valid_0 | tryToRead_10[1] & input_1_valid_0 | tryToRead_10[2] & input_2_valid_0 | tryToRead_10[3] & input_3_valid_0 | tryToRead_10[4] & input_4_valid_0 | tryToRead_10[5] & input_5_valid_0 | tryToRead_10[6]
    & input_6_valid_0 | tryToRead_10[7] & input_7_valid_0 | tryToRead_10[8] & input_8_valid_0 | tryToRead_10[9] & input_9_valid_0 | tryToRead_10[10] & input_10_valid_0 | tryToRead_10[11] & input_11_valid_0 | tryToRead_10[12]
    & input_12_valid_0 | tryToRead_10[13] & input_13_valid_0 | tryToRead_10[14] & input_14_valid_0 | tryToRead_10[15] & input_15_valid_0 | tryToRead_10[16] & input_16_valid_0 | tryToRead_10[17] & input_17_valid_0 | tryToRead_10[18]
    & input_18_valid_0 | tryToRead_10[19] & input_19_valid_0 | tryToRead_10[20] & input_20_valid_0 | tryToRead_10[21] & input_21_valid_0 | tryToRead_10[22] & input_22_valid_0 | tryToRead_10[23] & input_23_valid_0 | tryToRead_10[24]
    & input_24_valid_0 | tryToRead_10[25] & input_25_valid_0 | tryToRead_10[26] & input_26_valid_0 | tryToRead_10[27] & input_27_valid_0 | tryToRead_10[28] & input_28_valid_0 | tryToRead_10[29] & input_29_valid_0 | tryToRead_10[30]
    & input_30_valid_0 | tryToRead_10[31] & input_31_valid_0;
  wire        selectReq_10_ready =
    tryToRead_10[0] & input_0_ready_0 | tryToRead_10[1] & input_1_ready_0 | tryToRead_10[2] & input_2_ready_0 | tryToRead_10[3] & input_3_ready_0 | tryToRead_10[4] & input_4_ready_0 | tryToRead_10[5] & input_5_ready_0 | tryToRead_10[6]
    & input_6_ready_0 | tryToRead_10[7] & input_7_ready_0 | tryToRead_10[8] & input_8_ready_0 | tryToRead_10[9] & input_9_ready_0 | tryToRead_10[10] & input_10_ready_0 | tryToRead_10[11] & input_11_ready_0 | tryToRead_10[12]
    & input_12_ready_0 | tryToRead_10[13] & input_13_ready_0 | tryToRead_10[14] & input_14_ready_0 | tryToRead_10[15] & input_15_ready_0 | tryToRead_10[16] & input_16_ready_0 | tryToRead_10[17] & input_17_ready_0 | tryToRead_10[18]
    & input_18_ready_0 | tryToRead_10[19] & input_19_ready_0 | tryToRead_10[20] & input_20_ready_0 | tryToRead_10[21] & input_21_ready_0 | tryToRead_10[22] & input_22_ready_0 | tryToRead_10[23] & input_23_ready_0 | tryToRead_10[24]
    & input_24_ready_0 | tryToRead_10[25] & input_25_ready_0 | tryToRead_10[26] & input_26_ready_0 | tryToRead_10[27] & input_27_ready_0 | tryToRead_10[28] & input_28_ready_0 | tryToRead_10[29] & input_29_ready_0 | tryToRead_10[30]
    & input_30_ready_0 | tryToRead_10[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_11 = {inputSelect1H_1[11], inputSelect1H_0[11]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_11 = {inputSelect1H_3[11], inputSelect1H_2[11]};
  wire [3:0]  tryToRead_lo_lo_lo_11 = {tryToRead_lo_lo_lo_hi_11, tryToRead_lo_lo_lo_lo_11};
  wire [1:0]  tryToRead_lo_lo_hi_lo_11 = {inputSelect1H_5[11], inputSelect1H_4[11]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_11 = {inputSelect1H_7[11], inputSelect1H_6[11]};
  wire [3:0]  tryToRead_lo_lo_hi_11 = {tryToRead_lo_lo_hi_hi_11, tryToRead_lo_lo_hi_lo_11};
  wire [7:0]  tryToRead_lo_lo_11 = {tryToRead_lo_lo_hi_11, tryToRead_lo_lo_lo_11};
  wire [1:0]  tryToRead_lo_hi_lo_lo_11 = {inputSelect1H_9[11], inputSelect1H_8[11]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_11 = {inputSelect1H_11[11], inputSelect1H_10[11]};
  wire [3:0]  tryToRead_lo_hi_lo_11 = {tryToRead_lo_hi_lo_hi_11, tryToRead_lo_hi_lo_lo_11};
  wire [1:0]  tryToRead_lo_hi_hi_lo_11 = {inputSelect1H_13[11], inputSelect1H_12[11]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_11 = {inputSelect1H_15[11], inputSelect1H_14[11]};
  wire [3:0]  tryToRead_lo_hi_hi_11 = {tryToRead_lo_hi_hi_hi_11, tryToRead_lo_hi_hi_lo_11};
  wire [7:0]  tryToRead_lo_hi_11 = {tryToRead_lo_hi_hi_11, tryToRead_lo_hi_lo_11};
  wire [15:0] tryToRead_lo_11 = {tryToRead_lo_hi_11, tryToRead_lo_lo_11};
  wire [1:0]  tryToRead_hi_lo_lo_lo_11 = {inputSelect1H_17[11], inputSelect1H_16[11]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_11 = {inputSelect1H_19[11], inputSelect1H_18[11]};
  wire [3:0]  tryToRead_hi_lo_lo_11 = {tryToRead_hi_lo_lo_hi_11, tryToRead_hi_lo_lo_lo_11};
  wire [1:0]  tryToRead_hi_lo_hi_lo_11 = {inputSelect1H_21[11], inputSelect1H_20[11]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_11 = {inputSelect1H_23[11], inputSelect1H_22[11]};
  wire [3:0]  tryToRead_hi_lo_hi_11 = {tryToRead_hi_lo_hi_hi_11, tryToRead_hi_lo_hi_lo_11};
  wire [7:0]  tryToRead_hi_lo_11 = {tryToRead_hi_lo_hi_11, tryToRead_hi_lo_lo_11};
  wire [1:0]  tryToRead_hi_hi_lo_lo_11 = {inputSelect1H_25[11], inputSelect1H_24[11]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_11 = {inputSelect1H_27[11], inputSelect1H_26[11]};
  wire [3:0]  tryToRead_hi_hi_lo_11 = {tryToRead_hi_hi_lo_hi_11, tryToRead_hi_hi_lo_lo_11};
  wire [1:0]  tryToRead_hi_hi_hi_lo_11 = {inputSelect1H_29[11], inputSelect1H_28[11]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_11 = {inputSelect1H_31[11], inputSelect1H_30[11]};
  wire [3:0]  tryToRead_hi_hi_hi_11 = {tryToRead_hi_hi_hi_hi_11, tryToRead_hi_hi_hi_lo_11};
  wire [7:0]  tryToRead_hi_hi_11 = {tryToRead_hi_hi_hi_11, tryToRead_hi_hi_lo_11};
  wire [15:0] tryToRead_hi_11 = {tryToRead_hi_hi_11, tryToRead_hi_lo_11};
  wire [31:0] tryToRead_11 = {tryToRead_hi_11, tryToRead_lo_11};
  wire        output_11_valid_0 = |tryToRead_11;
  wire [4:0]  output_11_bits_vs_0 = selectReq_11_bits_vs;
  wire        output_11_bits_offset_0 = selectReq_11_bits_offset;
  wire [4:0]  output_11_bits_writeIndex_0 = selectReq_11_bits_requestIndex;
  wire [1:0]  output_11_bits_dataOffset_0 = selectReq_11_bits_dataOffset;
  assign selectReq_11_bits_dataOffset =
    (tryToRead_11[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_11[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_11[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_11[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_11[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_11[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_11[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_11[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_11[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_11[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_11[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_11[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_11[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_11[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_11[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_11[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_11[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_11[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_11[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_11[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_11[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_11[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_11[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_11[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_11[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_11_bits_requestIndex =
    {4'h0, tryToRead_11[1]} | {3'h0, tryToRead_11[2], 1'h0} | (tryToRead_11[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_11[4], 2'h0} | (tryToRead_11[5] ? 5'h5 : 5'h0) | (tryToRead_11[6] ? 5'h6 : 5'h0) | (tryToRead_11[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_11[8], 3'h0} | (tryToRead_11[9] ? 5'h9 : 5'h0) | (tryToRead_11[10] ? 5'hA : 5'h0) | (tryToRead_11[11] ? 5'hB : 5'h0) | (tryToRead_11[12] ? 5'hC : 5'h0) | (tryToRead_11[13] ? 5'hD : 5'h0)
    | (tryToRead_11[14] ? 5'hE : 5'h0) | (tryToRead_11[15] ? 5'hF : 5'h0) | {tryToRead_11[16], 4'h0} | (tryToRead_11[17] ? 5'h11 : 5'h0) | (tryToRead_11[18] ? 5'h12 : 5'h0) | (tryToRead_11[19] ? 5'h13 : 5'h0)
    | (tryToRead_11[20] ? 5'h14 : 5'h0) | (tryToRead_11[21] ? 5'h15 : 5'h0) | (tryToRead_11[22] ? 5'h16 : 5'h0) | (tryToRead_11[23] ? 5'h17 : 5'h0) | (tryToRead_11[24] ? 5'h18 : 5'h0) | (tryToRead_11[25] ? 5'h19 : 5'h0)
    | (tryToRead_11[26] ? 5'h1A : 5'h0) | (tryToRead_11[27] ? 5'h1B : 5'h0) | (tryToRead_11[28] ? 5'h1C : 5'h0) | (tryToRead_11[29] ? 5'h1D : 5'h0) | (tryToRead_11[30] ? 5'h1E : 5'h0) | {5{tryToRead_11[31]}};
  wire [4:0]  selectReq_11_bits_readLane =
    (tryToRead_11[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_11[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_11[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_11[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_11[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_11[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_11[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_11[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_11[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_11[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_11[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_11[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_11[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_11[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_11[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_11[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_11[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_11[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_11[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_11[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_11[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_11[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_11[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_11[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_11[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_11[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_11[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_11[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_11[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_11[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_11[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_11[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_11_bits_offset =
    tryToRead_11[0] & input_0_bits_offset_0 | tryToRead_11[1] & input_1_bits_offset_0 | tryToRead_11[2] & input_2_bits_offset_0 | tryToRead_11[3] & input_3_bits_offset_0 | tryToRead_11[4] & input_4_bits_offset_0 | tryToRead_11[5]
    & input_5_bits_offset_0 | tryToRead_11[6] & input_6_bits_offset_0 | tryToRead_11[7] & input_7_bits_offset_0 | tryToRead_11[8] & input_8_bits_offset_0 | tryToRead_11[9] & input_9_bits_offset_0 | tryToRead_11[10] & input_10_bits_offset_0
    | tryToRead_11[11] & input_11_bits_offset_0 | tryToRead_11[12] & input_12_bits_offset_0 | tryToRead_11[13] & input_13_bits_offset_0 | tryToRead_11[14] & input_14_bits_offset_0 | tryToRead_11[15] & input_15_bits_offset_0
    | tryToRead_11[16] & input_16_bits_offset_0 | tryToRead_11[17] & input_17_bits_offset_0 | tryToRead_11[18] & input_18_bits_offset_0 | tryToRead_11[19] & input_19_bits_offset_0 | tryToRead_11[20] & input_20_bits_offset_0
    | tryToRead_11[21] & input_21_bits_offset_0 | tryToRead_11[22] & input_22_bits_offset_0 | tryToRead_11[23] & input_23_bits_offset_0 | tryToRead_11[24] & input_24_bits_offset_0 | tryToRead_11[25] & input_25_bits_offset_0
    | tryToRead_11[26] & input_26_bits_offset_0 | tryToRead_11[27] & input_27_bits_offset_0 | tryToRead_11[28] & input_28_bits_offset_0 | tryToRead_11[29] & input_29_bits_offset_0 | tryToRead_11[30] & input_30_bits_offset_0
    | tryToRead_11[31] & input_31_bits_offset_0;
  assign selectReq_11_bits_vs =
    (tryToRead_11[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_11[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_11[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_11[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_11[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_11[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_11[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_11[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_11[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_11[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_11[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_11[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_11[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_11[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_11[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_11[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_11[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_11[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_11[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_11[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_11[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_11[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_11[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_11[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_11[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_11[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_11[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_11[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_11[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_11[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_11[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_11[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_11_valid =
    tryToRead_11[0] & input_0_valid_0 | tryToRead_11[1] & input_1_valid_0 | tryToRead_11[2] & input_2_valid_0 | tryToRead_11[3] & input_3_valid_0 | tryToRead_11[4] & input_4_valid_0 | tryToRead_11[5] & input_5_valid_0 | tryToRead_11[6]
    & input_6_valid_0 | tryToRead_11[7] & input_7_valid_0 | tryToRead_11[8] & input_8_valid_0 | tryToRead_11[9] & input_9_valid_0 | tryToRead_11[10] & input_10_valid_0 | tryToRead_11[11] & input_11_valid_0 | tryToRead_11[12]
    & input_12_valid_0 | tryToRead_11[13] & input_13_valid_0 | tryToRead_11[14] & input_14_valid_0 | tryToRead_11[15] & input_15_valid_0 | tryToRead_11[16] & input_16_valid_0 | tryToRead_11[17] & input_17_valid_0 | tryToRead_11[18]
    & input_18_valid_0 | tryToRead_11[19] & input_19_valid_0 | tryToRead_11[20] & input_20_valid_0 | tryToRead_11[21] & input_21_valid_0 | tryToRead_11[22] & input_22_valid_0 | tryToRead_11[23] & input_23_valid_0 | tryToRead_11[24]
    & input_24_valid_0 | tryToRead_11[25] & input_25_valid_0 | tryToRead_11[26] & input_26_valid_0 | tryToRead_11[27] & input_27_valid_0 | tryToRead_11[28] & input_28_valid_0 | tryToRead_11[29] & input_29_valid_0 | tryToRead_11[30]
    & input_30_valid_0 | tryToRead_11[31] & input_31_valid_0;
  wire        selectReq_11_ready =
    tryToRead_11[0] & input_0_ready_0 | tryToRead_11[1] & input_1_ready_0 | tryToRead_11[2] & input_2_ready_0 | tryToRead_11[3] & input_3_ready_0 | tryToRead_11[4] & input_4_ready_0 | tryToRead_11[5] & input_5_ready_0 | tryToRead_11[6]
    & input_6_ready_0 | tryToRead_11[7] & input_7_ready_0 | tryToRead_11[8] & input_8_ready_0 | tryToRead_11[9] & input_9_ready_0 | tryToRead_11[10] & input_10_ready_0 | tryToRead_11[11] & input_11_ready_0 | tryToRead_11[12]
    & input_12_ready_0 | tryToRead_11[13] & input_13_ready_0 | tryToRead_11[14] & input_14_ready_0 | tryToRead_11[15] & input_15_ready_0 | tryToRead_11[16] & input_16_ready_0 | tryToRead_11[17] & input_17_ready_0 | tryToRead_11[18]
    & input_18_ready_0 | tryToRead_11[19] & input_19_ready_0 | tryToRead_11[20] & input_20_ready_0 | tryToRead_11[21] & input_21_ready_0 | tryToRead_11[22] & input_22_ready_0 | tryToRead_11[23] & input_23_ready_0 | tryToRead_11[24]
    & input_24_ready_0 | tryToRead_11[25] & input_25_ready_0 | tryToRead_11[26] & input_26_ready_0 | tryToRead_11[27] & input_27_ready_0 | tryToRead_11[28] & input_28_ready_0 | tryToRead_11[29] & input_29_ready_0 | tryToRead_11[30]
    & input_30_ready_0 | tryToRead_11[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_12 = {inputSelect1H_1[12], inputSelect1H_0[12]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_12 = {inputSelect1H_3[12], inputSelect1H_2[12]};
  wire [3:0]  tryToRead_lo_lo_lo_12 = {tryToRead_lo_lo_lo_hi_12, tryToRead_lo_lo_lo_lo_12};
  wire [1:0]  tryToRead_lo_lo_hi_lo_12 = {inputSelect1H_5[12], inputSelect1H_4[12]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_12 = {inputSelect1H_7[12], inputSelect1H_6[12]};
  wire [3:0]  tryToRead_lo_lo_hi_12 = {tryToRead_lo_lo_hi_hi_12, tryToRead_lo_lo_hi_lo_12};
  wire [7:0]  tryToRead_lo_lo_12 = {tryToRead_lo_lo_hi_12, tryToRead_lo_lo_lo_12};
  wire [1:0]  tryToRead_lo_hi_lo_lo_12 = {inputSelect1H_9[12], inputSelect1H_8[12]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_12 = {inputSelect1H_11[12], inputSelect1H_10[12]};
  wire [3:0]  tryToRead_lo_hi_lo_12 = {tryToRead_lo_hi_lo_hi_12, tryToRead_lo_hi_lo_lo_12};
  wire [1:0]  tryToRead_lo_hi_hi_lo_12 = {inputSelect1H_13[12], inputSelect1H_12[12]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_12 = {inputSelect1H_15[12], inputSelect1H_14[12]};
  wire [3:0]  tryToRead_lo_hi_hi_12 = {tryToRead_lo_hi_hi_hi_12, tryToRead_lo_hi_hi_lo_12};
  wire [7:0]  tryToRead_lo_hi_12 = {tryToRead_lo_hi_hi_12, tryToRead_lo_hi_lo_12};
  wire [15:0] tryToRead_lo_12 = {tryToRead_lo_hi_12, tryToRead_lo_lo_12};
  wire [1:0]  tryToRead_hi_lo_lo_lo_12 = {inputSelect1H_17[12], inputSelect1H_16[12]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_12 = {inputSelect1H_19[12], inputSelect1H_18[12]};
  wire [3:0]  tryToRead_hi_lo_lo_12 = {tryToRead_hi_lo_lo_hi_12, tryToRead_hi_lo_lo_lo_12};
  wire [1:0]  tryToRead_hi_lo_hi_lo_12 = {inputSelect1H_21[12], inputSelect1H_20[12]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_12 = {inputSelect1H_23[12], inputSelect1H_22[12]};
  wire [3:0]  tryToRead_hi_lo_hi_12 = {tryToRead_hi_lo_hi_hi_12, tryToRead_hi_lo_hi_lo_12};
  wire [7:0]  tryToRead_hi_lo_12 = {tryToRead_hi_lo_hi_12, tryToRead_hi_lo_lo_12};
  wire [1:0]  tryToRead_hi_hi_lo_lo_12 = {inputSelect1H_25[12], inputSelect1H_24[12]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_12 = {inputSelect1H_27[12], inputSelect1H_26[12]};
  wire [3:0]  tryToRead_hi_hi_lo_12 = {tryToRead_hi_hi_lo_hi_12, tryToRead_hi_hi_lo_lo_12};
  wire [1:0]  tryToRead_hi_hi_hi_lo_12 = {inputSelect1H_29[12], inputSelect1H_28[12]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_12 = {inputSelect1H_31[12], inputSelect1H_30[12]};
  wire [3:0]  tryToRead_hi_hi_hi_12 = {tryToRead_hi_hi_hi_hi_12, tryToRead_hi_hi_hi_lo_12};
  wire [7:0]  tryToRead_hi_hi_12 = {tryToRead_hi_hi_hi_12, tryToRead_hi_hi_lo_12};
  wire [15:0] tryToRead_hi_12 = {tryToRead_hi_hi_12, tryToRead_hi_lo_12};
  wire [31:0] tryToRead_12 = {tryToRead_hi_12, tryToRead_lo_12};
  wire        output_12_valid_0 = |tryToRead_12;
  wire [4:0]  output_12_bits_vs_0 = selectReq_12_bits_vs;
  wire        output_12_bits_offset_0 = selectReq_12_bits_offset;
  wire [4:0]  output_12_bits_writeIndex_0 = selectReq_12_bits_requestIndex;
  wire [1:0]  output_12_bits_dataOffset_0 = selectReq_12_bits_dataOffset;
  assign selectReq_12_bits_dataOffset =
    (tryToRead_12[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_12[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_12[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_12[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_12[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_12[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_12[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_12[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_12[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_12[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_12[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_12[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_12[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_12[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_12[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_12[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_12[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_12[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_12[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_12[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_12[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_12[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_12[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_12[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_12[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_12_bits_requestIndex =
    {4'h0, tryToRead_12[1]} | {3'h0, tryToRead_12[2], 1'h0} | (tryToRead_12[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_12[4], 2'h0} | (tryToRead_12[5] ? 5'h5 : 5'h0) | (tryToRead_12[6] ? 5'h6 : 5'h0) | (tryToRead_12[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_12[8], 3'h0} | (tryToRead_12[9] ? 5'h9 : 5'h0) | (tryToRead_12[10] ? 5'hA : 5'h0) | (tryToRead_12[11] ? 5'hB : 5'h0) | (tryToRead_12[12] ? 5'hC : 5'h0) | (tryToRead_12[13] ? 5'hD : 5'h0)
    | (tryToRead_12[14] ? 5'hE : 5'h0) | (tryToRead_12[15] ? 5'hF : 5'h0) | {tryToRead_12[16], 4'h0} | (tryToRead_12[17] ? 5'h11 : 5'h0) | (tryToRead_12[18] ? 5'h12 : 5'h0) | (tryToRead_12[19] ? 5'h13 : 5'h0)
    | (tryToRead_12[20] ? 5'h14 : 5'h0) | (tryToRead_12[21] ? 5'h15 : 5'h0) | (tryToRead_12[22] ? 5'h16 : 5'h0) | (tryToRead_12[23] ? 5'h17 : 5'h0) | (tryToRead_12[24] ? 5'h18 : 5'h0) | (tryToRead_12[25] ? 5'h19 : 5'h0)
    | (tryToRead_12[26] ? 5'h1A : 5'h0) | (tryToRead_12[27] ? 5'h1B : 5'h0) | (tryToRead_12[28] ? 5'h1C : 5'h0) | (tryToRead_12[29] ? 5'h1D : 5'h0) | (tryToRead_12[30] ? 5'h1E : 5'h0) | {5{tryToRead_12[31]}};
  wire [4:0]  selectReq_12_bits_readLane =
    (tryToRead_12[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_12[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_12[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_12[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_12[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_12[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_12[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_12[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_12[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_12[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_12[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_12[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_12[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_12[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_12[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_12[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_12[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_12[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_12[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_12[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_12[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_12[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_12[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_12[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_12[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_12[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_12[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_12[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_12[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_12[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_12[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_12[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_12_bits_offset =
    tryToRead_12[0] & input_0_bits_offset_0 | tryToRead_12[1] & input_1_bits_offset_0 | tryToRead_12[2] & input_2_bits_offset_0 | tryToRead_12[3] & input_3_bits_offset_0 | tryToRead_12[4] & input_4_bits_offset_0 | tryToRead_12[5]
    & input_5_bits_offset_0 | tryToRead_12[6] & input_6_bits_offset_0 | tryToRead_12[7] & input_7_bits_offset_0 | tryToRead_12[8] & input_8_bits_offset_0 | tryToRead_12[9] & input_9_bits_offset_0 | tryToRead_12[10] & input_10_bits_offset_0
    | tryToRead_12[11] & input_11_bits_offset_0 | tryToRead_12[12] & input_12_bits_offset_0 | tryToRead_12[13] & input_13_bits_offset_0 | tryToRead_12[14] & input_14_bits_offset_0 | tryToRead_12[15] & input_15_bits_offset_0
    | tryToRead_12[16] & input_16_bits_offset_0 | tryToRead_12[17] & input_17_bits_offset_0 | tryToRead_12[18] & input_18_bits_offset_0 | tryToRead_12[19] & input_19_bits_offset_0 | tryToRead_12[20] & input_20_bits_offset_0
    | tryToRead_12[21] & input_21_bits_offset_0 | tryToRead_12[22] & input_22_bits_offset_0 | tryToRead_12[23] & input_23_bits_offset_0 | tryToRead_12[24] & input_24_bits_offset_0 | tryToRead_12[25] & input_25_bits_offset_0
    | tryToRead_12[26] & input_26_bits_offset_0 | tryToRead_12[27] & input_27_bits_offset_0 | tryToRead_12[28] & input_28_bits_offset_0 | tryToRead_12[29] & input_29_bits_offset_0 | tryToRead_12[30] & input_30_bits_offset_0
    | tryToRead_12[31] & input_31_bits_offset_0;
  assign selectReq_12_bits_vs =
    (tryToRead_12[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_12[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_12[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_12[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_12[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_12[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_12[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_12[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_12[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_12[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_12[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_12[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_12[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_12[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_12[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_12[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_12[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_12[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_12[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_12[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_12[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_12[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_12[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_12[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_12[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_12[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_12[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_12[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_12[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_12[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_12[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_12[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_12_valid =
    tryToRead_12[0] & input_0_valid_0 | tryToRead_12[1] & input_1_valid_0 | tryToRead_12[2] & input_2_valid_0 | tryToRead_12[3] & input_3_valid_0 | tryToRead_12[4] & input_4_valid_0 | tryToRead_12[5] & input_5_valid_0 | tryToRead_12[6]
    & input_6_valid_0 | tryToRead_12[7] & input_7_valid_0 | tryToRead_12[8] & input_8_valid_0 | tryToRead_12[9] & input_9_valid_0 | tryToRead_12[10] & input_10_valid_0 | tryToRead_12[11] & input_11_valid_0 | tryToRead_12[12]
    & input_12_valid_0 | tryToRead_12[13] & input_13_valid_0 | tryToRead_12[14] & input_14_valid_0 | tryToRead_12[15] & input_15_valid_0 | tryToRead_12[16] & input_16_valid_0 | tryToRead_12[17] & input_17_valid_0 | tryToRead_12[18]
    & input_18_valid_0 | tryToRead_12[19] & input_19_valid_0 | tryToRead_12[20] & input_20_valid_0 | tryToRead_12[21] & input_21_valid_0 | tryToRead_12[22] & input_22_valid_0 | tryToRead_12[23] & input_23_valid_0 | tryToRead_12[24]
    & input_24_valid_0 | tryToRead_12[25] & input_25_valid_0 | tryToRead_12[26] & input_26_valid_0 | tryToRead_12[27] & input_27_valid_0 | tryToRead_12[28] & input_28_valid_0 | tryToRead_12[29] & input_29_valid_0 | tryToRead_12[30]
    & input_30_valid_0 | tryToRead_12[31] & input_31_valid_0;
  wire        selectReq_12_ready =
    tryToRead_12[0] & input_0_ready_0 | tryToRead_12[1] & input_1_ready_0 | tryToRead_12[2] & input_2_ready_0 | tryToRead_12[3] & input_3_ready_0 | tryToRead_12[4] & input_4_ready_0 | tryToRead_12[5] & input_5_ready_0 | tryToRead_12[6]
    & input_6_ready_0 | tryToRead_12[7] & input_7_ready_0 | tryToRead_12[8] & input_8_ready_0 | tryToRead_12[9] & input_9_ready_0 | tryToRead_12[10] & input_10_ready_0 | tryToRead_12[11] & input_11_ready_0 | tryToRead_12[12]
    & input_12_ready_0 | tryToRead_12[13] & input_13_ready_0 | tryToRead_12[14] & input_14_ready_0 | tryToRead_12[15] & input_15_ready_0 | tryToRead_12[16] & input_16_ready_0 | tryToRead_12[17] & input_17_ready_0 | tryToRead_12[18]
    & input_18_ready_0 | tryToRead_12[19] & input_19_ready_0 | tryToRead_12[20] & input_20_ready_0 | tryToRead_12[21] & input_21_ready_0 | tryToRead_12[22] & input_22_ready_0 | tryToRead_12[23] & input_23_ready_0 | tryToRead_12[24]
    & input_24_ready_0 | tryToRead_12[25] & input_25_ready_0 | tryToRead_12[26] & input_26_ready_0 | tryToRead_12[27] & input_27_ready_0 | tryToRead_12[28] & input_28_ready_0 | tryToRead_12[29] & input_29_ready_0 | tryToRead_12[30]
    & input_30_ready_0 | tryToRead_12[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_13 = {inputSelect1H_1[13], inputSelect1H_0[13]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_13 = {inputSelect1H_3[13], inputSelect1H_2[13]};
  wire [3:0]  tryToRead_lo_lo_lo_13 = {tryToRead_lo_lo_lo_hi_13, tryToRead_lo_lo_lo_lo_13};
  wire [1:0]  tryToRead_lo_lo_hi_lo_13 = {inputSelect1H_5[13], inputSelect1H_4[13]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_13 = {inputSelect1H_7[13], inputSelect1H_6[13]};
  wire [3:0]  tryToRead_lo_lo_hi_13 = {tryToRead_lo_lo_hi_hi_13, tryToRead_lo_lo_hi_lo_13};
  wire [7:0]  tryToRead_lo_lo_13 = {tryToRead_lo_lo_hi_13, tryToRead_lo_lo_lo_13};
  wire [1:0]  tryToRead_lo_hi_lo_lo_13 = {inputSelect1H_9[13], inputSelect1H_8[13]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_13 = {inputSelect1H_11[13], inputSelect1H_10[13]};
  wire [3:0]  tryToRead_lo_hi_lo_13 = {tryToRead_lo_hi_lo_hi_13, tryToRead_lo_hi_lo_lo_13};
  wire [1:0]  tryToRead_lo_hi_hi_lo_13 = {inputSelect1H_13[13], inputSelect1H_12[13]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_13 = {inputSelect1H_15[13], inputSelect1H_14[13]};
  wire [3:0]  tryToRead_lo_hi_hi_13 = {tryToRead_lo_hi_hi_hi_13, tryToRead_lo_hi_hi_lo_13};
  wire [7:0]  tryToRead_lo_hi_13 = {tryToRead_lo_hi_hi_13, tryToRead_lo_hi_lo_13};
  wire [15:0] tryToRead_lo_13 = {tryToRead_lo_hi_13, tryToRead_lo_lo_13};
  wire [1:0]  tryToRead_hi_lo_lo_lo_13 = {inputSelect1H_17[13], inputSelect1H_16[13]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_13 = {inputSelect1H_19[13], inputSelect1H_18[13]};
  wire [3:0]  tryToRead_hi_lo_lo_13 = {tryToRead_hi_lo_lo_hi_13, tryToRead_hi_lo_lo_lo_13};
  wire [1:0]  tryToRead_hi_lo_hi_lo_13 = {inputSelect1H_21[13], inputSelect1H_20[13]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_13 = {inputSelect1H_23[13], inputSelect1H_22[13]};
  wire [3:0]  tryToRead_hi_lo_hi_13 = {tryToRead_hi_lo_hi_hi_13, tryToRead_hi_lo_hi_lo_13};
  wire [7:0]  tryToRead_hi_lo_13 = {tryToRead_hi_lo_hi_13, tryToRead_hi_lo_lo_13};
  wire [1:0]  tryToRead_hi_hi_lo_lo_13 = {inputSelect1H_25[13], inputSelect1H_24[13]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_13 = {inputSelect1H_27[13], inputSelect1H_26[13]};
  wire [3:0]  tryToRead_hi_hi_lo_13 = {tryToRead_hi_hi_lo_hi_13, tryToRead_hi_hi_lo_lo_13};
  wire [1:0]  tryToRead_hi_hi_hi_lo_13 = {inputSelect1H_29[13], inputSelect1H_28[13]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_13 = {inputSelect1H_31[13], inputSelect1H_30[13]};
  wire [3:0]  tryToRead_hi_hi_hi_13 = {tryToRead_hi_hi_hi_hi_13, tryToRead_hi_hi_hi_lo_13};
  wire [7:0]  tryToRead_hi_hi_13 = {tryToRead_hi_hi_hi_13, tryToRead_hi_hi_lo_13};
  wire [15:0] tryToRead_hi_13 = {tryToRead_hi_hi_13, tryToRead_hi_lo_13};
  wire [31:0] tryToRead_13 = {tryToRead_hi_13, tryToRead_lo_13};
  wire        output_13_valid_0 = |tryToRead_13;
  wire [4:0]  output_13_bits_vs_0 = selectReq_13_bits_vs;
  wire        output_13_bits_offset_0 = selectReq_13_bits_offset;
  wire [4:0]  output_13_bits_writeIndex_0 = selectReq_13_bits_requestIndex;
  wire [1:0]  output_13_bits_dataOffset_0 = selectReq_13_bits_dataOffset;
  assign selectReq_13_bits_dataOffset =
    (tryToRead_13[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_13[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_13[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_13[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_13[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_13[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_13[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_13[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_13[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_13[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_13[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_13[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_13[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_13[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_13[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_13[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_13[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_13[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_13[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_13[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_13[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_13[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_13[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_13[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_13[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_13_bits_requestIndex =
    {4'h0, tryToRead_13[1]} | {3'h0, tryToRead_13[2], 1'h0} | (tryToRead_13[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_13[4], 2'h0} | (tryToRead_13[5] ? 5'h5 : 5'h0) | (tryToRead_13[6] ? 5'h6 : 5'h0) | (tryToRead_13[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_13[8], 3'h0} | (tryToRead_13[9] ? 5'h9 : 5'h0) | (tryToRead_13[10] ? 5'hA : 5'h0) | (tryToRead_13[11] ? 5'hB : 5'h0) | (tryToRead_13[12] ? 5'hC : 5'h0) | (tryToRead_13[13] ? 5'hD : 5'h0)
    | (tryToRead_13[14] ? 5'hE : 5'h0) | (tryToRead_13[15] ? 5'hF : 5'h0) | {tryToRead_13[16], 4'h0} | (tryToRead_13[17] ? 5'h11 : 5'h0) | (tryToRead_13[18] ? 5'h12 : 5'h0) | (tryToRead_13[19] ? 5'h13 : 5'h0)
    | (tryToRead_13[20] ? 5'h14 : 5'h0) | (tryToRead_13[21] ? 5'h15 : 5'h0) | (tryToRead_13[22] ? 5'h16 : 5'h0) | (tryToRead_13[23] ? 5'h17 : 5'h0) | (tryToRead_13[24] ? 5'h18 : 5'h0) | (tryToRead_13[25] ? 5'h19 : 5'h0)
    | (tryToRead_13[26] ? 5'h1A : 5'h0) | (tryToRead_13[27] ? 5'h1B : 5'h0) | (tryToRead_13[28] ? 5'h1C : 5'h0) | (tryToRead_13[29] ? 5'h1D : 5'h0) | (tryToRead_13[30] ? 5'h1E : 5'h0) | {5{tryToRead_13[31]}};
  wire [4:0]  selectReq_13_bits_readLane =
    (tryToRead_13[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_13[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_13[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_13[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_13[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_13[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_13[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_13[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_13[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_13[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_13[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_13[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_13[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_13[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_13[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_13[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_13[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_13[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_13[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_13[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_13[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_13[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_13[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_13[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_13[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_13[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_13[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_13[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_13[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_13[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_13[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_13[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_13_bits_offset =
    tryToRead_13[0] & input_0_bits_offset_0 | tryToRead_13[1] & input_1_bits_offset_0 | tryToRead_13[2] & input_2_bits_offset_0 | tryToRead_13[3] & input_3_bits_offset_0 | tryToRead_13[4] & input_4_bits_offset_0 | tryToRead_13[5]
    & input_5_bits_offset_0 | tryToRead_13[6] & input_6_bits_offset_0 | tryToRead_13[7] & input_7_bits_offset_0 | tryToRead_13[8] & input_8_bits_offset_0 | tryToRead_13[9] & input_9_bits_offset_0 | tryToRead_13[10] & input_10_bits_offset_0
    | tryToRead_13[11] & input_11_bits_offset_0 | tryToRead_13[12] & input_12_bits_offset_0 | tryToRead_13[13] & input_13_bits_offset_0 | tryToRead_13[14] & input_14_bits_offset_0 | tryToRead_13[15] & input_15_bits_offset_0
    | tryToRead_13[16] & input_16_bits_offset_0 | tryToRead_13[17] & input_17_bits_offset_0 | tryToRead_13[18] & input_18_bits_offset_0 | tryToRead_13[19] & input_19_bits_offset_0 | tryToRead_13[20] & input_20_bits_offset_0
    | tryToRead_13[21] & input_21_bits_offset_0 | tryToRead_13[22] & input_22_bits_offset_0 | tryToRead_13[23] & input_23_bits_offset_0 | tryToRead_13[24] & input_24_bits_offset_0 | tryToRead_13[25] & input_25_bits_offset_0
    | tryToRead_13[26] & input_26_bits_offset_0 | tryToRead_13[27] & input_27_bits_offset_0 | tryToRead_13[28] & input_28_bits_offset_0 | tryToRead_13[29] & input_29_bits_offset_0 | tryToRead_13[30] & input_30_bits_offset_0
    | tryToRead_13[31] & input_31_bits_offset_0;
  assign selectReq_13_bits_vs =
    (tryToRead_13[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_13[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_13[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_13[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_13[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_13[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_13[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_13[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_13[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_13[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_13[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_13[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_13[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_13[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_13[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_13[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_13[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_13[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_13[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_13[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_13[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_13[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_13[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_13[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_13[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_13[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_13[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_13[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_13[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_13[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_13[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_13[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_13_valid =
    tryToRead_13[0] & input_0_valid_0 | tryToRead_13[1] & input_1_valid_0 | tryToRead_13[2] & input_2_valid_0 | tryToRead_13[3] & input_3_valid_0 | tryToRead_13[4] & input_4_valid_0 | tryToRead_13[5] & input_5_valid_0 | tryToRead_13[6]
    & input_6_valid_0 | tryToRead_13[7] & input_7_valid_0 | tryToRead_13[8] & input_8_valid_0 | tryToRead_13[9] & input_9_valid_0 | tryToRead_13[10] & input_10_valid_0 | tryToRead_13[11] & input_11_valid_0 | tryToRead_13[12]
    & input_12_valid_0 | tryToRead_13[13] & input_13_valid_0 | tryToRead_13[14] & input_14_valid_0 | tryToRead_13[15] & input_15_valid_0 | tryToRead_13[16] & input_16_valid_0 | tryToRead_13[17] & input_17_valid_0 | tryToRead_13[18]
    & input_18_valid_0 | tryToRead_13[19] & input_19_valid_0 | tryToRead_13[20] & input_20_valid_0 | tryToRead_13[21] & input_21_valid_0 | tryToRead_13[22] & input_22_valid_0 | tryToRead_13[23] & input_23_valid_0 | tryToRead_13[24]
    & input_24_valid_0 | tryToRead_13[25] & input_25_valid_0 | tryToRead_13[26] & input_26_valid_0 | tryToRead_13[27] & input_27_valid_0 | tryToRead_13[28] & input_28_valid_0 | tryToRead_13[29] & input_29_valid_0 | tryToRead_13[30]
    & input_30_valid_0 | tryToRead_13[31] & input_31_valid_0;
  wire        selectReq_13_ready =
    tryToRead_13[0] & input_0_ready_0 | tryToRead_13[1] & input_1_ready_0 | tryToRead_13[2] & input_2_ready_0 | tryToRead_13[3] & input_3_ready_0 | tryToRead_13[4] & input_4_ready_0 | tryToRead_13[5] & input_5_ready_0 | tryToRead_13[6]
    & input_6_ready_0 | tryToRead_13[7] & input_7_ready_0 | tryToRead_13[8] & input_8_ready_0 | tryToRead_13[9] & input_9_ready_0 | tryToRead_13[10] & input_10_ready_0 | tryToRead_13[11] & input_11_ready_0 | tryToRead_13[12]
    & input_12_ready_0 | tryToRead_13[13] & input_13_ready_0 | tryToRead_13[14] & input_14_ready_0 | tryToRead_13[15] & input_15_ready_0 | tryToRead_13[16] & input_16_ready_0 | tryToRead_13[17] & input_17_ready_0 | tryToRead_13[18]
    & input_18_ready_0 | tryToRead_13[19] & input_19_ready_0 | tryToRead_13[20] & input_20_ready_0 | tryToRead_13[21] & input_21_ready_0 | tryToRead_13[22] & input_22_ready_0 | tryToRead_13[23] & input_23_ready_0 | tryToRead_13[24]
    & input_24_ready_0 | tryToRead_13[25] & input_25_ready_0 | tryToRead_13[26] & input_26_ready_0 | tryToRead_13[27] & input_27_ready_0 | tryToRead_13[28] & input_28_ready_0 | tryToRead_13[29] & input_29_ready_0 | tryToRead_13[30]
    & input_30_ready_0 | tryToRead_13[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_14 = {inputSelect1H_1[14], inputSelect1H_0[14]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_14 = {inputSelect1H_3[14], inputSelect1H_2[14]};
  wire [3:0]  tryToRead_lo_lo_lo_14 = {tryToRead_lo_lo_lo_hi_14, tryToRead_lo_lo_lo_lo_14};
  wire [1:0]  tryToRead_lo_lo_hi_lo_14 = {inputSelect1H_5[14], inputSelect1H_4[14]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_14 = {inputSelect1H_7[14], inputSelect1H_6[14]};
  wire [3:0]  tryToRead_lo_lo_hi_14 = {tryToRead_lo_lo_hi_hi_14, tryToRead_lo_lo_hi_lo_14};
  wire [7:0]  tryToRead_lo_lo_14 = {tryToRead_lo_lo_hi_14, tryToRead_lo_lo_lo_14};
  wire [1:0]  tryToRead_lo_hi_lo_lo_14 = {inputSelect1H_9[14], inputSelect1H_8[14]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_14 = {inputSelect1H_11[14], inputSelect1H_10[14]};
  wire [3:0]  tryToRead_lo_hi_lo_14 = {tryToRead_lo_hi_lo_hi_14, tryToRead_lo_hi_lo_lo_14};
  wire [1:0]  tryToRead_lo_hi_hi_lo_14 = {inputSelect1H_13[14], inputSelect1H_12[14]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_14 = {inputSelect1H_15[14], inputSelect1H_14[14]};
  wire [3:0]  tryToRead_lo_hi_hi_14 = {tryToRead_lo_hi_hi_hi_14, tryToRead_lo_hi_hi_lo_14};
  wire [7:0]  tryToRead_lo_hi_14 = {tryToRead_lo_hi_hi_14, tryToRead_lo_hi_lo_14};
  wire [15:0] tryToRead_lo_14 = {tryToRead_lo_hi_14, tryToRead_lo_lo_14};
  wire [1:0]  tryToRead_hi_lo_lo_lo_14 = {inputSelect1H_17[14], inputSelect1H_16[14]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_14 = {inputSelect1H_19[14], inputSelect1H_18[14]};
  wire [3:0]  tryToRead_hi_lo_lo_14 = {tryToRead_hi_lo_lo_hi_14, tryToRead_hi_lo_lo_lo_14};
  wire [1:0]  tryToRead_hi_lo_hi_lo_14 = {inputSelect1H_21[14], inputSelect1H_20[14]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_14 = {inputSelect1H_23[14], inputSelect1H_22[14]};
  wire [3:0]  tryToRead_hi_lo_hi_14 = {tryToRead_hi_lo_hi_hi_14, tryToRead_hi_lo_hi_lo_14};
  wire [7:0]  tryToRead_hi_lo_14 = {tryToRead_hi_lo_hi_14, tryToRead_hi_lo_lo_14};
  wire [1:0]  tryToRead_hi_hi_lo_lo_14 = {inputSelect1H_25[14], inputSelect1H_24[14]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_14 = {inputSelect1H_27[14], inputSelect1H_26[14]};
  wire [3:0]  tryToRead_hi_hi_lo_14 = {tryToRead_hi_hi_lo_hi_14, tryToRead_hi_hi_lo_lo_14};
  wire [1:0]  tryToRead_hi_hi_hi_lo_14 = {inputSelect1H_29[14], inputSelect1H_28[14]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_14 = {inputSelect1H_31[14], inputSelect1H_30[14]};
  wire [3:0]  tryToRead_hi_hi_hi_14 = {tryToRead_hi_hi_hi_hi_14, tryToRead_hi_hi_hi_lo_14};
  wire [7:0]  tryToRead_hi_hi_14 = {tryToRead_hi_hi_hi_14, tryToRead_hi_hi_lo_14};
  wire [15:0] tryToRead_hi_14 = {tryToRead_hi_hi_14, tryToRead_hi_lo_14};
  wire [31:0] tryToRead_14 = {tryToRead_hi_14, tryToRead_lo_14};
  wire        output_14_valid_0 = |tryToRead_14;
  wire [4:0]  output_14_bits_vs_0 = selectReq_14_bits_vs;
  wire        output_14_bits_offset_0 = selectReq_14_bits_offset;
  wire [4:0]  output_14_bits_writeIndex_0 = selectReq_14_bits_requestIndex;
  wire [1:0]  output_14_bits_dataOffset_0 = selectReq_14_bits_dataOffset;
  assign selectReq_14_bits_dataOffset =
    (tryToRead_14[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_14[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_14[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_14[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_14[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_14[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_14[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_14[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_14[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_14[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_14[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_14[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_14[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_14[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_14[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_14[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_14[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_14[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_14[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_14[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_14[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_14[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_14[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_14[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_14[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_14_bits_requestIndex =
    {4'h0, tryToRead_14[1]} | {3'h0, tryToRead_14[2], 1'h0} | (tryToRead_14[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_14[4], 2'h0} | (tryToRead_14[5] ? 5'h5 : 5'h0) | (tryToRead_14[6] ? 5'h6 : 5'h0) | (tryToRead_14[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_14[8], 3'h0} | (tryToRead_14[9] ? 5'h9 : 5'h0) | (tryToRead_14[10] ? 5'hA : 5'h0) | (tryToRead_14[11] ? 5'hB : 5'h0) | (tryToRead_14[12] ? 5'hC : 5'h0) | (tryToRead_14[13] ? 5'hD : 5'h0)
    | (tryToRead_14[14] ? 5'hE : 5'h0) | (tryToRead_14[15] ? 5'hF : 5'h0) | {tryToRead_14[16], 4'h0} | (tryToRead_14[17] ? 5'h11 : 5'h0) | (tryToRead_14[18] ? 5'h12 : 5'h0) | (tryToRead_14[19] ? 5'h13 : 5'h0)
    | (tryToRead_14[20] ? 5'h14 : 5'h0) | (tryToRead_14[21] ? 5'h15 : 5'h0) | (tryToRead_14[22] ? 5'h16 : 5'h0) | (tryToRead_14[23] ? 5'h17 : 5'h0) | (tryToRead_14[24] ? 5'h18 : 5'h0) | (tryToRead_14[25] ? 5'h19 : 5'h0)
    | (tryToRead_14[26] ? 5'h1A : 5'h0) | (tryToRead_14[27] ? 5'h1B : 5'h0) | (tryToRead_14[28] ? 5'h1C : 5'h0) | (tryToRead_14[29] ? 5'h1D : 5'h0) | (tryToRead_14[30] ? 5'h1E : 5'h0) | {5{tryToRead_14[31]}};
  wire [4:0]  selectReq_14_bits_readLane =
    (tryToRead_14[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_14[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_14[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_14[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_14[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_14[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_14[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_14[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_14[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_14[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_14[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_14[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_14[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_14[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_14[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_14[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_14[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_14[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_14[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_14[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_14[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_14[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_14[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_14[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_14[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_14[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_14[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_14[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_14[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_14[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_14[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_14[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_14_bits_offset =
    tryToRead_14[0] & input_0_bits_offset_0 | tryToRead_14[1] & input_1_bits_offset_0 | tryToRead_14[2] & input_2_bits_offset_0 | tryToRead_14[3] & input_3_bits_offset_0 | tryToRead_14[4] & input_4_bits_offset_0 | tryToRead_14[5]
    & input_5_bits_offset_0 | tryToRead_14[6] & input_6_bits_offset_0 | tryToRead_14[7] & input_7_bits_offset_0 | tryToRead_14[8] & input_8_bits_offset_0 | tryToRead_14[9] & input_9_bits_offset_0 | tryToRead_14[10] & input_10_bits_offset_0
    | tryToRead_14[11] & input_11_bits_offset_0 | tryToRead_14[12] & input_12_bits_offset_0 | tryToRead_14[13] & input_13_bits_offset_0 | tryToRead_14[14] & input_14_bits_offset_0 | tryToRead_14[15] & input_15_bits_offset_0
    | tryToRead_14[16] & input_16_bits_offset_0 | tryToRead_14[17] & input_17_bits_offset_0 | tryToRead_14[18] & input_18_bits_offset_0 | tryToRead_14[19] & input_19_bits_offset_0 | tryToRead_14[20] & input_20_bits_offset_0
    | tryToRead_14[21] & input_21_bits_offset_0 | tryToRead_14[22] & input_22_bits_offset_0 | tryToRead_14[23] & input_23_bits_offset_0 | tryToRead_14[24] & input_24_bits_offset_0 | tryToRead_14[25] & input_25_bits_offset_0
    | tryToRead_14[26] & input_26_bits_offset_0 | tryToRead_14[27] & input_27_bits_offset_0 | tryToRead_14[28] & input_28_bits_offset_0 | tryToRead_14[29] & input_29_bits_offset_0 | tryToRead_14[30] & input_30_bits_offset_0
    | tryToRead_14[31] & input_31_bits_offset_0;
  assign selectReq_14_bits_vs =
    (tryToRead_14[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_14[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_14[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_14[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_14[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_14[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_14[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_14[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_14[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_14[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_14[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_14[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_14[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_14[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_14[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_14[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_14[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_14[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_14[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_14[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_14[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_14[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_14[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_14[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_14[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_14[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_14[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_14[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_14[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_14[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_14[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_14[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_14_valid =
    tryToRead_14[0] & input_0_valid_0 | tryToRead_14[1] & input_1_valid_0 | tryToRead_14[2] & input_2_valid_0 | tryToRead_14[3] & input_3_valid_0 | tryToRead_14[4] & input_4_valid_0 | tryToRead_14[5] & input_5_valid_0 | tryToRead_14[6]
    & input_6_valid_0 | tryToRead_14[7] & input_7_valid_0 | tryToRead_14[8] & input_8_valid_0 | tryToRead_14[9] & input_9_valid_0 | tryToRead_14[10] & input_10_valid_0 | tryToRead_14[11] & input_11_valid_0 | tryToRead_14[12]
    & input_12_valid_0 | tryToRead_14[13] & input_13_valid_0 | tryToRead_14[14] & input_14_valid_0 | tryToRead_14[15] & input_15_valid_0 | tryToRead_14[16] & input_16_valid_0 | tryToRead_14[17] & input_17_valid_0 | tryToRead_14[18]
    & input_18_valid_0 | tryToRead_14[19] & input_19_valid_0 | tryToRead_14[20] & input_20_valid_0 | tryToRead_14[21] & input_21_valid_0 | tryToRead_14[22] & input_22_valid_0 | tryToRead_14[23] & input_23_valid_0 | tryToRead_14[24]
    & input_24_valid_0 | tryToRead_14[25] & input_25_valid_0 | tryToRead_14[26] & input_26_valid_0 | tryToRead_14[27] & input_27_valid_0 | tryToRead_14[28] & input_28_valid_0 | tryToRead_14[29] & input_29_valid_0 | tryToRead_14[30]
    & input_30_valid_0 | tryToRead_14[31] & input_31_valid_0;
  wire        selectReq_14_ready =
    tryToRead_14[0] & input_0_ready_0 | tryToRead_14[1] & input_1_ready_0 | tryToRead_14[2] & input_2_ready_0 | tryToRead_14[3] & input_3_ready_0 | tryToRead_14[4] & input_4_ready_0 | tryToRead_14[5] & input_5_ready_0 | tryToRead_14[6]
    & input_6_ready_0 | tryToRead_14[7] & input_7_ready_0 | tryToRead_14[8] & input_8_ready_0 | tryToRead_14[9] & input_9_ready_0 | tryToRead_14[10] & input_10_ready_0 | tryToRead_14[11] & input_11_ready_0 | tryToRead_14[12]
    & input_12_ready_0 | tryToRead_14[13] & input_13_ready_0 | tryToRead_14[14] & input_14_ready_0 | tryToRead_14[15] & input_15_ready_0 | tryToRead_14[16] & input_16_ready_0 | tryToRead_14[17] & input_17_ready_0 | tryToRead_14[18]
    & input_18_ready_0 | tryToRead_14[19] & input_19_ready_0 | tryToRead_14[20] & input_20_ready_0 | tryToRead_14[21] & input_21_ready_0 | tryToRead_14[22] & input_22_ready_0 | tryToRead_14[23] & input_23_ready_0 | tryToRead_14[24]
    & input_24_ready_0 | tryToRead_14[25] & input_25_ready_0 | tryToRead_14[26] & input_26_ready_0 | tryToRead_14[27] & input_27_ready_0 | tryToRead_14[28] & input_28_ready_0 | tryToRead_14[29] & input_29_ready_0 | tryToRead_14[30]
    & input_30_ready_0 | tryToRead_14[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_15 = {inputSelect1H_1[15], inputSelect1H_0[15]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_15 = {inputSelect1H_3[15], inputSelect1H_2[15]};
  wire [3:0]  tryToRead_lo_lo_lo_15 = {tryToRead_lo_lo_lo_hi_15, tryToRead_lo_lo_lo_lo_15};
  wire [1:0]  tryToRead_lo_lo_hi_lo_15 = {inputSelect1H_5[15], inputSelect1H_4[15]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_15 = {inputSelect1H_7[15], inputSelect1H_6[15]};
  wire [3:0]  tryToRead_lo_lo_hi_15 = {tryToRead_lo_lo_hi_hi_15, tryToRead_lo_lo_hi_lo_15};
  wire [7:0]  tryToRead_lo_lo_15 = {tryToRead_lo_lo_hi_15, tryToRead_lo_lo_lo_15};
  wire [1:0]  tryToRead_lo_hi_lo_lo_15 = {inputSelect1H_9[15], inputSelect1H_8[15]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_15 = {inputSelect1H_11[15], inputSelect1H_10[15]};
  wire [3:0]  tryToRead_lo_hi_lo_15 = {tryToRead_lo_hi_lo_hi_15, tryToRead_lo_hi_lo_lo_15};
  wire [1:0]  tryToRead_lo_hi_hi_lo_15 = {inputSelect1H_13[15], inputSelect1H_12[15]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_15 = {inputSelect1H_15[15], inputSelect1H_14[15]};
  wire [3:0]  tryToRead_lo_hi_hi_15 = {tryToRead_lo_hi_hi_hi_15, tryToRead_lo_hi_hi_lo_15};
  wire [7:0]  tryToRead_lo_hi_15 = {tryToRead_lo_hi_hi_15, tryToRead_lo_hi_lo_15};
  wire [15:0] tryToRead_lo_15 = {tryToRead_lo_hi_15, tryToRead_lo_lo_15};
  wire [1:0]  tryToRead_hi_lo_lo_lo_15 = {inputSelect1H_17[15], inputSelect1H_16[15]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_15 = {inputSelect1H_19[15], inputSelect1H_18[15]};
  wire [3:0]  tryToRead_hi_lo_lo_15 = {tryToRead_hi_lo_lo_hi_15, tryToRead_hi_lo_lo_lo_15};
  wire [1:0]  tryToRead_hi_lo_hi_lo_15 = {inputSelect1H_21[15], inputSelect1H_20[15]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_15 = {inputSelect1H_23[15], inputSelect1H_22[15]};
  wire [3:0]  tryToRead_hi_lo_hi_15 = {tryToRead_hi_lo_hi_hi_15, tryToRead_hi_lo_hi_lo_15};
  wire [7:0]  tryToRead_hi_lo_15 = {tryToRead_hi_lo_hi_15, tryToRead_hi_lo_lo_15};
  wire [1:0]  tryToRead_hi_hi_lo_lo_15 = {inputSelect1H_25[15], inputSelect1H_24[15]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_15 = {inputSelect1H_27[15], inputSelect1H_26[15]};
  wire [3:0]  tryToRead_hi_hi_lo_15 = {tryToRead_hi_hi_lo_hi_15, tryToRead_hi_hi_lo_lo_15};
  wire [1:0]  tryToRead_hi_hi_hi_lo_15 = {inputSelect1H_29[15], inputSelect1H_28[15]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_15 = {inputSelect1H_31[15], inputSelect1H_30[15]};
  wire [3:0]  tryToRead_hi_hi_hi_15 = {tryToRead_hi_hi_hi_hi_15, tryToRead_hi_hi_hi_lo_15};
  wire [7:0]  tryToRead_hi_hi_15 = {tryToRead_hi_hi_hi_15, tryToRead_hi_hi_lo_15};
  wire [15:0] tryToRead_hi_15 = {tryToRead_hi_hi_15, tryToRead_hi_lo_15};
  wire [31:0] tryToRead_15 = {tryToRead_hi_15, tryToRead_lo_15};
  wire        output_15_valid_0 = |tryToRead_15;
  wire [4:0]  output_15_bits_vs_0 = selectReq_15_bits_vs;
  wire        output_15_bits_offset_0 = selectReq_15_bits_offset;
  wire [4:0]  output_15_bits_writeIndex_0 = selectReq_15_bits_requestIndex;
  wire [1:0]  output_15_bits_dataOffset_0 = selectReq_15_bits_dataOffset;
  assign selectReq_15_bits_dataOffset =
    (tryToRead_15[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_15[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_15[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_15[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_15[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_15[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_15[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_15[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_15[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_15[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_15[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_15[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_15[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_15[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_15[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_15[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_15[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_15[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_15[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_15[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_15[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_15[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_15[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_15[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_15[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_15_bits_requestIndex =
    {4'h0, tryToRead_15[1]} | {3'h0, tryToRead_15[2], 1'h0} | (tryToRead_15[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_15[4], 2'h0} | (tryToRead_15[5] ? 5'h5 : 5'h0) | (tryToRead_15[6] ? 5'h6 : 5'h0) | (tryToRead_15[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_15[8], 3'h0} | (tryToRead_15[9] ? 5'h9 : 5'h0) | (tryToRead_15[10] ? 5'hA : 5'h0) | (tryToRead_15[11] ? 5'hB : 5'h0) | (tryToRead_15[12] ? 5'hC : 5'h0) | (tryToRead_15[13] ? 5'hD : 5'h0)
    | (tryToRead_15[14] ? 5'hE : 5'h0) | (tryToRead_15[15] ? 5'hF : 5'h0) | {tryToRead_15[16], 4'h0} | (tryToRead_15[17] ? 5'h11 : 5'h0) | (tryToRead_15[18] ? 5'h12 : 5'h0) | (tryToRead_15[19] ? 5'h13 : 5'h0)
    | (tryToRead_15[20] ? 5'h14 : 5'h0) | (tryToRead_15[21] ? 5'h15 : 5'h0) | (tryToRead_15[22] ? 5'h16 : 5'h0) | (tryToRead_15[23] ? 5'h17 : 5'h0) | (tryToRead_15[24] ? 5'h18 : 5'h0) | (tryToRead_15[25] ? 5'h19 : 5'h0)
    | (tryToRead_15[26] ? 5'h1A : 5'h0) | (tryToRead_15[27] ? 5'h1B : 5'h0) | (tryToRead_15[28] ? 5'h1C : 5'h0) | (tryToRead_15[29] ? 5'h1D : 5'h0) | (tryToRead_15[30] ? 5'h1E : 5'h0) | {5{tryToRead_15[31]}};
  wire [4:0]  selectReq_15_bits_readLane =
    (tryToRead_15[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_15[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_15[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_15[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_15[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_15[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_15[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_15[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_15[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_15[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_15[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_15[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_15[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_15[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_15[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_15[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_15[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_15[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_15[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_15[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_15[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_15[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_15[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_15[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_15[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_15[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_15[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_15[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_15[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_15[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_15[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_15[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_15_bits_offset =
    tryToRead_15[0] & input_0_bits_offset_0 | tryToRead_15[1] & input_1_bits_offset_0 | tryToRead_15[2] & input_2_bits_offset_0 | tryToRead_15[3] & input_3_bits_offset_0 | tryToRead_15[4] & input_4_bits_offset_0 | tryToRead_15[5]
    & input_5_bits_offset_0 | tryToRead_15[6] & input_6_bits_offset_0 | tryToRead_15[7] & input_7_bits_offset_0 | tryToRead_15[8] & input_8_bits_offset_0 | tryToRead_15[9] & input_9_bits_offset_0 | tryToRead_15[10] & input_10_bits_offset_0
    | tryToRead_15[11] & input_11_bits_offset_0 | tryToRead_15[12] & input_12_bits_offset_0 | tryToRead_15[13] & input_13_bits_offset_0 | tryToRead_15[14] & input_14_bits_offset_0 | tryToRead_15[15] & input_15_bits_offset_0
    | tryToRead_15[16] & input_16_bits_offset_0 | tryToRead_15[17] & input_17_bits_offset_0 | tryToRead_15[18] & input_18_bits_offset_0 | tryToRead_15[19] & input_19_bits_offset_0 | tryToRead_15[20] & input_20_bits_offset_0
    | tryToRead_15[21] & input_21_bits_offset_0 | tryToRead_15[22] & input_22_bits_offset_0 | tryToRead_15[23] & input_23_bits_offset_0 | tryToRead_15[24] & input_24_bits_offset_0 | tryToRead_15[25] & input_25_bits_offset_0
    | tryToRead_15[26] & input_26_bits_offset_0 | tryToRead_15[27] & input_27_bits_offset_0 | tryToRead_15[28] & input_28_bits_offset_0 | tryToRead_15[29] & input_29_bits_offset_0 | tryToRead_15[30] & input_30_bits_offset_0
    | tryToRead_15[31] & input_31_bits_offset_0;
  assign selectReq_15_bits_vs =
    (tryToRead_15[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_15[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_15[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_15[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_15[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_15[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_15[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_15[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_15[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_15[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_15[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_15[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_15[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_15[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_15[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_15[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_15[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_15[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_15[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_15[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_15[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_15[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_15[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_15[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_15[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_15[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_15[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_15[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_15[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_15[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_15[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_15[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_15_valid =
    tryToRead_15[0] & input_0_valid_0 | tryToRead_15[1] & input_1_valid_0 | tryToRead_15[2] & input_2_valid_0 | tryToRead_15[3] & input_3_valid_0 | tryToRead_15[4] & input_4_valid_0 | tryToRead_15[5] & input_5_valid_0 | tryToRead_15[6]
    & input_6_valid_0 | tryToRead_15[7] & input_7_valid_0 | tryToRead_15[8] & input_8_valid_0 | tryToRead_15[9] & input_9_valid_0 | tryToRead_15[10] & input_10_valid_0 | tryToRead_15[11] & input_11_valid_0 | tryToRead_15[12]
    & input_12_valid_0 | tryToRead_15[13] & input_13_valid_0 | tryToRead_15[14] & input_14_valid_0 | tryToRead_15[15] & input_15_valid_0 | tryToRead_15[16] & input_16_valid_0 | tryToRead_15[17] & input_17_valid_0 | tryToRead_15[18]
    & input_18_valid_0 | tryToRead_15[19] & input_19_valid_0 | tryToRead_15[20] & input_20_valid_0 | tryToRead_15[21] & input_21_valid_0 | tryToRead_15[22] & input_22_valid_0 | tryToRead_15[23] & input_23_valid_0 | tryToRead_15[24]
    & input_24_valid_0 | tryToRead_15[25] & input_25_valid_0 | tryToRead_15[26] & input_26_valid_0 | tryToRead_15[27] & input_27_valid_0 | tryToRead_15[28] & input_28_valid_0 | tryToRead_15[29] & input_29_valid_0 | tryToRead_15[30]
    & input_30_valid_0 | tryToRead_15[31] & input_31_valid_0;
  wire        selectReq_15_ready =
    tryToRead_15[0] & input_0_ready_0 | tryToRead_15[1] & input_1_ready_0 | tryToRead_15[2] & input_2_ready_0 | tryToRead_15[3] & input_3_ready_0 | tryToRead_15[4] & input_4_ready_0 | tryToRead_15[5] & input_5_ready_0 | tryToRead_15[6]
    & input_6_ready_0 | tryToRead_15[7] & input_7_ready_0 | tryToRead_15[8] & input_8_ready_0 | tryToRead_15[9] & input_9_ready_0 | tryToRead_15[10] & input_10_ready_0 | tryToRead_15[11] & input_11_ready_0 | tryToRead_15[12]
    & input_12_ready_0 | tryToRead_15[13] & input_13_ready_0 | tryToRead_15[14] & input_14_ready_0 | tryToRead_15[15] & input_15_ready_0 | tryToRead_15[16] & input_16_ready_0 | tryToRead_15[17] & input_17_ready_0 | tryToRead_15[18]
    & input_18_ready_0 | tryToRead_15[19] & input_19_ready_0 | tryToRead_15[20] & input_20_ready_0 | tryToRead_15[21] & input_21_ready_0 | tryToRead_15[22] & input_22_ready_0 | tryToRead_15[23] & input_23_ready_0 | tryToRead_15[24]
    & input_24_ready_0 | tryToRead_15[25] & input_25_ready_0 | tryToRead_15[26] & input_26_ready_0 | tryToRead_15[27] & input_27_ready_0 | tryToRead_15[28] & input_28_ready_0 | tryToRead_15[29] & input_29_ready_0 | tryToRead_15[30]
    & input_30_ready_0 | tryToRead_15[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_16 = {inputSelect1H_1[16], inputSelect1H_0[16]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_16 = {inputSelect1H_3[16], inputSelect1H_2[16]};
  wire [3:0]  tryToRead_lo_lo_lo_16 = {tryToRead_lo_lo_lo_hi_16, tryToRead_lo_lo_lo_lo_16};
  wire [1:0]  tryToRead_lo_lo_hi_lo_16 = {inputSelect1H_5[16], inputSelect1H_4[16]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_16 = {inputSelect1H_7[16], inputSelect1H_6[16]};
  wire [3:0]  tryToRead_lo_lo_hi_16 = {tryToRead_lo_lo_hi_hi_16, tryToRead_lo_lo_hi_lo_16};
  wire [7:0]  tryToRead_lo_lo_16 = {tryToRead_lo_lo_hi_16, tryToRead_lo_lo_lo_16};
  wire [1:0]  tryToRead_lo_hi_lo_lo_16 = {inputSelect1H_9[16], inputSelect1H_8[16]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_16 = {inputSelect1H_11[16], inputSelect1H_10[16]};
  wire [3:0]  tryToRead_lo_hi_lo_16 = {tryToRead_lo_hi_lo_hi_16, tryToRead_lo_hi_lo_lo_16};
  wire [1:0]  tryToRead_lo_hi_hi_lo_16 = {inputSelect1H_13[16], inputSelect1H_12[16]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_16 = {inputSelect1H_15[16], inputSelect1H_14[16]};
  wire [3:0]  tryToRead_lo_hi_hi_16 = {tryToRead_lo_hi_hi_hi_16, tryToRead_lo_hi_hi_lo_16};
  wire [7:0]  tryToRead_lo_hi_16 = {tryToRead_lo_hi_hi_16, tryToRead_lo_hi_lo_16};
  wire [15:0] tryToRead_lo_16 = {tryToRead_lo_hi_16, tryToRead_lo_lo_16};
  wire [1:0]  tryToRead_hi_lo_lo_lo_16 = {inputSelect1H_17[16], inputSelect1H_16[16]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_16 = {inputSelect1H_19[16], inputSelect1H_18[16]};
  wire [3:0]  tryToRead_hi_lo_lo_16 = {tryToRead_hi_lo_lo_hi_16, tryToRead_hi_lo_lo_lo_16};
  wire [1:0]  tryToRead_hi_lo_hi_lo_16 = {inputSelect1H_21[16], inputSelect1H_20[16]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_16 = {inputSelect1H_23[16], inputSelect1H_22[16]};
  wire [3:0]  tryToRead_hi_lo_hi_16 = {tryToRead_hi_lo_hi_hi_16, tryToRead_hi_lo_hi_lo_16};
  wire [7:0]  tryToRead_hi_lo_16 = {tryToRead_hi_lo_hi_16, tryToRead_hi_lo_lo_16};
  wire [1:0]  tryToRead_hi_hi_lo_lo_16 = {inputSelect1H_25[16], inputSelect1H_24[16]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_16 = {inputSelect1H_27[16], inputSelect1H_26[16]};
  wire [3:0]  tryToRead_hi_hi_lo_16 = {tryToRead_hi_hi_lo_hi_16, tryToRead_hi_hi_lo_lo_16};
  wire [1:0]  tryToRead_hi_hi_hi_lo_16 = {inputSelect1H_29[16], inputSelect1H_28[16]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_16 = {inputSelect1H_31[16], inputSelect1H_30[16]};
  wire [3:0]  tryToRead_hi_hi_hi_16 = {tryToRead_hi_hi_hi_hi_16, tryToRead_hi_hi_hi_lo_16};
  wire [7:0]  tryToRead_hi_hi_16 = {tryToRead_hi_hi_hi_16, tryToRead_hi_hi_lo_16};
  wire [15:0] tryToRead_hi_16 = {tryToRead_hi_hi_16, tryToRead_hi_lo_16};
  wire [31:0] tryToRead_16 = {tryToRead_hi_16, tryToRead_lo_16};
  wire        output_16_valid_0 = |tryToRead_16;
  wire [4:0]  output_16_bits_vs_0 = selectReq_16_bits_vs;
  wire        output_16_bits_offset_0 = selectReq_16_bits_offset;
  wire [4:0]  output_16_bits_writeIndex_0 = selectReq_16_bits_requestIndex;
  wire [1:0]  output_16_bits_dataOffset_0 = selectReq_16_bits_dataOffset;
  assign selectReq_16_bits_dataOffset =
    (tryToRead_16[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_16[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_16[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_16[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_16[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_16[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_16[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_16[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_16[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_16[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_16[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_16[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_16[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_16[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_16[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_16[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_16[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_16[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_16[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_16[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_16[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_16[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_16[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_16[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_16[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_16[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_16_bits_requestIndex =
    {4'h0, tryToRead_16[1]} | {3'h0, tryToRead_16[2], 1'h0} | (tryToRead_16[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_16[4], 2'h0} | (tryToRead_16[5] ? 5'h5 : 5'h0) | (tryToRead_16[6] ? 5'h6 : 5'h0) | (tryToRead_16[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_16[8], 3'h0} | (tryToRead_16[9] ? 5'h9 : 5'h0) | (tryToRead_16[10] ? 5'hA : 5'h0) | (tryToRead_16[11] ? 5'hB : 5'h0) | (tryToRead_16[12] ? 5'hC : 5'h0) | (tryToRead_16[13] ? 5'hD : 5'h0)
    | (tryToRead_16[14] ? 5'hE : 5'h0) | (tryToRead_16[15] ? 5'hF : 5'h0) | {tryToRead_16[16], 4'h0} | (tryToRead_16[17] ? 5'h11 : 5'h0) | (tryToRead_16[18] ? 5'h12 : 5'h0) | (tryToRead_16[19] ? 5'h13 : 5'h0)
    | (tryToRead_16[20] ? 5'h14 : 5'h0) | (tryToRead_16[21] ? 5'h15 : 5'h0) | (tryToRead_16[22] ? 5'h16 : 5'h0) | (tryToRead_16[23] ? 5'h17 : 5'h0) | (tryToRead_16[24] ? 5'h18 : 5'h0) | (tryToRead_16[25] ? 5'h19 : 5'h0)
    | (tryToRead_16[26] ? 5'h1A : 5'h0) | (tryToRead_16[27] ? 5'h1B : 5'h0) | (tryToRead_16[28] ? 5'h1C : 5'h0) | (tryToRead_16[29] ? 5'h1D : 5'h0) | (tryToRead_16[30] ? 5'h1E : 5'h0) | {5{tryToRead_16[31]}};
  wire [4:0]  selectReq_16_bits_readLane =
    (tryToRead_16[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_16[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_16[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_16[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_16[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_16[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_16[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_16[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_16[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_16[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_16[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_16[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_16[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_16[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_16[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_16[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_16[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_16[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_16[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_16[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_16[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_16[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_16[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_16[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_16[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_16[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_16[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_16[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_16[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_16[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_16[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_16[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_16_bits_offset =
    tryToRead_16[0] & input_0_bits_offset_0 | tryToRead_16[1] & input_1_bits_offset_0 | tryToRead_16[2] & input_2_bits_offset_0 | tryToRead_16[3] & input_3_bits_offset_0 | tryToRead_16[4] & input_4_bits_offset_0 | tryToRead_16[5]
    & input_5_bits_offset_0 | tryToRead_16[6] & input_6_bits_offset_0 | tryToRead_16[7] & input_7_bits_offset_0 | tryToRead_16[8] & input_8_bits_offset_0 | tryToRead_16[9] & input_9_bits_offset_0 | tryToRead_16[10] & input_10_bits_offset_0
    | tryToRead_16[11] & input_11_bits_offset_0 | tryToRead_16[12] & input_12_bits_offset_0 | tryToRead_16[13] & input_13_bits_offset_0 | tryToRead_16[14] & input_14_bits_offset_0 | tryToRead_16[15] & input_15_bits_offset_0
    | tryToRead_16[16] & input_16_bits_offset_0 | tryToRead_16[17] & input_17_bits_offset_0 | tryToRead_16[18] & input_18_bits_offset_0 | tryToRead_16[19] & input_19_bits_offset_0 | tryToRead_16[20] & input_20_bits_offset_0
    | tryToRead_16[21] & input_21_bits_offset_0 | tryToRead_16[22] & input_22_bits_offset_0 | tryToRead_16[23] & input_23_bits_offset_0 | tryToRead_16[24] & input_24_bits_offset_0 | tryToRead_16[25] & input_25_bits_offset_0
    | tryToRead_16[26] & input_26_bits_offset_0 | tryToRead_16[27] & input_27_bits_offset_0 | tryToRead_16[28] & input_28_bits_offset_0 | tryToRead_16[29] & input_29_bits_offset_0 | tryToRead_16[30] & input_30_bits_offset_0
    | tryToRead_16[31] & input_31_bits_offset_0;
  assign selectReq_16_bits_vs =
    (tryToRead_16[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_16[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_16[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_16[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_16[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_16[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_16[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_16[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_16[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_16[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_16[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_16[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_16[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_16[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_16[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_16[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_16[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_16[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_16[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_16[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_16[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_16[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_16[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_16[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_16[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_16[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_16[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_16[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_16[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_16[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_16[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_16[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_16_valid =
    tryToRead_16[0] & input_0_valid_0 | tryToRead_16[1] & input_1_valid_0 | tryToRead_16[2] & input_2_valid_0 | tryToRead_16[3] & input_3_valid_0 | tryToRead_16[4] & input_4_valid_0 | tryToRead_16[5] & input_5_valid_0 | tryToRead_16[6]
    & input_6_valid_0 | tryToRead_16[7] & input_7_valid_0 | tryToRead_16[8] & input_8_valid_0 | tryToRead_16[9] & input_9_valid_0 | tryToRead_16[10] & input_10_valid_0 | tryToRead_16[11] & input_11_valid_0 | tryToRead_16[12]
    & input_12_valid_0 | tryToRead_16[13] & input_13_valid_0 | tryToRead_16[14] & input_14_valid_0 | tryToRead_16[15] & input_15_valid_0 | tryToRead_16[16] & input_16_valid_0 | tryToRead_16[17] & input_17_valid_0 | tryToRead_16[18]
    & input_18_valid_0 | tryToRead_16[19] & input_19_valid_0 | tryToRead_16[20] & input_20_valid_0 | tryToRead_16[21] & input_21_valid_0 | tryToRead_16[22] & input_22_valid_0 | tryToRead_16[23] & input_23_valid_0 | tryToRead_16[24]
    & input_24_valid_0 | tryToRead_16[25] & input_25_valid_0 | tryToRead_16[26] & input_26_valid_0 | tryToRead_16[27] & input_27_valid_0 | tryToRead_16[28] & input_28_valid_0 | tryToRead_16[29] & input_29_valid_0 | tryToRead_16[30]
    & input_30_valid_0 | tryToRead_16[31] & input_31_valid_0;
  wire        selectReq_16_ready =
    tryToRead_16[0] & input_0_ready_0 | tryToRead_16[1] & input_1_ready_0 | tryToRead_16[2] & input_2_ready_0 | tryToRead_16[3] & input_3_ready_0 | tryToRead_16[4] & input_4_ready_0 | tryToRead_16[5] & input_5_ready_0 | tryToRead_16[6]
    & input_6_ready_0 | tryToRead_16[7] & input_7_ready_0 | tryToRead_16[8] & input_8_ready_0 | tryToRead_16[9] & input_9_ready_0 | tryToRead_16[10] & input_10_ready_0 | tryToRead_16[11] & input_11_ready_0 | tryToRead_16[12]
    & input_12_ready_0 | tryToRead_16[13] & input_13_ready_0 | tryToRead_16[14] & input_14_ready_0 | tryToRead_16[15] & input_15_ready_0 | tryToRead_16[16] & input_16_ready_0 | tryToRead_16[17] & input_17_ready_0 | tryToRead_16[18]
    & input_18_ready_0 | tryToRead_16[19] & input_19_ready_0 | tryToRead_16[20] & input_20_ready_0 | tryToRead_16[21] & input_21_ready_0 | tryToRead_16[22] & input_22_ready_0 | tryToRead_16[23] & input_23_ready_0 | tryToRead_16[24]
    & input_24_ready_0 | tryToRead_16[25] & input_25_ready_0 | tryToRead_16[26] & input_26_ready_0 | tryToRead_16[27] & input_27_ready_0 | tryToRead_16[28] & input_28_ready_0 | tryToRead_16[29] & input_29_ready_0 | tryToRead_16[30]
    & input_30_ready_0 | tryToRead_16[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_17 = {inputSelect1H_1[17], inputSelect1H_0[17]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_17 = {inputSelect1H_3[17], inputSelect1H_2[17]};
  wire [3:0]  tryToRead_lo_lo_lo_17 = {tryToRead_lo_lo_lo_hi_17, tryToRead_lo_lo_lo_lo_17};
  wire [1:0]  tryToRead_lo_lo_hi_lo_17 = {inputSelect1H_5[17], inputSelect1H_4[17]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_17 = {inputSelect1H_7[17], inputSelect1H_6[17]};
  wire [3:0]  tryToRead_lo_lo_hi_17 = {tryToRead_lo_lo_hi_hi_17, tryToRead_lo_lo_hi_lo_17};
  wire [7:0]  tryToRead_lo_lo_17 = {tryToRead_lo_lo_hi_17, tryToRead_lo_lo_lo_17};
  wire [1:0]  tryToRead_lo_hi_lo_lo_17 = {inputSelect1H_9[17], inputSelect1H_8[17]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_17 = {inputSelect1H_11[17], inputSelect1H_10[17]};
  wire [3:0]  tryToRead_lo_hi_lo_17 = {tryToRead_lo_hi_lo_hi_17, tryToRead_lo_hi_lo_lo_17};
  wire [1:0]  tryToRead_lo_hi_hi_lo_17 = {inputSelect1H_13[17], inputSelect1H_12[17]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_17 = {inputSelect1H_15[17], inputSelect1H_14[17]};
  wire [3:0]  tryToRead_lo_hi_hi_17 = {tryToRead_lo_hi_hi_hi_17, tryToRead_lo_hi_hi_lo_17};
  wire [7:0]  tryToRead_lo_hi_17 = {tryToRead_lo_hi_hi_17, tryToRead_lo_hi_lo_17};
  wire [15:0] tryToRead_lo_17 = {tryToRead_lo_hi_17, tryToRead_lo_lo_17};
  wire [1:0]  tryToRead_hi_lo_lo_lo_17 = {inputSelect1H_17[17], inputSelect1H_16[17]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_17 = {inputSelect1H_19[17], inputSelect1H_18[17]};
  wire [3:0]  tryToRead_hi_lo_lo_17 = {tryToRead_hi_lo_lo_hi_17, tryToRead_hi_lo_lo_lo_17};
  wire [1:0]  tryToRead_hi_lo_hi_lo_17 = {inputSelect1H_21[17], inputSelect1H_20[17]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_17 = {inputSelect1H_23[17], inputSelect1H_22[17]};
  wire [3:0]  tryToRead_hi_lo_hi_17 = {tryToRead_hi_lo_hi_hi_17, tryToRead_hi_lo_hi_lo_17};
  wire [7:0]  tryToRead_hi_lo_17 = {tryToRead_hi_lo_hi_17, tryToRead_hi_lo_lo_17};
  wire [1:0]  tryToRead_hi_hi_lo_lo_17 = {inputSelect1H_25[17], inputSelect1H_24[17]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_17 = {inputSelect1H_27[17], inputSelect1H_26[17]};
  wire [3:0]  tryToRead_hi_hi_lo_17 = {tryToRead_hi_hi_lo_hi_17, tryToRead_hi_hi_lo_lo_17};
  wire [1:0]  tryToRead_hi_hi_hi_lo_17 = {inputSelect1H_29[17], inputSelect1H_28[17]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_17 = {inputSelect1H_31[17], inputSelect1H_30[17]};
  wire [3:0]  tryToRead_hi_hi_hi_17 = {tryToRead_hi_hi_hi_hi_17, tryToRead_hi_hi_hi_lo_17};
  wire [7:0]  tryToRead_hi_hi_17 = {tryToRead_hi_hi_hi_17, tryToRead_hi_hi_lo_17};
  wire [15:0] tryToRead_hi_17 = {tryToRead_hi_hi_17, tryToRead_hi_lo_17};
  wire [31:0] tryToRead_17 = {tryToRead_hi_17, tryToRead_lo_17};
  wire        output_17_valid_0 = |tryToRead_17;
  wire [4:0]  output_17_bits_vs_0 = selectReq_17_bits_vs;
  wire        output_17_bits_offset_0 = selectReq_17_bits_offset;
  wire [4:0]  output_17_bits_writeIndex_0 = selectReq_17_bits_requestIndex;
  wire [1:0]  output_17_bits_dataOffset_0 = selectReq_17_bits_dataOffset;
  assign selectReq_17_bits_dataOffset =
    (tryToRead_17[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_17[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_17[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_17[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_17[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_17[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_17[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_17[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_17[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_17[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_17[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_17[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_17[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_17[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_17[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_17[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_17[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_17[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_17[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_17[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_17[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_17[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_17[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_17[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_17[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_17[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_17_bits_requestIndex =
    {4'h0, tryToRead_17[1]} | {3'h0, tryToRead_17[2], 1'h0} | (tryToRead_17[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_17[4], 2'h0} | (tryToRead_17[5] ? 5'h5 : 5'h0) | (tryToRead_17[6] ? 5'h6 : 5'h0) | (tryToRead_17[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_17[8], 3'h0} | (tryToRead_17[9] ? 5'h9 : 5'h0) | (tryToRead_17[10] ? 5'hA : 5'h0) | (tryToRead_17[11] ? 5'hB : 5'h0) | (tryToRead_17[12] ? 5'hC : 5'h0) | (tryToRead_17[13] ? 5'hD : 5'h0)
    | (tryToRead_17[14] ? 5'hE : 5'h0) | (tryToRead_17[15] ? 5'hF : 5'h0) | {tryToRead_17[16], 4'h0} | (tryToRead_17[17] ? 5'h11 : 5'h0) | (tryToRead_17[18] ? 5'h12 : 5'h0) | (tryToRead_17[19] ? 5'h13 : 5'h0)
    | (tryToRead_17[20] ? 5'h14 : 5'h0) | (tryToRead_17[21] ? 5'h15 : 5'h0) | (tryToRead_17[22] ? 5'h16 : 5'h0) | (tryToRead_17[23] ? 5'h17 : 5'h0) | (tryToRead_17[24] ? 5'h18 : 5'h0) | (tryToRead_17[25] ? 5'h19 : 5'h0)
    | (tryToRead_17[26] ? 5'h1A : 5'h0) | (tryToRead_17[27] ? 5'h1B : 5'h0) | (tryToRead_17[28] ? 5'h1C : 5'h0) | (tryToRead_17[29] ? 5'h1D : 5'h0) | (tryToRead_17[30] ? 5'h1E : 5'h0) | {5{tryToRead_17[31]}};
  wire [4:0]  selectReq_17_bits_readLane =
    (tryToRead_17[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_17[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_17[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_17[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_17[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_17[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_17[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_17[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_17[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_17[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_17[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_17[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_17[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_17[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_17[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_17[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_17[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_17[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_17[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_17[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_17[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_17[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_17[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_17[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_17[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_17[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_17[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_17[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_17[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_17[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_17[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_17[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_17_bits_offset =
    tryToRead_17[0] & input_0_bits_offset_0 | tryToRead_17[1] & input_1_bits_offset_0 | tryToRead_17[2] & input_2_bits_offset_0 | tryToRead_17[3] & input_3_bits_offset_0 | tryToRead_17[4] & input_4_bits_offset_0 | tryToRead_17[5]
    & input_5_bits_offset_0 | tryToRead_17[6] & input_6_bits_offset_0 | tryToRead_17[7] & input_7_bits_offset_0 | tryToRead_17[8] & input_8_bits_offset_0 | tryToRead_17[9] & input_9_bits_offset_0 | tryToRead_17[10] & input_10_bits_offset_0
    | tryToRead_17[11] & input_11_bits_offset_0 | tryToRead_17[12] & input_12_bits_offset_0 | tryToRead_17[13] & input_13_bits_offset_0 | tryToRead_17[14] & input_14_bits_offset_0 | tryToRead_17[15] & input_15_bits_offset_0
    | tryToRead_17[16] & input_16_bits_offset_0 | tryToRead_17[17] & input_17_bits_offset_0 | tryToRead_17[18] & input_18_bits_offset_0 | tryToRead_17[19] & input_19_bits_offset_0 | tryToRead_17[20] & input_20_bits_offset_0
    | tryToRead_17[21] & input_21_bits_offset_0 | tryToRead_17[22] & input_22_bits_offset_0 | tryToRead_17[23] & input_23_bits_offset_0 | tryToRead_17[24] & input_24_bits_offset_0 | tryToRead_17[25] & input_25_bits_offset_0
    | tryToRead_17[26] & input_26_bits_offset_0 | tryToRead_17[27] & input_27_bits_offset_0 | tryToRead_17[28] & input_28_bits_offset_0 | tryToRead_17[29] & input_29_bits_offset_0 | tryToRead_17[30] & input_30_bits_offset_0
    | tryToRead_17[31] & input_31_bits_offset_0;
  assign selectReq_17_bits_vs =
    (tryToRead_17[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_17[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_17[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_17[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_17[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_17[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_17[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_17[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_17[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_17[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_17[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_17[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_17[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_17[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_17[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_17[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_17[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_17[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_17[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_17[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_17[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_17[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_17[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_17[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_17[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_17[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_17[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_17[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_17[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_17[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_17[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_17[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_17_valid =
    tryToRead_17[0] & input_0_valid_0 | tryToRead_17[1] & input_1_valid_0 | tryToRead_17[2] & input_2_valid_0 | tryToRead_17[3] & input_3_valid_0 | tryToRead_17[4] & input_4_valid_0 | tryToRead_17[5] & input_5_valid_0 | tryToRead_17[6]
    & input_6_valid_0 | tryToRead_17[7] & input_7_valid_0 | tryToRead_17[8] & input_8_valid_0 | tryToRead_17[9] & input_9_valid_0 | tryToRead_17[10] & input_10_valid_0 | tryToRead_17[11] & input_11_valid_0 | tryToRead_17[12]
    & input_12_valid_0 | tryToRead_17[13] & input_13_valid_0 | tryToRead_17[14] & input_14_valid_0 | tryToRead_17[15] & input_15_valid_0 | tryToRead_17[16] & input_16_valid_0 | tryToRead_17[17] & input_17_valid_0 | tryToRead_17[18]
    & input_18_valid_0 | tryToRead_17[19] & input_19_valid_0 | tryToRead_17[20] & input_20_valid_0 | tryToRead_17[21] & input_21_valid_0 | tryToRead_17[22] & input_22_valid_0 | tryToRead_17[23] & input_23_valid_0 | tryToRead_17[24]
    & input_24_valid_0 | tryToRead_17[25] & input_25_valid_0 | tryToRead_17[26] & input_26_valid_0 | tryToRead_17[27] & input_27_valid_0 | tryToRead_17[28] & input_28_valid_0 | tryToRead_17[29] & input_29_valid_0 | tryToRead_17[30]
    & input_30_valid_0 | tryToRead_17[31] & input_31_valid_0;
  wire        selectReq_17_ready =
    tryToRead_17[0] & input_0_ready_0 | tryToRead_17[1] & input_1_ready_0 | tryToRead_17[2] & input_2_ready_0 | tryToRead_17[3] & input_3_ready_0 | tryToRead_17[4] & input_4_ready_0 | tryToRead_17[5] & input_5_ready_0 | tryToRead_17[6]
    & input_6_ready_0 | tryToRead_17[7] & input_7_ready_0 | tryToRead_17[8] & input_8_ready_0 | tryToRead_17[9] & input_9_ready_0 | tryToRead_17[10] & input_10_ready_0 | tryToRead_17[11] & input_11_ready_0 | tryToRead_17[12]
    & input_12_ready_0 | tryToRead_17[13] & input_13_ready_0 | tryToRead_17[14] & input_14_ready_0 | tryToRead_17[15] & input_15_ready_0 | tryToRead_17[16] & input_16_ready_0 | tryToRead_17[17] & input_17_ready_0 | tryToRead_17[18]
    & input_18_ready_0 | tryToRead_17[19] & input_19_ready_0 | tryToRead_17[20] & input_20_ready_0 | tryToRead_17[21] & input_21_ready_0 | tryToRead_17[22] & input_22_ready_0 | tryToRead_17[23] & input_23_ready_0 | tryToRead_17[24]
    & input_24_ready_0 | tryToRead_17[25] & input_25_ready_0 | tryToRead_17[26] & input_26_ready_0 | tryToRead_17[27] & input_27_ready_0 | tryToRead_17[28] & input_28_ready_0 | tryToRead_17[29] & input_29_ready_0 | tryToRead_17[30]
    & input_30_ready_0 | tryToRead_17[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_18 = {inputSelect1H_1[18], inputSelect1H_0[18]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_18 = {inputSelect1H_3[18], inputSelect1H_2[18]};
  wire [3:0]  tryToRead_lo_lo_lo_18 = {tryToRead_lo_lo_lo_hi_18, tryToRead_lo_lo_lo_lo_18};
  wire [1:0]  tryToRead_lo_lo_hi_lo_18 = {inputSelect1H_5[18], inputSelect1H_4[18]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_18 = {inputSelect1H_7[18], inputSelect1H_6[18]};
  wire [3:0]  tryToRead_lo_lo_hi_18 = {tryToRead_lo_lo_hi_hi_18, tryToRead_lo_lo_hi_lo_18};
  wire [7:0]  tryToRead_lo_lo_18 = {tryToRead_lo_lo_hi_18, tryToRead_lo_lo_lo_18};
  wire [1:0]  tryToRead_lo_hi_lo_lo_18 = {inputSelect1H_9[18], inputSelect1H_8[18]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_18 = {inputSelect1H_11[18], inputSelect1H_10[18]};
  wire [3:0]  tryToRead_lo_hi_lo_18 = {tryToRead_lo_hi_lo_hi_18, tryToRead_lo_hi_lo_lo_18};
  wire [1:0]  tryToRead_lo_hi_hi_lo_18 = {inputSelect1H_13[18], inputSelect1H_12[18]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_18 = {inputSelect1H_15[18], inputSelect1H_14[18]};
  wire [3:0]  tryToRead_lo_hi_hi_18 = {tryToRead_lo_hi_hi_hi_18, tryToRead_lo_hi_hi_lo_18};
  wire [7:0]  tryToRead_lo_hi_18 = {tryToRead_lo_hi_hi_18, tryToRead_lo_hi_lo_18};
  wire [15:0] tryToRead_lo_18 = {tryToRead_lo_hi_18, tryToRead_lo_lo_18};
  wire [1:0]  tryToRead_hi_lo_lo_lo_18 = {inputSelect1H_17[18], inputSelect1H_16[18]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_18 = {inputSelect1H_19[18], inputSelect1H_18[18]};
  wire [3:0]  tryToRead_hi_lo_lo_18 = {tryToRead_hi_lo_lo_hi_18, tryToRead_hi_lo_lo_lo_18};
  wire [1:0]  tryToRead_hi_lo_hi_lo_18 = {inputSelect1H_21[18], inputSelect1H_20[18]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_18 = {inputSelect1H_23[18], inputSelect1H_22[18]};
  wire [3:0]  tryToRead_hi_lo_hi_18 = {tryToRead_hi_lo_hi_hi_18, tryToRead_hi_lo_hi_lo_18};
  wire [7:0]  tryToRead_hi_lo_18 = {tryToRead_hi_lo_hi_18, tryToRead_hi_lo_lo_18};
  wire [1:0]  tryToRead_hi_hi_lo_lo_18 = {inputSelect1H_25[18], inputSelect1H_24[18]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_18 = {inputSelect1H_27[18], inputSelect1H_26[18]};
  wire [3:0]  tryToRead_hi_hi_lo_18 = {tryToRead_hi_hi_lo_hi_18, tryToRead_hi_hi_lo_lo_18};
  wire [1:0]  tryToRead_hi_hi_hi_lo_18 = {inputSelect1H_29[18], inputSelect1H_28[18]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_18 = {inputSelect1H_31[18], inputSelect1H_30[18]};
  wire [3:0]  tryToRead_hi_hi_hi_18 = {tryToRead_hi_hi_hi_hi_18, tryToRead_hi_hi_hi_lo_18};
  wire [7:0]  tryToRead_hi_hi_18 = {tryToRead_hi_hi_hi_18, tryToRead_hi_hi_lo_18};
  wire [15:0] tryToRead_hi_18 = {tryToRead_hi_hi_18, tryToRead_hi_lo_18};
  wire [31:0] tryToRead_18 = {tryToRead_hi_18, tryToRead_lo_18};
  wire        output_18_valid_0 = |tryToRead_18;
  wire [4:0]  output_18_bits_vs_0 = selectReq_18_bits_vs;
  wire        output_18_bits_offset_0 = selectReq_18_bits_offset;
  wire [4:0]  output_18_bits_writeIndex_0 = selectReq_18_bits_requestIndex;
  wire [1:0]  output_18_bits_dataOffset_0 = selectReq_18_bits_dataOffset;
  assign selectReq_18_bits_dataOffset =
    (tryToRead_18[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_18[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_18[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_18[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_18[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_18[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_18[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_18[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_18[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_18[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_18[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_18[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_18[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_18[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_18[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_18[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_18[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_18[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_18[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_18[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_18[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_18[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_18[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_18[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_18[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_18[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_18_bits_requestIndex =
    {4'h0, tryToRead_18[1]} | {3'h0, tryToRead_18[2], 1'h0} | (tryToRead_18[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_18[4], 2'h0} | (tryToRead_18[5] ? 5'h5 : 5'h0) | (tryToRead_18[6] ? 5'h6 : 5'h0) | (tryToRead_18[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_18[8], 3'h0} | (tryToRead_18[9] ? 5'h9 : 5'h0) | (tryToRead_18[10] ? 5'hA : 5'h0) | (tryToRead_18[11] ? 5'hB : 5'h0) | (tryToRead_18[12] ? 5'hC : 5'h0) | (tryToRead_18[13] ? 5'hD : 5'h0)
    | (tryToRead_18[14] ? 5'hE : 5'h0) | (tryToRead_18[15] ? 5'hF : 5'h0) | {tryToRead_18[16], 4'h0} | (tryToRead_18[17] ? 5'h11 : 5'h0) | (tryToRead_18[18] ? 5'h12 : 5'h0) | (tryToRead_18[19] ? 5'h13 : 5'h0)
    | (tryToRead_18[20] ? 5'h14 : 5'h0) | (tryToRead_18[21] ? 5'h15 : 5'h0) | (tryToRead_18[22] ? 5'h16 : 5'h0) | (tryToRead_18[23] ? 5'h17 : 5'h0) | (tryToRead_18[24] ? 5'h18 : 5'h0) | (tryToRead_18[25] ? 5'h19 : 5'h0)
    | (tryToRead_18[26] ? 5'h1A : 5'h0) | (tryToRead_18[27] ? 5'h1B : 5'h0) | (tryToRead_18[28] ? 5'h1C : 5'h0) | (tryToRead_18[29] ? 5'h1D : 5'h0) | (tryToRead_18[30] ? 5'h1E : 5'h0) | {5{tryToRead_18[31]}};
  wire [4:0]  selectReq_18_bits_readLane =
    (tryToRead_18[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_18[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_18[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_18[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_18[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_18[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_18[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_18[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_18[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_18[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_18[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_18[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_18[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_18[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_18[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_18[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_18[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_18[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_18[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_18[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_18[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_18[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_18[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_18[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_18[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_18[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_18[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_18[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_18[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_18[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_18[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_18[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_18_bits_offset =
    tryToRead_18[0] & input_0_bits_offset_0 | tryToRead_18[1] & input_1_bits_offset_0 | tryToRead_18[2] & input_2_bits_offset_0 | tryToRead_18[3] & input_3_bits_offset_0 | tryToRead_18[4] & input_4_bits_offset_0 | tryToRead_18[5]
    & input_5_bits_offset_0 | tryToRead_18[6] & input_6_bits_offset_0 | tryToRead_18[7] & input_7_bits_offset_0 | tryToRead_18[8] & input_8_bits_offset_0 | tryToRead_18[9] & input_9_bits_offset_0 | tryToRead_18[10] & input_10_bits_offset_0
    | tryToRead_18[11] & input_11_bits_offset_0 | tryToRead_18[12] & input_12_bits_offset_0 | tryToRead_18[13] & input_13_bits_offset_0 | tryToRead_18[14] & input_14_bits_offset_0 | tryToRead_18[15] & input_15_bits_offset_0
    | tryToRead_18[16] & input_16_bits_offset_0 | tryToRead_18[17] & input_17_bits_offset_0 | tryToRead_18[18] & input_18_bits_offset_0 | tryToRead_18[19] & input_19_bits_offset_0 | tryToRead_18[20] & input_20_bits_offset_0
    | tryToRead_18[21] & input_21_bits_offset_0 | tryToRead_18[22] & input_22_bits_offset_0 | tryToRead_18[23] & input_23_bits_offset_0 | tryToRead_18[24] & input_24_bits_offset_0 | tryToRead_18[25] & input_25_bits_offset_0
    | tryToRead_18[26] & input_26_bits_offset_0 | tryToRead_18[27] & input_27_bits_offset_0 | tryToRead_18[28] & input_28_bits_offset_0 | tryToRead_18[29] & input_29_bits_offset_0 | tryToRead_18[30] & input_30_bits_offset_0
    | tryToRead_18[31] & input_31_bits_offset_0;
  assign selectReq_18_bits_vs =
    (tryToRead_18[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_18[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_18[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_18[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_18[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_18[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_18[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_18[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_18[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_18[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_18[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_18[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_18[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_18[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_18[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_18[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_18[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_18[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_18[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_18[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_18[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_18[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_18[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_18[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_18[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_18[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_18[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_18[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_18[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_18[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_18[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_18[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_18_valid =
    tryToRead_18[0] & input_0_valid_0 | tryToRead_18[1] & input_1_valid_0 | tryToRead_18[2] & input_2_valid_0 | tryToRead_18[3] & input_3_valid_0 | tryToRead_18[4] & input_4_valid_0 | tryToRead_18[5] & input_5_valid_0 | tryToRead_18[6]
    & input_6_valid_0 | tryToRead_18[7] & input_7_valid_0 | tryToRead_18[8] & input_8_valid_0 | tryToRead_18[9] & input_9_valid_0 | tryToRead_18[10] & input_10_valid_0 | tryToRead_18[11] & input_11_valid_0 | tryToRead_18[12]
    & input_12_valid_0 | tryToRead_18[13] & input_13_valid_0 | tryToRead_18[14] & input_14_valid_0 | tryToRead_18[15] & input_15_valid_0 | tryToRead_18[16] & input_16_valid_0 | tryToRead_18[17] & input_17_valid_0 | tryToRead_18[18]
    & input_18_valid_0 | tryToRead_18[19] & input_19_valid_0 | tryToRead_18[20] & input_20_valid_0 | tryToRead_18[21] & input_21_valid_0 | tryToRead_18[22] & input_22_valid_0 | tryToRead_18[23] & input_23_valid_0 | tryToRead_18[24]
    & input_24_valid_0 | tryToRead_18[25] & input_25_valid_0 | tryToRead_18[26] & input_26_valid_0 | tryToRead_18[27] & input_27_valid_0 | tryToRead_18[28] & input_28_valid_0 | tryToRead_18[29] & input_29_valid_0 | tryToRead_18[30]
    & input_30_valid_0 | tryToRead_18[31] & input_31_valid_0;
  wire        selectReq_18_ready =
    tryToRead_18[0] & input_0_ready_0 | tryToRead_18[1] & input_1_ready_0 | tryToRead_18[2] & input_2_ready_0 | tryToRead_18[3] & input_3_ready_0 | tryToRead_18[4] & input_4_ready_0 | tryToRead_18[5] & input_5_ready_0 | tryToRead_18[6]
    & input_6_ready_0 | tryToRead_18[7] & input_7_ready_0 | tryToRead_18[8] & input_8_ready_0 | tryToRead_18[9] & input_9_ready_0 | tryToRead_18[10] & input_10_ready_0 | tryToRead_18[11] & input_11_ready_0 | tryToRead_18[12]
    & input_12_ready_0 | tryToRead_18[13] & input_13_ready_0 | tryToRead_18[14] & input_14_ready_0 | tryToRead_18[15] & input_15_ready_0 | tryToRead_18[16] & input_16_ready_0 | tryToRead_18[17] & input_17_ready_0 | tryToRead_18[18]
    & input_18_ready_0 | tryToRead_18[19] & input_19_ready_0 | tryToRead_18[20] & input_20_ready_0 | tryToRead_18[21] & input_21_ready_0 | tryToRead_18[22] & input_22_ready_0 | tryToRead_18[23] & input_23_ready_0 | tryToRead_18[24]
    & input_24_ready_0 | tryToRead_18[25] & input_25_ready_0 | tryToRead_18[26] & input_26_ready_0 | tryToRead_18[27] & input_27_ready_0 | tryToRead_18[28] & input_28_ready_0 | tryToRead_18[29] & input_29_ready_0 | tryToRead_18[30]
    & input_30_ready_0 | tryToRead_18[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_19 = {inputSelect1H_1[19], inputSelect1H_0[19]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_19 = {inputSelect1H_3[19], inputSelect1H_2[19]};
  wire [3:0]  tryToRead_lo_lo_lo_19 = {tryToRead_lo_lo_lo_hi_19, tryToRead_lo_lo_lo_lo_19};
  wire [1:0]  tryToRead_lo_lo_hi_lo_19 = {inputSelect1H_5[19], inputSelect1H_4[19]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_19 = {inputSelect1H_7[19], inputSelect1H_6[19]};
  wire [3:0]  tryToRead_lo_lo_hi_19 = {tryToRead_lo_lo_hi_hi_19, tryToRead_lo_lo_hi_lo_19};
  wire [7:0]  tryToRead_lo_lo_19 = {tryToRead_lo_lo_hi_19, tryToRead_lo_lo_lo_19};
  wire [1:0]  tryToRead_lo_hi_lo_lo_19 = {inputSelect1H_9[19], inputSelect1H_8[19]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_19 = {inputSelect1H_11[19], inputSelect1H_10[19]};
  wire [3:0]  tryToRead_lo_hi_lo_19 = {tryToRead_lo_hi_lo_hi_19, tryToRead_lo_hi_lo_lo_19};
  wire [1:0]  tryToRead_lo_hi_hi_lo_19 = {inputSelect1H_13[19], inputSelect1H_12[19]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_19 = {inputSelect1H_15[19], inputSelect1H_14[19]};
  wire [3:0]  tryToRead_lo_hi_hi_19 = {tryToRead_lo_hi_hi_hi_19, tryToRead_lo_hi_hi_lo_19};
  wire [7:0]  tryToRead_lo_hi_19 = {tryToRead_lo_hi_hi_19, tryToRead_lo_hi_lo_19};
  wire [15:0] tryToRead_lo_19 = {tryToRead_lo_hi_19, tryToRead_lo_lo_19};
  wire [1:0]  tryToRead_hi_lo_lo_lo_19 = {inputSelect1H_17[19], inputSelect1H_16[19]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_19 = {inputSelect1H_19[19], inputSelect1H_18[19]};
  wire [3:0]  tryToRead_hi_lo_lo_19 = {tryToRead_hi_lo_lo_hi_19, tryToRead_hi_lo_lo_lo_19};
  wire [1:0]  tryToRead_hi_lo_hi_lo_19 = {inputSelect1H_21[19], inputSelect1H_20[19]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_19 = {inputSelect1H_23[19], inputSelect1H_22[19]};
  wire [3:0]  tryToRead_hi_lo_hi_19 = {tryToRead_hi_lo_hi_hi_19, tryToRead_hi_lo_hi_lo_19};
  wire [7:0]  tryToRead_hi_lo_19 = {tryToRead_hi_lo_hi_19, tryToRead_hi_lo_lo_19};
  wire [1:0]  tryToRead_hi_hi_lo_lo_19 = {inputSelect1H_25[19], inputSelect1H_24[19]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_19 = {inputSelect1H_27[19], inputSelect1H_26[19]};
  wire [3:0]  tryToRead_hi_hi_lo_19 = {tryToRead_hi_hi_lo_hi_19, tryToRead_hi_hi_lo_lo_19};
  wire [1:0]  tryToRead_hi_hi_hi_lo_19 = {inputSelect1H_29[19], inputSelect1H_28[19]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_19 = {inputSelect1H_31[19], inputSelect1H_30[19]};
  wire [3:0]  tryToRead_hi_hi_hi_19 = {tryToRead_hi_hi_hi_hi_19, tryToRead_hi_hi_hi_lo_19};
  wire [7:0]  tryToRead_hi_hi_19 = {tryToRead_hi_hi_hi_19, tryToRead_hi_hi_lo_19};
  wire [15:0] tryToRead_hi_19 = {tryToRead_hi_hi_19, tryToRead_hi_lo_19};
  wire [31:0] tryToRead_19 = {tryToRead_hi_19, tryToRead_lo_19};
  wire        output_19_valid_0 = |tryToRead_19;
  wire [4:0]  output_19_bits_vs_0 = selectReq_19_bits_vs;
  wire        output_19_bits_offset_0 = selectReq_19_bits_offset;
  wire [4:0]  output_19_bits_writeIndex_0 = selectReq_19_bits_requestIndex;
  wire [1:0]  output_19_bits_dataOffset_0 = selectReq_19_bits_dataOffset;
  assign selectReq_19_bits_dataOffset =
    (tryToRead_19[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_19[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_19[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_19[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_19[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_19[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_19[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_19[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_19[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_19[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_19[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_19[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_19[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_19[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_19[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_19[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_19[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_19[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_19[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_19[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_19[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_19[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_19[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_19[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_19[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_19[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_19_bits_requestIndex =
    {4'h0, tryToRead_19[1]} | {3'h0, tryToRead_19[2], 1'h0} | (tryToRead_19[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_19[4], 2'h0} | (tryToRead_19[5] ? 5'h5 : 5'h0) | (tryToRead_19[6] ? 5'h6 : 5'h0) | (tryToRead_19[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_19[8], 3'h0} | (tryToRead_19[9] ? 5'h9 : 5'h0) | (tryToRead_19[10] ? 5'hA : 5'h0) | (tryToRead_19[11] ? 5'hB : 5'h0) | (tryToRead_19[12] ? 5'hC : 5'h0) | (tryToRead_19[13] ? 5'hD : 5'h0)
    | (tryToRead_19[14] ? 5'hE : 5'h0) | (tryToRead_19[15] ? 5'hF : 5'h0) | {tryToRead_19[16], 4'h0} | (tryToRead_19[17] ? 5'h11 : 5'h0) | (tryToRead_19[18] ? 5'h12 : 5'h0) | (tryToRead_19[19] ? 5'h13 : 5'h0)
    | (tryToRead_19[20] ? 5'h14 : 5'h0) | (tryToRead_19[21] ? 5'h15 : 5'h0) | (tryToRead_19[22] ? 5'h16 : 5'h0) | (tryToRead_19[23] ? 5'h17 : 5'h0) | (tryToRead_19[24] ? 5'h18 : 5'h0) | (tryToRead_19[25] ? 5'h19 : 5'h0)
    | (tryToRead_19[26] ? 5'h1A : 5'h0) | (tryToRead_19[27] ? 5'h1B : 5'h0) | (tryToRead_19[28] ? 5'h1C : 5'h0) | (tryToRead_19[29] ? 5'h1D : 5'h0) | (tryToRead_19[30] ? 5'h1E : 5'h0) | {5{tryToRead_19[31]}};
  wire [4:0]  selectReq_19_bits_readLane =
    (tryToRead_19[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_19[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_19[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_19[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_19[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_19[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_19[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_19[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_19[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_19[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_19[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_19[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_19[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_19[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_19[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_19[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_19[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_19[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_19[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_19[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_19[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_19[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_19[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_19[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_19[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_19[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_19[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_19[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_19[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_19[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_19[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_19[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_19_bits_offset =
    tryToRead_19[0] & input_0_bits_offset_0 | tryToRead_19[1] & input_1_bits_offset_0 | tryToRead_19[2] & input_2_bits_offset_0 | tryToRead_19[3] & input_3_bits_offset_0 | tryToRead_19[4] & input_4_bits_offset_0 | tryToRead_19[5]
    & input_5_bits_offset_0 | tryToRead_19[6] & input_6_bits_offset_0 | tryToRead_19[7] & input_7_bits_offset_0 | tryToRead_19[8] & input_8_bits_offset_0 | tryToRead_19[9] & input_9_bits_offset_0 | tryToRead_19[10] & input_10_bits_offset_0
    | tryToRead_19[11] & input_11_bits_offset_0 | tryToRead_19[12] & input_12_bits_offset_0 | tryToRead_19[13] & input_13_bits_offset_0 | tryToRead_19[14] & input_14_bits_offset_0 | tryToRead_19[15] & input_15_bits_offset_0
    | tryToRead_19[16] & input_16_bits_offset_0 | tryToRead_19[17] & input_17_bits_offset_0 | tryToRead_19[18] & input_18_bits_offset_0 | tryToRead_19[19] & input_19_bits_offset_0 | tryToRead_19[20] & input_20_bits_offset_0
    | tryToRead_19[21] & input_21_bits_offset_0 | tryToRead_19[22] & input_22_bits_offset_0 | tryToRead_19[23] & input_23_bits_offset_0 | tryToRead_19[24] & input_24_bits_offset_0 | tryToRead_19[25] & input_25_bits_offset_0
    | tryToRead_19[26] & input_26_bits_offset_0 | tryToRead_19[27] & input_27_bits_offset_0 | tryToRead_19[28] & input_28_bits_offset_0 | tryToRead_19[29] & input_29_bits_offset_0 | tryToRead_19[30] & input_30_bits_offset_0
    | tryToRead_19[31] & input_31_bits_offset_0;
  assign selectReq_19_bits_vs =
    (tryToRead_19[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_19[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_19[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_19[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_19[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_19[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_19[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_19[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_19[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_19[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_19[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_19[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_19[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_19[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_19[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_19[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_19[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_19[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_19[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_19[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_19[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_19[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_19[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_19[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_19[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_19[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_19[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_19[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_19[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_19[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_19[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_19[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_19_valid =
    tryToRead_19[0] & input_0_valid_0 | tryToRead_19[1] & input_1_valid_0 | tryToRead_19[2] & input_2_valid_0 | tryToRead_19[3] & input_3_valid_0 | tryToRead_19[4] & input_4_valid_0 | tryToRead_19[5] & input_5_valid_0 | tryToRead_19[6]
    & input_6_valid_0 | tryToRead_19[7] & input_7_valid_0 | tryToRead_19[8] & input_8_valid_0 | tryToRead_19[9] & input_9_valid_0 | tryToRead_19[10] & input_10_valid_0 | tryToRead_19[11] & input_11_valid_0 | tryToRead_19[12]
    & input_12_valid_0 | tryToRead_19[13] & input_13_valid_0 | tryToRead_19[14] & input_14_valid_0 | tryToRead_19[15] & input_15_valid_0 | tryToRead_19[16] & input_16_valid_0 | tryToRead_19[17] & input_17_valid_0 | tryToRead_19[18]
    & input_18_valid_0 | tryToRead_19[19] & input_19_valid_0 | tryToRead_19[20] & input_20_valid_0 | tryToRead_19[21] & input_21_valid_0 | tryToRead_19[22] & input_22_valid_0 | tryToRead_19[23] & input_23_valid_0 | tryToRead_19[24]
    & input_24_valid_0 | tryToRead_19[25] & input_25_valid_0 | tryToRead_19[26] & input_26_valid_0 | tryToRead_19[27] & input_27_valid_0 | tryToRead_19[28] & input_28_valid_0 | tryToRead_19[29] & input_29_valid_0 | tryToRead_19[30]
    & input_30_valid_0 | tryToRead_19[31] & input_31_valid_0;
  wire        selectReq_19_ready =
    tryToRead_19[0] & input_0_ready_0 | tryToRead_19[1] & input_1_ready_0 | tryToRead_19[2] & input_2_ready_0 | tryToRead_19[3] & input_3_ready_0 | tryToRead_19[4] & input_4_ready_0 | tryToRead_19[5] & input_5_ready_0 | tryToRead_19[6]
    & input_6_ready_0 | tryToRead_19[7] & input_7_ready_0 | tryToRead_19[8] & input_8_ready_0 | tryToRead_19[9] & input_9_ready_0 | tryToRead_19[10] & input_10_ready_0 | tryToRead_19[11] & input_11_ready_0 | tryToRead_19[12]
    & input_12_ready_0 | tryToRead_19[13] & input_13_ready_0 | tryToRead_19[14] & input_14_ready_0 | tryToRead_19[15] & input_15_ready_0 | tryToRead_19[16] & input_16_ready_0 | tryToRead_19[17] & input_17_ready_0 | tryToRead_19[18]
    & input_18_ready_0 | tryToRead_19[19] & input_19_ready_0 | tryToRead_19[20] & input_20_ready_0 | tryToRead_19[21] & input_21_ready_0 | tryToRead_19[22] & input_22_ready_0 | tryToRead_19[23] & input_23_ready_0 | tryToRead_19[24]
    & input_24_ready_0 | tryToRead_19[25] & input_25_ready_0 | tryToRead_19[26] & input_26_ready_0 | tryToRead_19[27] & input_27_ready_0 | tryToRead_19[28] & input_28_ready_0 | tryToRead_19[29] & input_29_ready_0 | tryToRead_19[30]
    & input_30_ready_0 | tryToRead_19[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_20 = {inputSelect1H_1[20], inputSelect1H_0[20]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_20 = {inputSelect1H_3[20], inputSelect1H_2[20]};
  wire [3:0]  tryToRead_lo_lo_lo_20 = {tryToRead_lo_lo_lo_hi_20, tryToRead_lo_lo_lo_lo_20};
  wire [1:0]  tryToRead_lo_lo_hi_lo_20 = {inputSelect1H_5[20], inputSelect1H_4[20]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_20 = {inputSelect1H_7[20], inputSelect1H_6[20]};
  wire [3:0]  tryToRead_lo_lo_hi_20 = {tryToRead_lo_lo_hi_hi_20, tryToRead_lo_lo_hi_lo_20};
  wire [7:0]  tryToRead_lo_lo_20 = {tryToRead_lo_lo_hi_20, tryToRead_lo_lo_lo_20};
  wire [1:0]  tryToRead_lo_hi_lo_lo_20 = {inputSelect1H_9[20], inputSelect1H_8[20]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_20 = {inputSelect1H_11[20], inputSelect1H_10[20]};
  wire [3:0]  tryToRead_lo_hi_lo_20 = {tryToRead_lo_hi_lo_hi_20, tryToRead_lo_hi_lo_lo_20};
  wire [1:0]  tryToRead_lo_hi_hi_lo_20 = {inputSelect1H_13[20], inputSelect1H_12[20]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_20 = {inputSelect1H_15[20], inputSelect1H_14[20]};
  wire [3:0]  tryToRead_lo_hi_hi_20 = {tryToRead_lo_hi_hi_hi_20, tryToRead_lo_hi_hi_lo_20};
  wire [7:0]  tryToRead_lo_hi_20 = {tryToRead_lo_hi_hi_20, tryToRead_lo_hi_lo_20};
  wire [15:0] tryToRead_lo_20 = {tryToRead_lo_hi_20, tryToRead_lo_lo_20};
  wire [1:0]  tryToRead_hi_lo_lo_lo_20 = {inputSelect1H_17[20], inputSelect1H_16[20]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_20 = {inputSelect1H_19[20], inputSelect1H_18[20]};
  wire [3:0]  tryToRead_hi_lo_lo_20 = {tryToRead_hi_lo_lo_hi_20, tryToRead_hi_lo_lo_lo_20};
  wire [1:0]  tryToRead_hi_lo_hi_lo_20 = {inputSelect1H_21[20], inputSelect1H_20[20]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_20 = {inputSelect1H_23[20], inputSelect1H_22[20]};
  wire [3:0]  tryToRead_hi_lo_hi_20 = {tryToRead_hi_lo_hi_hi_20, tryToRead_hi_lo_hi_lo_20};
  wire [7:0]  tryToRead_hi_lo_20 = {tryToRead_hi_lo_hi_20, tryToRead_hi_lo_lo_20};
  wire [1:0]  tryToRead_hi_hi_lo_lo_20 = {inputSelect1H_25[20], inputSelect1H_24[20]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_20 = {inputSelect1H_27[20], inputSelect1H_26[20]};
  wire [3:0]  tryToRead_hi_hi_lo_20 = {tryToRead_hi_hi_lo_hi_20, tryToRead_hi_hi_lo_lo_20};
  wire [1:0]  tryToRead_hi_hi_hi_lo_20 = {inputSelect1H_29[20], inputSelect1H_28[20]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_20 = {inputSelect1H_31[20], inputSelect1H_30[20]};
  wire [3:0]  tryToRead_hi_hi_hi_20 = {tryToRead_hi_hi_hi_hi_20, tryToRead_hi_hi_hi_lo_20};
  wire [7:0]  tryToRead_hi_hi_20 = {tryToRead_hi_hi_hi_20, tryToRead_hi_hi_lo_20};
  wire [15:0] tryToRead_hi_20 = {tryToRead_hi_hi_20, tryToRead_hi_lo_20};
  wire [31:0] tryToRead_20 = {tryToRead_hi_20, tryToRead_lo_20};
  wire        output_20_valid_0 = |tryToRead_20;
  wire [4:0]  output_20_bits_vs_0 = selectReq_20_bits_vs;
  wire        output_20_bits_offset_0 = selectReq_20_bits_offset;
  wire [4:0]  output_20_bits_writeIndex_0 = selectReq_20_bits_requestIndex;
  wire [1:0]  output_20_bits_dataOffset_0 = selectReq_20_bits_dataOffset;
  assign selectReq_20_bits_dataOffset =
    (tryToRead_20[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_20[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_20[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_20[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_20[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_20[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_20[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_20[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_20[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_20[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_20[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_20[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_20[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_20[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_20[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_20[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_20[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_20[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_20[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_20[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_20[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_20[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_20[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_20[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_20[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_20[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_20_bits_requestIndex =
    {4'h0, tryToRead_20[1]} | {3'h0, tryToRead_20[2], 1'h0} | (tryToRead_20[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_20[4], 2'h0} | (tryToRead_20[5] ? 5'h5 : 5'h0) | (tryToRead_20[6] ? 5'h6 : 5'h0) | (tryToRead_20[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_20[8], 3'h0} | (tryToRead_20[9] ? 5'h9 : 5'h0) | (tryToRead_20[10] ? 5'hA : 5'h0) | (tryToRead_20[11] ? 5'hB : 5'h0) | (tryToRead_20[12] ? 5'hC : 5'h0) | (tryToRead_20[13] ? 5'hD : 5'h0)
    | (tryToRead_20[14] ? 5'hE : 5'h0) | (tryToRead_20[15] ? 5'hF : 5'h0) | {tryToRead_20[16], 4'h0} | (tryToRead_20[17] ? 5'h11 : 5'h0) | (tryToRead_20[18] ? 5'h12 : 5'h0) | (tryToRead_20[19] ? 5'h13 : 5'h0)
    | (tryToRead_20[20] ? 5'h14 : 5'h0) | (tryToRead_20[21] ? 5'h15 : 5'h0) | (tryToRead_20[22] ? 5'h16 : 5'h0) | (tryToRead_20[23] ? 5'h17 : 5'h0) | (tryToRead_20[24] ? 5'h18 : 5'h0) | (tryToRead_20[25] ? 5'h19 : 5'h0)
    | (tryToRead_20[26] ? 5'h1A : 5'h0) | (tryToRead_20[27] ? 5'h1B : 5'h0) | (tryToRead_20[28] ? 5'h1C : 5'h0) | (tryToRead_20[29] ? 5'h1D : 5'h0) | (tryToRead_20[30] ? 5'h1E : 5'h0) | {5{tryToRead_20[31]}};
  wire [4:0]  selectReq_20_bits_readLane =
    (tryToRead_20[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_20[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_20[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_20[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_20[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_20[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_20[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_20[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_20[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_20[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_20[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_20[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_20[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_20[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_20[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_20[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_20[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_20[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_20[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_20[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_20[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_20[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_20[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_20[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_20[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_20[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_20[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_20[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_20[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_20[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_20[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_20[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_20_bits_offset =
    tryToRead_20[0] & input_0_bits_offset_0 | tryToRead_20[1] & input_1_bits_offset_0 | tryToRead_20[2] & input_2_bits_offset_0 | tryToRead_20[3] & input_3_bits_offset_0 | tryToRead_20[4] & input_4_bits_offset_0 | tryToRead_20[5]
    & input_5_bits_offset_0 | tryToRead_20[6] & input_6_bits_offset_0 | tryToRead_20[7] & input_7_bits_offset_0 | tryToRead_20[8] & input_8_bits_offset_0 | tryToRead_20[9] & input_9_bits_offset_0 | tryToRead_20[10] & input_10_bits_offset_0
    | tryToRead_20[11] & input_11_bits_offset_0 | tryToRead_20[12] & input_12_bits_offset_0 | tryToRead_20[13] & input_13_bits_offset_0 | tryToRead_20[14] & input_14_bits_offset_0 | tryToRead_20[15] & input_15_bits_offset_0
    | tryToRead_20[16] & input_16_bits_offset_0 | tryToRead_20[17] & input_17_bits_offset_0 | tryToRead_20[18] & input_18_bits_offset_0 | tryToRead_20[19] & input_19_bits_offset_0 | tryToRead_20[20] & input_20_bits_offset_0
    | tryToRead_20[21] & input_21_bits_offset_0 | tryToRead_20[22] & input_22_bits_offset_0 | tryToRead_20[23] & input_23_bits_offset_0 | tryToRead_20[24] & input_24_bits_offset_0 | tryToRead_20[25] & input_25_bits_offset_0
    | tryToRead_20[26] & input_26_bits_offset_0 | tryToRead_20[27] & input_27_bits_offset_0 | tryToRead_20[28] & input_28_bits_offset_0 | tryToRead_20[29] & input_29_bits_offset_0 | tryToRead_20[30] & input_30_bits_offset_0
    | tryToRead_20[31] & input_31_bits_offset_0;
  assign selectReq_20_bits_vs =
    (tryToRead_20[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_20[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_20[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_20[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_20[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_20[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_20[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_20[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_20[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_20[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_20[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_20[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_20[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_20[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_20[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_20[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_20[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_20[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_20[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_20[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_20[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_20[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_20[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_20[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_20[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_20[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_20[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_20[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_20[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_20[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_20[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_20[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_20_valid =
    tryToRead_20[0] & input_0_valid_0 | tryToRead_20[1] & input_1_valid_0 | tryToRead_20[2] & input_2_valid_0 | tryToRead_20[3] & input_3_valid_0 | tryToRead_20[4] & input_4_valid_0 | tryToRead_20[5] & input_5_valid_0 | tryToRead_20[6]
    & input_6_valid_0 | tryToRead_20[7] & input_7_valid_0 | tryToRead_20[8] & input_8_valid_0 | tryToRead_20[9] & input_9_valid_0 | tryToRead_20[10] & input_10_valid_0 | tryToRead_20[11] & input_11_valid_0 | tryToRead_20[12]
    & input_12_valid_0 | tryToRead_20[13] & input_13_valid_0 | tryToRead_20[14] & input_14_valid_0 | tryToRead_20[15] & input_15_valid_0 | tryToRead_20[16] & input_16_valid_0 | tryToRead_20[17] & input_17_valid_0 | tryToRead_20[18]
    & input_18_valid_0 | tryToRead_20[19] & input_19_valid_0 | tryToRead_20[20] & input_20_valid_0 | tryToRead_20[21] & input_21_valid_0 | tryToRead_20[22] & input_22_valid_0 | tryToRead_20[23] & input_23_valid_0 | tryToRead_20[24]
    & input_24_valid_0 | tryToRead_20[25] & input_25_valid_0 | tryToRead_20[26] & input_26_valid_0 | tryToRead_20[27] & input_27_valid_0 | tryToRead_20[28] & input_28_valid_0 | tryToRead_20[29] & input_29_valid_0 | tryToRead_20[30]
    & input_30_valid_0 | tryToRead_20[31] & input_31_valid_0;
  wire        selectReq_20_ready =
    tryToRead_20[0] & input_0_ready_0 | tryToRead_20[1] & input_1_ready_0 | tryToRead_20[2] & input_2_ready_0 | tryToRead_20[3] & input_3_ready_0 | tryToRead_20[4] & input_4_ready_0 | tryToRead_20[5] & input_5_ready_0 | tryToRead_20[6]
    & input_6_ready_0 | tryToRead_20[7] & input_7_ready_0 | tryToRead_20[8] & input_8_ready_0 | tryToRead_20[9] & input_9_ready_0 | tryToRead_20[10] & input_10_ready_0 | tryToRead_20[11] & input_11_ready_0 | tryToRead_20[12]
    & input_12_ready_0 | tryToRead_20[13] & input_13_ready_0 | tryToRead_20[14] & input_14_ready_0 | tryToRead_20[15] & input_15_ready_0 | tryToRead_20[16] & input_16_ready_0 | tryToRead_20[17] & input_17_ready_0 | tryToRead_20[18]
    & input_18_ready_0 | tryToRead_20[19] & input_19_ready_0 | tryToRead_20[20] & input_20_ready_0 | tryToRead_20[21] & input_21_ready_0 | tryToRead_20[22] & input_22_ready_0 | tryToRead_20[23] & input_23_ready_0 | tryToRead_20[24]
    & input_24_ready_0 | tryToRead_20[25] & input_25_ready_0 | tryToRead_20[26] & input_26_ready_0 | tryToRead_20[27] & input_27_ready_0 | tryToRead_20[28] & input_28_ready_0 | tryToRead_20[29] & input_29_ready_0 | tryToRead_20[30]
    & input_30_ready_0 | tryToRead_20[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_21 = {inputSelect1H_1[21], inputSelect1H_0[21]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_21 = {inputSelect1H_3[21], inputSelect1H_2[21]};
  wire [3:0]  tryToRead_lo_lo_lo_21 = {tryToRead_lo_lo_lo_hi_21, tryToRead_lo_lo_lo_lo_21};
  wire [1:0]  tryToRead_lo_lo_hi_lo_21 = {inputSelect1H_5[21], inputSelect1H_4[21]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_21 = {inputSelect1H_7[21], inputSelect1H_6[21]};
  wire [3:0]  tryToRead_lo_lo_hi_21 = {tryToRead_lo_lo_hi_hi_21, tryToRead_lo_lo_hi_lo_21};
  wire [7:0]  tryToRead_lo_lo_21 = {tryToRead_lo_lo_hi_21, tryToRead_lo_lo_lo_21};
  wire [1:0]  tryToRead_lo_hi_lo_lo_21 = {inputSelect1H_9[21], inputSelect1H_8[21]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_21 = {inputSelect1H_11[21], inputSelect1H_10[21]};
  wire [3:0]  tryToRead_lo_hi_lo_21 = {tryToRead_lo_hi_lo_hi_21, tryToRead_lo_hi_lo_lo_21};
  wire [1:0]  tryToRead_lo_hi_hi_lo_21 = {inputSelect1H_13[21], inputSelect1H_12[21]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_21 = {inputSelect1H_15[21], inputSelect1H_14[21]};
  wire [3:0]  tryToRead_lo_hi_hi_21 = {tryToRead_lo_hi_hi_hi_21, tryToRead_lo_hi_hi_lo_21};
  wire [7:0]  tryToRead_lo_hi_21 = {tryToRead_lo_hi_hi_21, tryToRead_lo_hi_lo_21};
  wire [15:0] tryToRead_lo_21 = {tryToRead_lo_hi_21, tryToRead_lo_lo_21};
  wire [1:0]  tryToRead_hi_lo_lo_lo_21 = {inputSelect1H_17[21], inputSelect1H_16[21]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_21 = {inputSelect1H_19[21], inputSelect1H_18[21]};
  wire [3:0]  tryToRead_hi_lo_lo_21 = {tryToRead_hi_lo_lo_hi_21, tryToRead_hi_lo_lo_lo_21};
  wire [1:0]  tryToRead_hi_lo_hi_lo_21 = {inputSelect1H_21[21], inputSelect1H_20[21]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_21 = {inputSelect1H_23[21], inputSelect1H_22[21]};
  wire [3:0]  tryToRead_hi_lo_hi_21 = {tryToRead_hi_lo_hi_hi_21, tryToRead_hi_lo_hi_lo_21};
  wire [7:0]  tryToRead_hi_lo_21 = {tryToRead_hi_lo_hi_21, tryToRead_hi_lo_lo_21};
  wire [1:0]  tryToRead_hi_hi_lo_lo_21 = {inputSelect1H_25[21], inputSelect1H_24[21]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_21 = {inputSelect1H_27[21], inputSelect1H_26[21]};
  wire [3:0]  tryToRead_hi_hi_lo_21 = {tryToRead_hi_hi_lo_hi_21, tryToRead_hi_hi_lo_lo_21};
  wire [1:0]  tryToRead_hi_hi_hi_lo_21 = {inputSelect1H_29[21], inputSelect1H_28[21]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_21 = {inputSelect1H_31[21], inputSelect1H_30[21]};
  wire [3:0]  tryToRead_hi_hi_hi_21 = {tryToRead_hi_hi_hi_hi_21, tryToRead_hi_hi_hi_lo_21};
  wire [7:0]  tryToRead_hi_hi_21 = {tryToRead_hi_hi_hi_21, tryToRead_hi_hi_lo_21};
  wire [15:0] tryToRead_hi_21 = {tryToRead_hi_hi_21, tryToRead_hi_lo_21};
  wire [31:0] tryToRead_21 = {tryToRead_hi_21, tryToRead_lo_21};
  wire        output_21_valid_0 = |tryToRead_21;
  wire [4:0]  output_21_bits_vs_0 = selectReq_21_bits_vs;
  wire        output_21_bits_offset_0 = selectReq_21_bits_offset;
  wire [4:0]  output_21_bits_writeIndex_0 = selectReq_21_bits_requestIndex;
  wire [1:0]  output_21_bits_dataOffset_0 = selectReq_21_bits_dataOffset;
  assign selectReq_21_bits_dataOffset =
    (tryToRead_21[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_21[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_21[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_21[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_21[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_21[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_21[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_21[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_21[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_21[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_21[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_21[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_21[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_21[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_21[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_21[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_21[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_21[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_21[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_21[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_21[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_21[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_21[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_21[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_21[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_21[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_21_bits_requestIndex =
    {4'h0, tryToRead_21[1]} | {3'h0, tryToRead_21[2], 1'h0} | (tryToRead_21[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_21[4], 2'h0} | (tryToRead_21[5] ? 5'h5 : 5'h0) | (tryToRead_21[6] ? 5'h6 : 5'h0) | (tryToRead_21[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_21[8], 3'h0} | (tryToRead_21[9] ? 5'h9 : 5'h0) | (tryToRead_21[10] ? 5'hA : 5'h0) | (tryToRead_21[11] ? 5'hB : 5'h0) | (tryToRead_21[12] ? 5'hC : 5'h0) | (tryToRead_21[13] ? 5'hD : 5'h0)
    | (tryToRead_21[14] ? 5'hE : 5'h0) | (tryToRead_21[15] ? 5'hF : 5'h0) | {tryToRead_21[16], 4'h0} | (tryToRead_21[17] ? 5'h11 : 5'h0) | (tryToRead_21[18] ? 5'h12 : 5'h0) | (tryToRead_21[19] ? 5'h13 : 5'h0)
    | (tryToRead_21[20] ? 5'h14 : 5'h0) | (tryToRead_21[21] ? 5'h15 : 5'h0) | (tryToRead_21[22] ? 5'h16 : 5'h0) | (tryToRead_21[23] ? 5'h17 : 5'h0) | (tryToRead_21[24] ? 5'h18 : 5'h0) | (tryToRead_21[25] ? 5'h19 : 5'h0)
    | (tryToRead_21[26] ? 5'h1A : 5'h0) | (tryToRead_21[27] ? 5'h1B : 5'h0) | (tryToRead_21[28] ? 5'h1C : 5'h0) | (tryToRead_21[29] ? 5'h1D : 5'h0) | (tryToRead_21[30] ? 5'h1E : 5'h0) | {5{tryToRead_21[31]}};
  wire [4:0]  selectReq_21_bits_readLane =
    (tryToRead_21[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_21[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_21[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_21[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_21[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_21[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_21[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_21[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_21[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_21[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_21[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_21[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_21[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_21[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_21[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_21[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_21[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_21[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_21[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_21[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_21[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_21[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_21[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_21[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_21[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_21[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_21[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_21[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_21[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_21[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_21[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_21[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_21_bits_offset =
    tryToRead_21[0] & input_0_bits_offset_0 | tryToRead_21[1] & input_1_bits_offset_0 | tryToRead_21[2] & input_2_bits_offset_0 | tryToRead_21[3] & input_3_bits_offset_0 | tryToRead_21[4] & input_4_bits_offset_0 | tryToRead_21[5]
    & input_5_bits_offset_0 | tryToRead_21[6] & input_6_bits_offset_0 | tryToRead_21[7] & input_7_bits_offset_0 | tryToRead_21[8] & input_8_bits_offset_0 | tryToRead_21[9] & input_9_bits_offset_0 | tryToRead_21[10] & input_10_bits_offset_0
    | tryToRead_21[11] & input_11_bits_offset_0 | tryToRead_21[12] & input_12_bits_offset_0 | tryToRead_21[13] & input_13_bits_offset_0 | tryToRead_21[14] & input_14_bits_offset_0 | tryToRead_21[15] & input_15_bits_offset_0
    | tryToRead_21[16] & input_16_bits_offset_0 | tryToRead_21[17] & input_17_bits_offset_0 | tryToRead_21[18] & input_18_bits_offset_0 | tryToRead_21[19] & input_19_bits_offset_0 | tryToRead_21[20] & input_20_bits_offset_0
    | tryToRead_21[21] & input_21_bits_offset_0 | tryToRead_21[22] & input_22_bits_offset_0 | tryToRead_21[23] & input_23_bits_offset_0 | tryToRead_21[24] & input_24_bits_offset_0 | tryToRead_21[25] & input_25_bits_offset_0
    | tryToRead_21[26] & input_26_bits_offset_0 | tryToRead_21[27] & input_27_bits_offset_0 | tryToRead_21[28] & input_28_bits_offset_0 | tryToRead_21[29] & input_29_bits_offset_0 | tryToRead_21[30] & input_30_bits_offset_0
    | tryToRead_21[31] & input_31_bits_offset_0;
  assign selectReq_21_bits_vs =
    (tryToRead_21[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_21[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_21[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_21[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_21[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_21[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_21[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_21[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_21[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_21[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_21[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_21[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_21[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_21[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_21[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_21[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_21[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_21[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_21[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_21[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_21[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_21[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_21[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_21[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_21[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_21[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_21[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_21[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_21[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_21[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_21[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_21[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_21_valid =
    tryToRead_21[0] & input_0_valid_0 | tryToRead_21[1] & input_1_valid_0 | tryToRead_21[2] & input_2_valid_0 | tryToRead_21[3] & input_3_valid_0 | tryToRead_21[4] & input_4_valid_0 | tryToRead_21[5] & input_5_valid_0 | tryToRead_21[6]
    & input_6_valid_0 | tryToRead_21[7] & input_7_valid_0 | tryToRead_21[8] & input_8_valid_0 | tryToRead_21[9] & input_9_valid_0 | tryToRead_21[10] & input_10_valid_0 | tryToRead_21[11] & input_11_valid_0 | tryToRead_21[12]
    & input_12_valid_0 | tryToRead_21[13] & input_13_valid_0 | tryToRead_21[14] & input_14_valid_0 | tryToRead_21[15] & input_15_valid_0 | tryToRead_21[16] & input_16_valid_0 | tryToRead_21[17] & input_17_valid_0 | tryToRead_21[18]
    & input_18_valid_0 | tryToRead_21[19] & input_19_valid_0 | tryToRead_21[20] & input_20_valid_0 | tryToRead_21[21] & input_21_valid_0 | tryToRead_21[22] & input_22_valid_0 | tryToRead_21[23] & input_23_valid_0 | tryToRead_21[24]
    & input_24_valid_0 | tryToRead_21[25] & input_25_valid_0 | tryToRead_21[26] & input_26_valid_0 | tryToRead_21[27] & input_27_valid_0 | tryToRead_21[28] & input_28_valid_0 | tryToRead_21[29] & input_29_valid_0 | tryToRead_21[30]
    & input_30_valid_0 | tryToRead_21[31] & input_31_valid_0;
  wire        selectReq_21_ready =
    tryToRead_21[0] & input_0_ready_0 | tryToRead_21[1] & input_1_ready_0 | tryToRead_21[2] & input_2_ready_0 | tryToRead_21[3] & input_3_ready_0 | tryToRead_21[4] & input_4_ready_0 | tryToRead_21[5] & input_5_ready_0 | tryToRead_21[6]
    & input_6_ready_0 | tryToRead_21[7] & input_7_ready_0 | tryToRead_21[8] & input_8_ready_0 | tryToRead_21[9] & input_9_ready_0 | tryToRead_21[10] & input_10_ready_0 | tryToRead_21[11] & input_11_ready_0 | tryToRead_21[12]
    & input_12_ready_0 | tryToRead_21[13] & input_13_ready_0 | tryToRead_21[14] & input_14_ready_0 | tryToRead_21[15] & input_15_ready_0 | tryToRead_21[16] & input_16_ready_0 | tryToRead_21[17] & input_17_ready_0 | tryToRead_21[18]
    & input_18_ready_0 | tryToRead_21[19] & input_19_ready_0 | tryToRead_21[20] & input_20_ready_0 | tryToRead_21[21] & input_21_ready_0 | tryToRead_21[22] & input_22_ready_0 | tryToRead_21[23] & input_23_ready_0 | tryToRead_21[24]
    & input_24_ready_0 | tryToRead_21[25] & input_25_ready_0 | tryToRead_21[26] & input_26_ready_0 | tryToRead_21[27] & input_27_ready_0 | tryToRead_21[28] & input_28_ready_0 | tryToRead_21[29] & input_29_ready_0 | tryToRead_21[30]
    & input_30_ready_0 | tryToRead_21[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_22 = {inputSelect1H_1[22], inputSelect1H_0[22]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_22 = {inputSelect1H_3[22], inputSelect1H_2[22]};
  wire [3:0]  tryToRead_lo_lo_lo_22 = {tryToRead_lo_lo_lo_hi_22, tryToRead_lo_lo_lo_lo_22};
  wire [1:0]  tryToRead_lo_lo_hi_lo_22 = {inputSelect1H_5[22], inputSelect1H_4[22]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_22 = {inputSelect1H_7[22], inputSelect1H_6[22]};
  wire [3:0]  tryToRead_lo_lo_hi_22 = {tryToRead_lo_lo_hi_hi_22, tryToRead_lo_lo_hi_lo_22};
  wire [7:0]  tryToRead_lo_lo_22 = {tryToRead_lo_lo_hi_22, tryToRead_lo_lo_lo_22};
  wire [1:0]  tryToRead_lo_hi_lo_lo_22 = {inputSelect1H_9[22], inputSelect1H_8[22]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_22 = {inputSelect1H_11[22], inputSelect1H_10[22]};
  wire [3:0]  tryToRead_lo_hi_lo_22 = {tryToRead_lo_hi_lo_hi_22, tryToRead_lo_hi_lo_lo_22};
  wire [1:0]  tryToRead_lo_hi_hi_lo_22 = {inputSelect1H_13[22], inputSelect1H_12[22]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_22 = {inputSelect1H_15[22], inputSelect1H_14[22]};
  wire [3:0]  tryToRead_lo_hi_hi_22 = {tryToRead_lo_hi_hi_hi_22, tryToRead_lo_hi_hi_lo_22};
  wire [7:0]  tryToRead_lo_hi_22 = {tryToRead_lo_hi_hi_22, tryToRead_lo_hi_lo_22};
  wire [15:0] tryToRead_lo_22 = {tryToRead_lo_hi_22, tryToRead_lo_lo_22};
  wire [1:0]  tryToRead_hi_lo_lo_lo_22 = {inputSelect1H_17[22], inputSelect1H_16[22]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_22 = {inputSelect1H_19[22], inputSelect1H_18[22]};
  wire [3:0]  tryToRead_hi_lo_lo_22 = {tryToRead_hi_lo_lo_hi_22, tryToRead_hi_lo_lo_lo_22};
  wire [1:0]  tryToRead_hi_lo_hi_lo_22 = {inputSelect1H_21[22], inputSelect1H_20[22]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_22 = {inputSelect1H_23[22], inputSelect1H_22[22]};
  wire [3:0]  tryToRead_hi_lo_hi_22 = {tryToRead_hi_lo_hi_hi_22, tryToRead_hi_lo_hi_lo_22};
  wire [7:0]  tryToRead_hi_lo_22 = {tryToRead_hi_lo_hi_22, tryToRead_hi_lo_lo_22};
  wire [1:0]  tryToRead_hi_hi_lo_lo_22 = {inputSelect1H_25[22], inputSelect1H_24[22]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_22 = {inputSelect1H_27[22], inputSelect1H_26[22]};
  wire [3:0]  tryToRead_hi_hi_lo_22 = {tryToRead_hi_hi_lo_hi_22, tryToRead_hi_hi_lo_lo_22};
  wire [1:0]  tryToRead_hi_hi_hi_lo_22 = {inputSelect1H_29[22], inputSelect1H_28[22]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_22 = {inputSelect1H_31[22], inputSelect1H_30[22]};
  wire [3:0]  tryToRead_hi_hi_hi_22 = {tryToRead_hi_hi_hi_hi_22, tryToRead_hi_hi_hi_lo_22};
  wire [7:0]  tryToRead_hi_hi_22 = {tryToRead_hi_hi_hi_22, tryToRead_hi_hi_lo_22};
  wire [15:0] tryToRead_hi_22 = {tryToRead_hi_hi_22, tryToRead_hi_lo_22};
  wire [31:0] tryToRead_22 = {tryToRead_hi_22, tryToRead_lo_22};
  wire        output_22_valid_0 = |tryToRead_22;
  wire [4:0]  output_22_bits_vs_0 = selectReq_22_bits_vs;
  wire        output_22_bits_offset_0 = selectReq_22_bits_offset;
  wire [4:0]  output_22_bits_writeIndex_0 = selectReq_22_bits_requestIndex;
  wire [1:0]  output_22_bits_dataOffset_0 = selectReq_22_bits_dataOffset;
  assign selectReq_22_bits_dataOffset =
    (tryToRead_22[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_22[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_22[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_22[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_22[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_22[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_22[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_22[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_22[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_22[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_22[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_22[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_22[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_22[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_22[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_22[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_22[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_22[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_22[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_22[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_22[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_22[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_22[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_22[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_22[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_22[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_22_bits_requestIndex =
    {4'h0, tryToRead_22[1]} | {3'h0, tryToRead_22[2], 1'h0} | (tryToRead_22[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_22[4], 2'h0} | (tryToRead_22[5] ? 5'h5 : 5'h0) | (tryToRead_22[6] ? 5'h6 : 5'h0) | (tryToRead_22[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_22[8], 3'h0} | (tryToRead_22[9] ? 5'h9 : 5'h0) | (tryToRead_22[10] ? 5'hA : 5'h0) | (tryToRead_22[11] ? 5'hB : 5'h0) | (tryToRead_22[12] ? 5'hC : 5'h0) | (tryToRead_22[13] ? 5'hD : 5'h0)
    | (tryToRead_22[14] ? 5'hE : 5'h0) | (tryToRead_22[15] ? 5'hF : 5'h0) | {tryToRead_22[16], 4'h0} | (tryToRead_22[17] ? 5'h11 : 5'h0) | (tryToRead_22[18] ? 5'h12 : 5'h0) | (tryToRead_22[19] ? 5'h13 : 5'h0)
    | (tryToRead_22[20] ? 5'h14 : 5'h0) | (tryToRead_22[21] ? 5'h15 : 5'h0) | (tryToRead_22[22] ? 5'h16 : 5'h0) | (tryToRead_22[23] ? 5'h17 : 5'h0) | (tryToRead_22[24] ? 5'h18 : 5'h0) | (tryToRead_22[25] ? 5'h19 : 5'h0)
    | (tryToRead_22[26] ? 5'h1A : 5'h0) | (tryToRead_22[27] ? 5'h1B : 5'h0) | (tryToRead_22[28] ? 5'h1C : 5'h0) | (tryToRead_22[29] ? 5'h1D : 5'h0) | (tryToRead_22[30] ? 5'h1E : 5'h0) | {5{tryToRead_22[31]}};
  wire [4:0]  selectReq_22_bits_readLane =
    (tryToRead_22[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_22[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_22[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_22[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_22[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_22[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_22[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_22[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_22[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_22[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_22[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_22[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_22[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_22[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_22[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_22[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_22[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_22[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_22[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_22[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_22[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_22[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_22[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_22[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_22[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_22[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_22[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_22[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_22[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_22[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_22[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_22[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_22_bits_offset =
    tryToRead_22[0] & input_0_bits_offset_0 | tryToRead_22[1] & input_1_bits_offset_0 | tryToRead_22[2] & input_2_bits_offset_0 | tryToRead_22[3] & input_3_bits_offset_0 | tryToRead_22[4] & input_4_bits_offset_0 | tryToRead_22[5]
    & input_5_bits_offset_0 | tryToRead_22[6] & input_6_bits_offset_0 | tryToRead_22[7] & input_7_bits_offset_0 | tryToRead_22[8] & input_8_bits_offset_0 | tryToRead_22[9] & input_9_bits_offset_0 | tryToRead_22[10] & input_10_bits_offset_0
    | tryToRead_22[11] & input_11_bits_offset_0 | tryToRead_22[12] & input_12_bits_offset_0 | tryToRead_22[13] & input_13_bits_offset_0 | tryToRead_22[14] & input_14_bits_offset_0 | tryToRead_22[15] & input_15_bits_offset_0
    | tryToRead_22[16] & input_16_bits_offset_0 | tryToRead_22[17] & input_17_bits_offset_0 | tryToRead_22[18] & input_18_bits_offset_0 | tryToRead_22[19] & input_19_bits_offset_0 | tryToRead_22[20] & input_20_bits_offset_0
    | tryToRead_22[21] & input_21_bits_offset_0 | tryToRead_22[22] & input_22_bits_offset_0 | tryToRead_22[23] & input_23_bits_offset_0 | tryToRead_22[24] & input_24_bits_offset_0 | tryToRead_22[25] & input_25_bits_offset_0
    | tryToRead_22[26] & input_26_bits_offset_0 | tryToRead_22[27] & input_27_bits_offset_0 | tryToRead_22[28] & input_28_bits_offset_0 | tryToRead_22[29] & input_29_bits_offset_0 | tryToRead_22[30] & input_30_bits_offset_0
    | tryToRead_22[31] & input_31_bits_offset_0;
  assign selectReq_22_bits_vs =
    (tryToRead_22[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_22[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_22[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_22[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_22[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_22[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_22[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_22[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_22[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_22[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_22[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_22[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_22[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_22[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_22[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_22[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_22[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_22[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_22[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_22[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_22[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_22[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_22[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_22[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_22[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_22[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_22[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_22[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_22[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_22[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_22[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_22[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_22_valid =
    tryToRead_22[0] & input_0_valid_0 | tryToRead_22[1] & input_1_valid_0 | tryToRead_22[2] & input_2_valid_0 | tryToRead_22[3] & input_3_valid_0 | tryToRead_22[4] & input_4_valid_0 | tryToRead_22[5] & input_5_valid_0 | tryToRead_22[6]
    & input_6_valid_0 | tryToRead_22[7] & input_7_valid_0 | tryToRead_22[8] & input_8_valid_0 | tryToRead_22[9] & input_9_valid_0 | tryToRead_22[10] & input_10_valid_0 | tryToRead_22[11] & input_11_valid_0 | tryToRead_22[12]
    & input_12_valid_0 | tryToRead_22[13] & input_13_valid_0 | tryToRead_22[14] & input_14_valid_0 | tryToRead_22[15] & input_15_valid_0 | tryToRead_22[16] & input_16_valid_0 | tryToRead_22[17] & input_17_valid_0 | tryToRead_22[18]
    & input_18_valid_0 | tryToRead_22[19] & input_19_valid_0 | tryToRead_22[20] & input_20_valid_0 | tryToRead_22[21] & input_21_valid_0 | tryToRead_22[22] & input_22_valid_0 | tryToRead_22[23] & input_23_valid_0 | tryToRead_22[24]
    & input_24_valid_0 | tryToRead_22[25] & input_25_valid_0 | tryToRead_22[26] & input_26_valid_0 | tryToRead_22[27] & input_27_valid_0 | tryToRead_22[28] & input_28_valid_0 | tryToRead_22[29] & input_29_valid_0 | tryToRead_22[30]
    & input_30_valid_0 | tryToRead_22[31] & input_31_valid_0;
  wire        selectReq_22_ready =
    tryToRead_22[0] & input_0_ready_0 | tryToRead_22[1] & input_1_ready_0 | tryToRead_22[2] & input_2_ready_0 | tryToRead_22[3] & input_3_ready_0 | tryToRead_22[4] & input_4_ready_0 | tryToRead_22[5] & input_5_ready_0 | tryToRead_22[6]
    & input_6_ready_0 | tryToRead_22[7] & input_7_ready_0 | tryToRead_22[8] & input_8_ready_0 | tryToRead_22[9] & input_9_ready_0 | tryToRead_22[10] & input_10_ready_0 | tryToRead_22[11] & input_11_ready_0 | tryToRead_22[12]
    & input_12_ready_0 | tryToRead_22[13] & input_13_ready_0 | tryToRead_22[14] & input_14_ready_0 | tryToRead_22[15] & input_15_ready_0 | tryToRead_22[16] & input_16_ready_0 | tryToRead_22[17] & input_17_ready_0 | tryToRead_22[18]
    & input_18_ready_0 | tryToRead_22[19] & input_19_ready_0 | tryToRead_22[20] & input_20_ready_0 | tryToRead_22[21] & input_21_ready_0 | tryToRead_22[22] & input_22_ready_0 | tryToRead_22[23] & input_23_ready_0 | tryToRead_22[24]
    & input_24_ready_0 | tryToRead_22[25] & input_25_ready_0 | tryToRead_22[26] & input_26_ready_0 | tryToRead_22[27] & input_27_ready_0 | tryToRead_22[28] & input_28_ready_0 | tryToRead_22[29] & input_29_ready_0 | tryToRead_22[30]
    & input_30_ready_0 | tryToRead_22[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_23 = {inputSelect1H_1[23], inputSelect1H_0[23]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_23 = {inputSelect1H_3[23], inputSelect1H_2[23]};
  wire [3:0]  tryToRead_lo_lo_lo_23 = {tryToRead_lo_lo_lo_hi_23, tryToRead_lo_lo_lo_lo_23};
  wire [1:0]  tryToRead_lo_lo_hi_lo_23 = {inputSelect1H_5[23], inputSelect1H_4[23]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_23 = {inputSelect1H_7[23], inputSelect1H_6[23]};
  wire [3:0]  tryToRead_lo_lo_hi_23 = {tryToRead_lo_lo_hi_hi_23, tryToRead_lo_lo_hi_lo_23};
  wire [7:0]  tryToRead_lo_lo_23 = {tryToRead_lo_lo_hi_23, tryToRead_lo_lo_lo_23};
  wire [1:0]  tryToRead_lo_hi_lo_lo_23 = {inputSelect1H_9[23], inputSelect1H_8[23]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_23 = {inputSelect1H_11[23], inputSelect1H_10[23]};
  wire [3:0]  tryToRead_lo_hi_lo_23 = {tryToRead_lo_hi_lo_hi_23, tryToRead_lo_hi_lo_lo_23};
  wire [1:0]  tryToRead_lo_hi_hi_lo_23 = {inputSelect1H_13[23], inputSelect1H_12[23]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_23 = {inputSelect1H_15[23], inputSelect1H_14[23]};
  wire [3:0]  tryToRead_lo_hi_hi_23 = {tryToRead_lo_hi_hi_hi_23, tryToRead_lo_hi_hi_lo_23};
  wire [7:0]  tryToRead_lo_hi_23 = {tryToRead_lo_hi_hi_23, tryToRead_lo_hi_lo_23};
  wire [15:0] tryToRead_lo_23 = {tryToRead_lo_hi_23, tryToRead_lo_lo_23};
  wire [1:0]  tryToRead_hi_lo_lo_lo_23 = {inputSelect1H_17[23], inputSelect1H_16[23]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_23 = {inputSelect1H_19[23], inputSelect1H_18[23]};
  wire [3:0]  tryToRead_hi_lo_lo_23 = {tryToRead_hi_lo_lo_hi_23, tryToRead_hi_lo_lo_lo_23};
  wire [1:0]  tryToRead_hi_lo_hi_lo_23 = {inputSelect1H_21[23], inputSelect1H_20[23]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_23 = {inputSelect1H_23[23], inputSelect1H_22[23]};
  wire [3:0]  tryToRead_hi_lo_hi_23 = {tryToRead_hi_lo_hi_hi_23, tryToRead_hi_lo_hi_lo_23};
  wire [7:0]  tryToRead_hi_lo_23 = {tryToRead_hi_lo_hi_23, tryToRead_hi_lo_lo_23};
  wire [1:0]  tryToRead_hi_hi_lo_lo_23 = {inputSelect1H_25[23], inputSelect1H_24[23]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_23 = {inputSelect1H_27[23], inputSelect1H_26[23]};
  wire [3:0]  tryToRead_hi_hi_lo_23 = {tryToRead_hi_hi_lo_hi_23, tryToRead_hi_hi_lo_lo_23};
  wire [1:0]  tryToRead_hi_hi_hi_lo_23 = {inputSelect1H_29[23], inputSelect1H_28[23]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_23 = {inputSelect1H_31[23], inputSelect1H_30[23]};
  wire [3:0]  tryToRead_hi_hi_hi_23 = {tryToRead_hi_hi_hi_hi_23, tryToRead_hi_hi_hi_lo_23};
  wire [7:0]  tryToRead_hi_hi_23 = {tryToRead_hi_hi_hi_23, tryToRead_hi_hi_lo_23};
  wire [15:0] tryToRead_hi_23 = {tryToRead_hi_hi_23, tryToRead_hi_lo_23};
  wire [31:0] tryToRead_23 = {tryToRead_hi_23, tryToRead_lo_23};
  wire        output_23_valid_0 = |tryToRead_23;
  wire [4:0]  output_23_bits_vs_0 = selectReq_23_bits_vs;
  wire        output_23_bits_offset_0 = selectReq_23_bits_offset;
  wire [4:0]  output_23_bits_writeIndex_0 = selectReq_23_bits_requestIndex;
  wire [1:0]  output_23_bits_dataOffset_0 = selectReq_23_bits_dataOffset;
  assign selectReq_23_bits_dataOffset =
    (tryToRead_23[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_23[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_23[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_23[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_23[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_23[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_23[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_23[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_23[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_23[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_23[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_23[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_23[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_23[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_23[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_23[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_23[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_23[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_23[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_23[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_23[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_23[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_23[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_23[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_23[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_23[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_23_bits_requestIndex =
    {4'h0, tryToRead_23[1]} | {3'h0, tryToRead_23[2], 1'h0} | (tryToRead_23[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_23[4], 2'h0} | (tryToRead_23[5] ? 5'h5 : 5'h0) | (tryToRead_23[6] ? 5'h6 : 5'h0) | (tryToRead_23[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_23[8], 3'h0} | (tryToRead_23[9] ? 5'h9 : 5'h0) | (tryToRead_23[10] ? 5'hA : 5'h0) | (tryToRead_23[11] ? 5'hB : 5'h0) | (tryToRead_23[12] ? 5'hC : 5'h0) | (tryToRead_23[13] ? 5'hD : 5'h0)
    | (tryToRead_23[14] ? 5'hE : 5'h0) | (tryToRead_23[15] ? 5'hF : 5'h0) | {tryToRead_23[16], 4'h0} | (tryToRead_23[17] ? 5'h11 : 5'h0) | (tryToRead_23[18] ? 5'h12 : 5'h0) | (tryToRead_23[19] ? 5'h13 : 5'h0)
    | (tryToRead_23[20] ? 5'h14 : 5'h0) | (tryToRead_23[21] ? 5'h15 : 5'h0) | (tryToRead_23[22] ? 5'h16 : 5'h0) | (tryToRead_23[23] ? 5'h17 : 5'h0) | (tryToRead_23[24] ? 5'h18 : 5'h0) | (tryToRead_23[25] ? 5'h19 : 5'h0)
    | (tryToRead_23[26] ? 5'h1A : 5'h0) | (tryToRead_23[27] ? 5'h1B : 5'h0) | (tryToRead_23[28] ? 5'h1C : 5'h0) | (tryToRead_23[29] ? 5'h1D : 5'h0) | (tryToRead_23[30] ? 5'h1E : 5'h0) | {5{tryToRead_23[31]}};
  wire [4:0]  selectReq_23_bits_readLane =
    (tryToRead_23[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_23[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_23[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_23[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_23[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_23[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_23[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_23[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_23[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_23[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_23[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_23[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_23[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_23[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_23[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_23[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_23[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_23[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_23[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_23[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_23[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_23[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_23[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_23[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_23[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_23[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_23[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_23[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_23[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_23[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_23[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_23[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_23_bits_offset =
    tryToRead_23[0] & input_0_bits_offset_0 | tryToRead_23[1] & input_1_bits_offset_0 | tryToRead_23[2] & input_2_bits_offset_0 | tryToRead_23[3] & input_3_bits_offset_0 | tryToRead_23[4] & input_4_bits_offset_0 | tryToRead_23[5]
    & input_5_bits_offset_0 | tryToRead_23[6] & input_6_bits_offset_0 | tryToRead_23[7] & input_7_bits_offset_0 | tryToRead_23[8] & input_8_bits_offset_0 | tryToRead_23[9] & input_9_bits_offset_0 | tryToRead_23[10] & input_10_bits_offset_0
    | tryToRead_23[11] & input_11_bits_offset_0 | tryToRead_23[12] & input_12_bits_offset_0 | tryToRead_23[13] & input_13_bits_offset_0 | tryToRead_23[14] & input_14_bits_offset_0 | tryToRead_23[15] & input_15_bits_offset_0
    | tryToRead_23[16] & input_16_bits_offset_0 | tryToRead_23[17] & input_17_bits_offset_0 | tryToRead_23[18] & input_18_bits_offset_0 | tryToRead_23[19] & input_19_bits_offset_0 | tryToRead_23[20] & input_20_bits_offset_0
    | tryToRead_23[21] & input_21_bits_offset_0 | tryToRead_23[22] & input_22_bits_offset_0 | tryToRead_23[23] & input_23_bits_offset_0 | tryToRead_23[24] & input_24_bits_offset_0 | tryToRead_23[25] & input_25_bits_offset_0
    | tryToRead_23[26] & input_26_bits_offset_0 | tryToRead_23[27] & input_27_bits_offset_0 | tryToRead_23[28] & input_28_bits_offset_0 | tryToRead_23[29] & input_29_bits_offset_0 | tryToRead_23[30] & input_30_bits_offset_0
    | tryToRead_23[31] & input_31_bits_offset_0;
  assign selectReq_23_bits_vs =
    (tryToRead_23[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_23[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_23[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_23[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_23[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_23[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_23[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_23[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_23[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_23[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_23[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_23[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_23[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_23[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_23[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_23[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_23[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_23[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_23[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_23[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_23[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_23[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_23[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_23[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_23[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_23[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_23[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_23[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_23[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_23[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_23[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_23[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_23_valid =
    tryToRead_23[0] & input_0_valid_0 | tryToRead_23[1] & input_1_valid_0 | tryToRead_23[2] & input_2_valid_0 | tryToRead_23[3] & input_3_valid_0 | tryToRead_23[4] & input_4_valid_0 | tryToRead_23[5] & input_5_valid_0 | tryToRead_23[6]
    & input_6_valid_0 | tryToRead_23[7] & input_7_valid_0 | tryToRead_23[8] & input_8_valid_0 | tryToRead_23[9] & input_9_valid_0 | tryToRead_23[10] & input_10_valid_0 | tryToRead_23[11] & input_11_valid_0 | tryToRead_23[12]
    & input_12_valid_0 | tryToRead_23[13] & input_13_valid_0 | tryToRead_23[14] & input_14_valid_0 | tryToRead_23[15] & input_15_valid_0 | tryToRead_23[16] & input_16_valid_0 | tryToRead_23[17] & input_17_valid_0 | tryToRead_23[18]
    & input_18_valid_0 | tryToRead_23[19] & input_19_valid_0 | tryToRead_23[20] & input_20_valid_0 | tryToRead_23[21] & input_21_valid_0 | tryToRead_23[22] & input_22_valid_0 | tryToRead_23[23] & input_23_valid_0 | tryToRead_23[24]
    & input_24_valid_0 | tryToRead_23[25] & input_25_valid_0 | tryToRead_23[26] & input_26_valid_0 | tryToRead_23[27] & input_27_valid_0 | tryToRead_23[28] & input_28_valid_0 | tryToRead_23[29] & input_29_valid_0 | tryToRead_23[30]
    & input_30_valid_0 | tryToRead_23[31] & input_31_valid_0;
  wire        selectReq_23_ready =
    tryToRead_23[0] & input_0_ready_0 | tryToRead_23[1] & input_1_ready_0 | tryToRead_23[2] & input_2_ready_0 | tryToRead_23[3] & input_3_ready_0 | tryToRead_23[4] & input_4_ready_0 | tryToRead_23[5] & input_5_ready_0 | tryToRead_23[6]
    & input_6_ready_0 | tryToRead_23[7] & input_7_ready_0 | tryToRead_23[8] & input_8_ready_0 | tryToRead_23[9] & input_9_ready_0 | tryToRead_23[10] & input_10_ready_0 | tryToRead_23[11] & input_11_ready_0 | tryToRead_23[12]
    & input_12_ready_0 | tryToRead_23[13] & input_13_ready_0 | tryToRead_23[14] & input_14_ready_0 | tryToRead_23[15] & input_15_ready_0 | tryToRead_23[16] & input_16_ready_0 | tryToRead_23[17] & input_17_ready_0 | tryToRead_23[18]
    & input_18_ready_0 | tryToRead_23[19] & input_19_ready_0 | tryToRead_23[20] & input_20_ready_0 | tryToRead_23[21] & input_21_ready_0 | tryToRead_23[22] & input_22_ready_0 | tryToRead_23[23] & input_23_ready_0 | tryToRead_23[24]
    & input_24_ready_0 | tryToRead_23[25] & input_25_ready_0 | tryToRead_23[26] & input_26_ready_0 | tryToRead_23[27] & input_27_ready_0 | tryToRead_23[28] & input_28_ready_0 | tryToRead_23[29] & input_29_ready_0 | tryToRead_23[30]
    & input_30_ready_0 | tryToRead_23[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_24 = {inputSelect1H_1[24], inputSelect1H_0[24]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_24 = {inputSelect1H_3[24], inputSelect1H_2[24]};
  wire [3:0]  tryToRead_lo_lo_lo_24 = {tryToRead_lo_lo_lo_hi_24, tryToRead_lo_lo_lo_lo_24};
  wire [1:0]  tryToRead_lo_lo_hi_lo_24 = {inputSelect1H_5[24], inputSelect1H_4[24]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_24 = {inputSelect1H_7[24], inputSelect1H_6[24]};
  wire [3:0]  tryToRead_lo_lo_hi_24 = {tryToRead_lo_lo_hi_hi_24, tryToRead_lo_lo_hi_lo_24};
  wire [7:0]  tryToRead_lo_lo_24 = {tryToRead_lo_lo_hi_24, tryToRead_lo_lo_lo_24};
  wire [1:0]  tryToRead_lo_hi_lo_lo_24 = {inputSelect1H_9[24], inputSelect1H_8[24]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_24 = {inputSelect1H_11[24], inputSelect1H_10[24]};
  wire [3:0]  tryToRead_lo_hi_lo_24 = {tryToRead_lo_hi_lo_hi_24, tryToRead_lo_hi_lo_lo_24};
  wire [1:0]  tryToRead_lo_hi_hi_lo_24 = {inputSelect1H_13[24], inputSelect1H_12[24]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_24 = {inputSelect1H_15[24], inputSelect1H_14[24]};
  wire [3:0]  tryToRead_lo_hi_hi_24 = {tryToRead_lo_hi_hi_hi_24, tryToRead_lo_hi_hi_lo_24};
  wire [7:0]  tryToRead_lo_hi_24 = {tryToRead_lo_hi_hi_24, tryToRead_lo_hi_lo_24};
  wire [15:0] tryToRead_lo_24 = {tryToRead_lo_hi_24, tryToRead_lo_lo_24};
  wire [1:0]  tryToRead_hi_lo_lo_lo_24 = {inputSelect1H_17[24], inputSelect1H_16[24]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_24 = {inputSelect1H_19[24], inputSelect1H_18[24]};
  wire [3:0]  tryToRead_hi_lo_lo_24 = {tryToRead_hi_lo_lo_hi_24, tryToRead_hi_lo_lo_lo_24};
  wire [1:0]  tryToRead_hi_lo_hi_lo_24 = {inputSelect1H_21[24], inputSelect1H_20[24]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_24 = {inputSelect1H_23[24], inputSelect1H_22[24]};
  wire [3:0]  tryToRead_hi_lo_hi_24 = {tryToRead_hi_lo_hi_hi_24, tryToRead_hi_lo_hi_lo_24};
  wire [7:0]  tryToRead_hi_lo_24 = {tryToRead_hi_lo_hi_24, tryToRead_hi_lo_lo_24};
  wire [1:0]  tryToRead_hi_hi_lo_lo_24 = {inputSelect1H_25[24], inputSelect1H_24[24]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_24 = {inputSelect1H_27[24], inputSelect1H_26[24]};
  wire [3:0]  tryToRead_hi_hi_lo_24 = {tryToRead_hi_hi_lo_hi_24, tryToRead_hi_hi_lo_lo_24};
  wire [1:0]  tryToRead_hi_hi_hi_lo_24 = {inputSelect1H_29[24], inputSelect1H_28[24]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_24 = {inputSelect1H_31[24], inputSelect1H_30[24]};
  wire [3:0]  tryToRead_hi_hi_hi_24 = {tryToRead_hi_hi_hi_hi_24, tryToRead_hi_hi_hi_lo_24};
  wire [7:0]  tryToRead_hi_hi_24 = {tryToRead_hi_hi_hi_24, tryToRead_hi_hi_lo_24};
  wire [15:0] tryToRead_hi_24 = {tryToRead_hi_hi_24, tryToRead_hi_lo_24};
  wire [31:0] tryToRead_24 = {tryToRead_hi_24, tryToRead_lo_24};
  wire        output_24_valid_0 = |tryToRead_24;
  wire [4:0]  output_24_bits_vs_0 = selectReq_24_bits_vs;
  wire        output_24_bits_offset_0 = selectReq_24_bits_offset;
  wire [4:0]  output_24_bits_writeIndex_0 = selectReq_24_bits_requestIndex;
  wire [1:0]  output_24_bits_dataOffset_0 = selectReq_24_bits_dataOffset;
  assign selectReq_24_bits_dataOffset =
    (tryToRead_24[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_24[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_24[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_24[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_24[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_24[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_24[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_24[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_24[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_24[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_24[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_24[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_24[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_24[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_24[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_24[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_24[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_24[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_24[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_24[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_24[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_24[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_24[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_24[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_24[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_24[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_24_bits_requestIndex =
    {4'h0, tryToRead_24[1]} | {3'h0, tryToRead_24[2], 1'h0} | (tryToRead_24[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_24[4], 2'h0} | (tryToRead_24[5] ? 5'h5 : 5'h0) | (tryToRead_24[6] ? 5'h6 : 5'h0) | (tryToRead_24[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_24[8], 3'h0} | (tryToRead_24[9] ? 5'h9 : 5'h0) | (tryToRead_24[10] ? 5'hA : 5'h0) | (tryToRead_24[11] ? 5'hB : 5'h0) | (tryToRead_24[12] ? 5'hC : 5'h0) | (tryToRead_24[13] ? 5'hD : 5'h0)
    | (tryToRead_24[14] ? 5'hE : 5'h0) | (tryToRead_24[15] ? 5'hF : 5'h0) | {tryToRead_24[16], 4'h0} | (tryToRead_24[17] ? 5'h11 : 5'h0) | (tryToRead_24[18] ? 5'h12 : 5'h0) | (tryToRead_24[19] ? 5'h13 : 5'h0)
    | (tryToRead_24[20] ? 5'h14 : 5'h0) | (tryToRead_24[21] ? 5'h15 : 5'h0) | (tryToRead_24[22] ? 5'h16 : 5'h0) | (tryToRead_24[23] ? 5'h17 : 5'h0) | (tryToRead_24[24] ? 5'h18 : 5'h0) | (tryToRead_24[25] ? 5'h19 : 5'h0)
    | (tryToRead_24[26] ? 5'h1A : 5'h0) | (tryToRead_24[27] ? 5'h1B : 5'h0) | (tryToRead_24[28] ? 5'h1C : 5'h0) | (tryToRead_24[29] ? 5'h1D : 5'h0) | (tryToRead_24[30] ? 5'h1E : 5'h0) | {5{tryToRead_24[31]}};
  wire [4:0]  selectReq_24_bits_readLane =
    (tryToRead_24[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_24[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_24[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_24[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_24[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_24[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_24[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_24[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_24[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_24[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_24[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_24[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_24[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_24[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_24[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_24[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_24[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_24[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_24[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_24[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_24[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_24[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_24[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_24[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_24[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_24[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_24[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_24[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_24[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_24[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_24[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_24[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_24_bits_offset =
    tryToRead_24[0] & input_0_bits_offset_0 | tryToRead_24[1] & input_1_bits_offset_0 | tryToRead_24[2] & input_2_bits_offset_0 | tryToRead_24[3] & input_3_bits_offset_0 | tryToRead_24[4] & input_4_bits_offset_0 | tryToRead_24[5]
    & input_5_bits_offset_0 | tryToRead_24[6] & input_6_bits_offset_0 | tryToRead_24[7] & input_7_bits_offset_0 | tryToRead_24[8] & input_8_bits_offset_0 | tryToRead_24[9] & input_9_bits_offset_0 | tryToRead_24[10] & input_10_bits_offset_0
    | tryToRead_24[11] & input_11_bits_offset_0 | tryToRead_24[12] & input_12_bits_offset_0 | tryToRead_24[13] & input_13_bits_offset_0 | tryToRead_24[14] & input_14_bits_offset_0 | tryToRead_24[15] & input_15_bits_offset_0
    | tryToRead_24[16] & input_16_bits_offset_0 | tryToRead_24[17] & input_17_bits_offset_0 | tryToRead_24[18] & input_18_bits_offset_0 | tryToRead_24[19] & input_19_bits_offset_0 | tryToRead_24[20] & input_20_bits_offset_0
    | tryToRead_24[21] & input_21_bits_offset_0 | tryToRead_24[22] & input_22_bits_offset_0 | tryToRead_24[23] & input_23_bits_offset_0 | tryToRead_24[24] & input_24_bits_offset_0 | tryToRead_24[25] & input_25_bits_offset_0
    | tryToRead_24[26] & input_26_bits_offset_0 | tryToRead_24[27] & input_27_bits_offset_0 | tryToRead_24[28] & input_28_bits_offset_0 | tryToRead_24[29] & input_29_bits_offset_0 | tryToRead_24[30] & input_30_bits_offset_0
    | tryToRead_24[31] & input_31_bits_offset_0;
  assign selectReq_24_bits_vs =
    (tryToRead_24[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_24[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_24[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_24[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_24[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_24[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_24[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_24[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_24[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_24[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_24[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_24[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_24[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_24[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_24[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_24[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_24[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_24[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_24[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_24[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_24[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_24[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_24[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_24[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_24[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_24[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_24[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_24[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_24[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_24[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_24[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_24[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_24_valid =
    tryToRead_24[0] & input_0_valid_0 | tryToRead_24[1] & input_1_valid_0 | tryToRead_24[2] & input_2_valid_0 | tryToRead_24[3] & input_3_valid_0 | tryToRead_24[4] & input_4_valid_0 | tryToRead_24[5] & input_5_valid_0 | tryToRead_24[6]
    & input_6_valid_0 | tryToRead_24[7] & input_7_valid_0 | tryToRead_24[8] & input_8_valid_0 | tryToRead_24[9] & input_9_valid_0 | tryToRead_24[10] & input_10_valid_0 | tryToRead_24[11] & input_11_valid_0 | tryToRead_24[12]
    & input_12_valid_0 | tryToRead_24[13] & input_13_valid_0 | tryToRead_24[14] & input_14_valid_0 | tryToRead_24[15] & input_15_valid_0 | tryToRead_24[16] & input_16_valid_0 | tryToRead_24[17] & input_17_valid_0 | tryToRead_24[18]
    & input_18_valid_0 | tryToRead_24[19] & input_19_valid_0 | tryToRead_24[20] & input_20_valid_0 | tryToRead_24[21] & input_21_valid_0 | tryToRead_24[22] & input_22_valid_0 | tryToRead_24[23] & input_23_valid_0 | tryToRead_24[24]
    & input_24_valid_0 | tryToRead_24[25] & input_25_valid_0 | tryToRead_24[26] & input_26_valid_0 | tryToRead_24[27] & input_27_valid_0 | tryToRead_24[28] & input_28_valid_0 | tryToRead_24[29] & input_29_valid_0 | tryToRead_24[30]
    & input_30_valid_0 | tryToRead_24[31] & input_31_valid_0;
  wire        selectReq_24_ready =
    tryToRead_24[0] & input_0_ready_0 | tryToRead_24[1] & input_1_ready_0 | tryToRead_24[2] & input_2_ready_0 | tryToRead_24[3] & input_3_ready_0 | tryToRead_24[4] & input_4_ready_0 | tryToRead_24[5] & input_5_ready_0 | tryToRead_24[6]
    & input_6_ready_0 | tryToRead_24[7] & input_7_ready_0 | tryToRead_24[8] & input_8_ready_0 | tryToRead_24[9] & input_9_ready_0 | tryToRead_24[10] & input_10_ready_0 | tryToRead_24[11] & input_11_ready_0 | tryToRead_24[12]
    & input_12_ready_0 | tryToRead_24[13] & input_13_ready_0 | tryToRead_24[14] & input_14_ready_0 | tryToRead_24[15] & input_15_ready_0 | tryToRead_24[16] & input_16_ready_0 | tryToRead_24[17] & input_17_ready_0 | tryToRead_24[18]
    & input_18_ready_0 | tryToRead_24[19] & input_19_ready_0 | tryToRead_24[20] & input_20_ready_0 | tryToRead_24[21] & input_21_ready_0 | tryToRead_24[22] & input_22_ready_0 | tryToRead_24[23] & input_23_ready_0 | tryToRead_24[24]
    & input_24_ready_0 | tryToRead_24[25] & input_25_ready_0 | tryToRead_24[26] & input_26_ready_0 | tryToRead_24[27] & input_27_ready_0 | tryToRead_24[28] & input_28_ready_0 | tryToRead_24[29] & input_29_ready_0 | tryToRead_24[30]
    & input_30_ready_0 | tryToRead_24[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_25 = {inputSelect1H_1[25], inputSelect1H_0[25]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_25 = {inputSelect1H_3[25], inputSelect1H_2[25]};
  wire [3:0]  tryToRead_lo_lo_lo_25 = {tryToRead_lo_lo_lo_hi_25, tryToRead_lo_lo_lo_lo_25};
  wire [1:0]  tryToRead_lo_lo_hi_lo_25 = {inputSelect1H_5[25], inputSelect1H_4[25]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_25 = {inputSelect1H_7[25], inputSelect1H_6[25]};
  wire [3:0]  tryToRead_lo_lo_hi_25 = {tryToRead_lo_lo_hi_hi_25, tryToRead_lo_lo_hi_lo_25};
  wire [7:0]  tryToRead_lo_lo_25 = {tryToRead_lo_lo_hi_25, tryToRead_lo_lo_lo_25};
  wire [1:0]  tryToRead_lo_hi_lo_lo_25 = {inputSelect1H_9[25], inputSelect1H_8[25]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_25 = {inputSelect1H_11[25], inputSelect1H_10[25]};
  wire [3:0]  tryToRead_lo_hi_lo_25 = {tryToRead_lo_hi_lo_hi_25, tryToRead_lo_hi_lo_lo_25};
  wire [1:0]  tryToRead_lo_hi_hi_lo_25 = {inputSelect1H_13[25], inputSelect1H_12[25]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_25 = {inputSelect1H_15[25], inputSelect1H_14[25]};
  wire [3:0]  tryToRead_lo_hi_hi_25 = {tryToRead_lo_hi_hi_hi_25, tryToRead_lo_hi_hi_lo_25};
  wire [7:0]  tryToRead_lo_hi_25 = {tryToRead_lo_hi_hi_25, tryToRead_lo_hi_lo_25};
  wire [15:0] tryToRead_lo_25 = {tryToRead_lo_hi_25, tryToRead_lo_lo_25};
  wire [1:0]  tryToRead_hi_lo_lo_lo_25 = {inputSelect1H_17[25], inputSelect1H_16[25]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_25 = {inputSelect1H_19[25], inputSelect1H_18[25]};
  wire [3:0]  tryToRead_hi_lo_lo_25 = {tryToRead_hi_lo_lo_hi_25, tryToRead_hi_lo_lo_lo_25};
  wire [1:0]  tryToRead_hi_lo_hi_lo_25 = {inputSelect1H_21[25], inputSelect1H_20[25]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_25 = {inputSelect1H_23[25], inputSelect1H_22[25]};
  wire [3:0]  tryToRead_hi_lo_hi_25 = {tryToRead_hi_lo_hi_hi_25, tryToRead_hi_lo_hi_lo_25};
  wire [7:0]  tryToRead_hi_lo_25 = {tryToRead_hi_lo_hi_25, tryToRead_hi_lo_lo_25};
  wire [1:0]  tryToRead_hi_hi_lo_lo_25 = {inputSelect1H_25[25], inputSelect1H_24[25]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_25 = {inputSelect1H_27[25], inputSelect1H_26[25]};
  wire [3:0]  tryToRead_hi_hi_lo_25 = {tryToRead_hi_hi_lo_hi_25, tryToRead_hi_hi_lo_lo_25};
  wire [1:0]  tryToRead_hi_hi_hi_lo_25 = {inputSelect1H_29[25], inputSelect1H_28[25]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_25 = {inputSelect1H_31[25], inputSelect1H_30[25]};
  wire [3:0]  tryToRead_hi_hi_hi_25 = {tryToRead_hi_hi_hi_hi_25, tryToRead_hi_hi_hi_lo_25};
  wire [7:0]  tryToRead_hi_hi_25 = {tryToRead_hi_hi_hi_25, tryToRead_hi_hi_lo_25};
  wire [15:0] tryToRead_hi_25 = {tryToRead_hi_hi_25, tryToRead_hi_lo_25};
  wire [31:0] tryToRead_25 = {tryToRead_hi_25, tryToRead_lo_25};
  wire        output_25_valid_0 = |tryToRead_25;
  wire [4:0]  output_25_bits_vs_0 = selectReq_25_bits_vs;
  wire        output_25_bits_offset_0 = selectReq_25_bits_offset;
  wire [4:0]  output_25_bits_writeIndex_0 = selectReq_25_bits_requestIndex;
  wire [1:0]  output_25_bits_dataOffset_0 = selectReq_25_bits_dataOffset;
  assign selectReq_25_bits_dataOffset =
    (tryToRead_25[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_25[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_25[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_25[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_25[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_25[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_25[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_25[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_25[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_25[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_25[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_25[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_25[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_25[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_25[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_25[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_25[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_25[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_25[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_25[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_25[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_25[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_25[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_25[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_25[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_25[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_25_bits_requestIndex =
    {4'h0, tryToRead_25[1]} | {3'h0, tryToRead_25[2], 1'h0} | (tryToRead_25[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_25[4], 2'h0} | (tryToRead_25[5] ? 5'h5 : 5'h0) | (tryToRead_25[6] ? 5'h6 : 5'h0) | (tryToRead_25[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_25[8], 3'h0} | (tryToRead_25[9] ? 5'h9 : 5'h0) | (tryToRead_25[10] ? 5'hA : 5'h0) | (tryToRead_25[11] ? 5'hB : 5'h0) | (tryToRead_25[12] ? 5'hC : 5'h0) | (tryToRead_25[13] ? 5'hD : 5'h0)
    | (tryToRead_25[14] ? 5'hE : 5'h0) | (tryToRead_25[15] ? 5'hF : 5'h0) | {tryToRead_25[16], 4'h0} | (tryToRead_25[17] ? 5'h11 : 5'h0) | (tryToRead_25[18] ? 5'h12 : 5'h0) | (tryToRead_25[19] ? 5'h13 : 5'h0)
    | (tryToRead_25[20] ? 5'h14 : 5'h0) | (tryToRead_25[21] ? 5'h15 : 5'h0) | (tryToRead_25[22] ? 5'h16 : 5'h0) | (tryToRead_25[23] ? 5'h17 : 5'h0) | (tryToRead_25[24] ? 5'h18 : 5'h0) | (tryToRead_25[25] ? 5'h19 : 5'h0)
    | (tryToRead_25[26] ? 5'h1A : 5'h0) | (tryToRead_25[27] ? 5'h1B : 5'h0) | (tryToRead_25[28] ? 5'h1C : 5'h0) | (tryToRead_25[29] ? 5'h1D : 5'h0) | (tryToRead_25[30] ? 5'h1E : 5'h0) | {5{tryToRead_25[31]}};
  wire [4:0]  selectReq_25_bits_readLane =
    (tryToRead_25[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_25[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_25[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_25[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_25[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_25[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_25[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_25[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_25[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_25[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_25[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_25[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_25[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_25[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_25[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_25[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_25[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_25[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_25[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_25[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_25[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_25[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_25[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_25[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_25[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_25[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_25[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_25[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_25[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_25[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_25[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_25[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_25_bits_offset =
    tryToRead_25[0] & input_0_bits_offset_0 | tryToRead_25[1] & input_1_bits_offset_0 | tryToRead_25[2] & input_2_bits_offset_0 | tryToRead_25[3] & input_3_bits_offset_0 | tryToRead_25[4] & input_4_bits_offset_0 | tryToRead_25[5]
    & input_5_bits_offset_0 | tryToRead_25[6] & input_6_bits_offset_0 | tryToRead_25[7] & input_7_bits_offset_0 | tryToRead_25[8] & input_8_bits_offset_0 | tryToRead_25[9] & input_9_bits_offset_0 | tryToRead_25[10] & input_10_bits_offset_0
    | tryToRead_25[11] & input_11_bits_offset_0 | tryToRead_25[12] & input_12_bits_offset_0 | tryToRead_25[13] & input_13_bits_offset_0 | tryToRead_25[14] & input_14_bits_offset_0 | tryToRead_25[15] & input_15_bits_offset_0
    | tryToRead_25[16] & input_16_bits_offset_0 | tryToRead_25[17] & input_17_bits_offset_0 | tryToRead_25[18] & input_18_bits_offset_0 | tryToRead_25[19] & input_19_bits_offset_0 | tryToRead_25[20] & input_20_bits_offset_0
    | tryToRead_25[21] & input_21_bits_offset_0 | tryToRead_25[22] & input_22_bits_offset_0 | tryToRead_25[23] & input_23_bits_offset_0 | tryToRead_25[24] & input_24_bits_offset_0 | tryToRead_25[25] & input_25_bits_offset_0
    | tryToRead_25[26] & input_26_bits_offset_0 | tryToRead_25[27] & input_27_bits_offset_0 | tryToRead_25[28] & input_28_bits_offset_0 | tryToRead_25[29] & input_29_bits_offset_0 | tryToRead_25[30] & input_30_bits_offset_0
    | tryToRead_25[31] & input_31_bits_offset_0;
  assign selectReq_25_bits_vs =
    (tryToRead_25[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_25[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_25[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_25[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_25[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_25[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_25[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_25[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_25[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_25[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_25[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_25[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_25[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_25[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_25[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_25[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_25[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_25[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_25[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_25[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_25[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_25[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_25[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_25[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_25[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_25[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_25[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_25[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_25[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_25[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_25[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_25[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_25_valid =
    tryToRead_25[0] & input_0_valid_0 | tryToRead_25[1] & input_1_valid_0 | tryToRead_25[2] & input_2_valid_0 | tryToRead_25[3] & input_3_valid_0 | tryToRead_25[4] & input_4_valid_0 | tryToRead_25[5] & input_5_valid_0 | tryToRead_25[6]
    & input_6_valid_0 | tryToRead_25[7] & input_7_valid_0 | tryToRead_25[8] & input_8_valid_0 | tryToRead_25[9] & input_9_valid_0 | tryToRead_25[10] & input_10_valid_0 | tryToRead_25[11] & input_11_valid_0 | tryToRead_25[12]
    & input_12_valid_0 | tryToRead_25[13] & input_13_valid_0 | tryToRead_25[14] & input_14_valid_0 | tryToRead_25[15] & input_15_valid_0 | tryToRead_25[16] & input_16_valid_0 | tryToRead_25[17] & input_17_valid_0 | tryToRead_25[18]
    & input_18_valid_0 | tryToRead_25[19] & input_19_valid_0 | tryToRead_25[20] & input_20_valid_0 | tryToRead_25[21] & input_21_valid_0 | tryToRead_25[22] & input_22_valid_0 | tryToRead_25[23] & input_23_valid_0 | tryToRead_25[24]
    & input_24_valid_0 | tryToRead_25[25] & input_25_valid_0 | tryToRead_25[26] & input_26_valid_0 | tryToRead_25[27] & input_27_valid_0 | tryToRead_25[28] & input_28_valid_0 | tryToRead_25[29] & input_29_valid_0 | tryToRead_25[30]
    & input_30_valid_0 | tryToRead_25[31] & input_31_valid_0;
  wire        selectReq_25_ready =
    tryToRead_25[0] & input_0_ready_0 | tryToRead_25[1] & input_1_ready_0 | tryToRead_25[2] & input_2_ready_0 | tryToRead_25[3] & input_3_ready_0 | tryToRead_25[4] & input_4_ready_0 | tryToRead_25[5] & input_5_ready_0 | tryToRead_25[6]
    & input_6_ready_0 | tryToRead_25[7] & input_7_ready_0 | tryToRead_25[8] & input_8_ready_0 | tryToRead_25[9] & input_9_ready_0 | tryToRead_25[10] & input_10_ready_0 | tryToRead_25[11] & input_11_ready_0 | tryToRead_25[12]
    & input_12_ready_0 | tryToRead_25[13] & input_13_ready_0 | tryToRead_25[14] & input_14_ready_0 | tryToRead_25[15] & input_15_ready_0 | tryToRead_25[16] & input_16_ready_0 | tryToRead_25[17] & input_17_ready_0 | tryToRead_25[18]
    & input_18_ready_0 | tryToRead_25[19] & input_19_ready_0 | tryToRead_25[20] & input_20_ready_0 | tryToRead_25[21] & input_21_ready_0 | tryToRead_25[22] & input_22_ready_0 | tryToRead_25[23] & input_23_ready_0 | tryToRead_25[24]
    & input_24_ready_0 | tryToRead_25[25] & input_25_ready_0 | tryToRead_25[26] & input_26_ready_0 | tryToRead_25[27] & input_27_ready_0 | tryToRead_25[28] & input_28_ready_0 | tryToRead_25[29] & input_29_ready_0 | tryToRead_25[30]
    & input_30_ready_0 | tryToRead_25[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_26 = {inputSelect1H_1[26], inputSelect1H_0[26]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_26 = {inputSelect1H_3[26], inputSelect1H_2[26]};
  wire [3:0]  tryToRead_lo_lo_lo_26 = {tryToRead_lo_lo_lo_hi_26, tryToRead_lo_lo_lo_lo_26};
  wire [1:0]  tryToRead_lo_lo_hi_lo_26 = {inputSelect1H_5[26], inputSelect1H_4[26]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_26 = {inputSelect1H_7[26], inputSelect1H_6[26]};
  wire [3:0]  tryToRead_lo_lo_hi_26 = {tryToRead_lo_lo_hi_hi_26, tryToRead_lo_lo_hi_lo_26};
  wire [7:0]  tryToRead_lo_lo_26 = {tryToRead_lo_lo_hi_26, tryToRead_lo_lo_lo_26};
  wire [1:0]  tryToRead_lo_hi_lo_lo_26 = {inputSelect1H_9[26], inputSelect1H_8[26]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_26 = {inputSelect1H_11[26], inputSelect1H_10[26]};
  wire [3:0]  tryToRead_lo_hi_lo_26 = {tryToRead_lo_hi_lo_hi_26, tryToRead_lo_hi_lo_lo_26};
  wire [1:0]  tryToRead_lo_hi_hi_lo_26 = {inputSelect1H_13[26], inputSelect1H_12[26]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_26 = {inputSelect1H_15[26], inputSelect1H_14[26]};
  wire [3:0]  tryToRead_lo_hi_hi_26 = {tryToRead_lo_hi_hi_hi_26, tryToRead_lo_hi_hi_lo_26};
  wire [7:0]  tryToRead_lo_hi_26 = {tryToRead_lo_hi_hi_26, tryToRead_lo_hi_lo_26};
  wire [15:0] tryToRead_lo_26 = {tryToRead_lo_hi_26, tryToRead_lo_lo_26};
  wire [1:0]  tryToRead_hi_lo_lo_lo_26 = {inputSelect1H_17[26], inputSelect1H_16[26]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_26 = {inputSelect1H_19[26], inputSelect1H_18[26]};
  wire [3:0]  tryToRead_hi_lo_lo_26 = {tryToRead_hi_lo_lo_hi_26, tryToRead_hi_lo_lo_lo_26};
  wire [1:0]  tryToRead_hi_lo_hi_lo_26 = {inputSelect1H_21[26], inputSelect1H_20[26]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_26 = {inputSelect1H_23[26], inputSelect1H_22[26]};
  wire [3:0]  tryToRead_hi_lo_hi_26 = {tryToRead_hi_lo_hi_hi_26, tryToRead_hi_lo_hi_lo_26};
  wire [7:0]  tryToRead_hi_lo_26 = {tryToRead_hi_lo_hi_26, tryToRead_hi_lo_lo_26};
  wire [1:0]  tryToRead_hi_hi_lo_lo_26 = {inputSelect1H_25[26], inputSelect1H_24[26]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_26 = {inputSelect1H_27[26], inputSelect1H_26[26]};
  wire [3:0]  tryToRead_hi_hi_lo_26 = {tryToRead_hi_hi_lo_hi_26, tryToRead_hi_hi_lo_lo_26};
  wire [1:0]  tryToRead_hi_hi_hi_lo_26 = {inputSelect1H_29[26], inputSelect1H_28[26]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_26 = {inputSelect1H_31[26], inputSelect1H_30[26]};
  wire [3:0]  tryToRead_hi_hi_hi_26 = {tryToRead_hi_hi_hi_hi_26, tryToRead_hi_hi_hi_lo_26};
  wire [7:0]  tryToRead_hi_hi_26 = {tryToRead_hi_hi_hi_26, tryToRead_hi_hi_lo_26};
  wire [15:0] tryToRead_hi_26 = {tryToRead_hi_hi_26, tryToRead_hi_lo_26};
  wire [31:0] tryToRead_26 = {tryToRead_hi_26, tryToRead_lo_26};
  wire        output_26_valid_0 = |tryToRead_26;
  wire [4:0]  output_26_bits_vs_0 = selectReq_26_bits_vs;
  wire        output_26_bits_offset_0 = selectReq_26_bits_offset;
  wire [4:0]  output_26_bits_writeIndex_0 = selectReq_26_bits_requestIndex;
  wire [1:0]  output_26_bits_dataOffset_0 = selectReq_26_bits_dataOffset;
  assign selectReq_26_bits_dataOffset =
    (tryToRead_26[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_26[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_26[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_26[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_26[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_26[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_26[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_26[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_26[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_26[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_26[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_26[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_26[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_26[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_26[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_26[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_26[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_26[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_26[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_26[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_26[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_26[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_26[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_26[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_26[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_26[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_26_bits_requestIndex =
    {4'h0, tryToRead_26[1]} | {3'h0, tryToRead_26[2], 1'h0} | (tryToRead_26[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_26[4], 2'h0} | (tryToRead_26[5] ? 5'h5 : 5'h0) | (tryToRead_26[6] ? 5'h6 : 5'h0) | (tryToRead_26[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_26[8], 3'h0} | (tryToRead_26[9] ? 5'h9 : 5'h0) | (tryToRead_26[10] ? 5'hA : 5'h0) | (tryToRead_26[11] ? 5'hB : 5'h0) | (tryToRead_26[12] ? 5'hC : 5'h0) | (tryToRead_26[13] ? 5'hD : 5'h0)
    | (tryToRead_26[14] ? 5'hE : 5'h0) | (tryToRead_26[15] ? 5'hF : 5'h0) | {tryToRead_26[16], 4'h0} | (tryToRead_26[17] ? 5'h11 : 5'h0) | (tryToRead_26[18] ? 5'h12 : 5'h0) | (tryToRead_26[19] ? 5'h13 : 5'h0)
    | (tryToRead_26[20] ? 5'h14 : 5'h0) | (tryToRead_26[21] ? 5'h15 : 5'h0) | (tryToRead_26[22] ? 5'h16 : 5'h0) | (tryToRead_26[23] ? 5'h17 : 5'h0) | (tryToRead_26[24] ? 5'h18 : 5'h0) | (tryToRead_26[25] ? 5'h19 : 5'h0)
    | (tryToRead_26[26] ? 5'h1A : 5'h0) | (tryToRead_26[27] ? 5'h1B : 5'h0) | (tryToRead_26[28] ? 5'h1C : 5'h0) | (tryToRead_26[29] ? 5'h1D : 5'h0) | (tryToRead_26[30] ? 5'h1E : 5'h0) | {5{tryToRead_26[31]}};
  wire [4:0]  selectReq_26_bits_readLane =
    (tryToRead_26[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_26[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_26[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_26[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_26[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_26[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_26[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_26[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_26[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_26[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_26[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_26[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_26[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_26[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_26[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_26[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_26[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_26[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_26[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_26[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_26[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_26[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_26[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_26[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_26[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_26[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_26[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_26[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_26[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_26[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_26[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_26[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_26_bits_offset =
    tryToRead_26[0] & input_0_bits_offset_0 | tryToRead_26[1] & input_1_bits_offset_0 | tryToRead_26[2] & input_2_bits_offset_0 | tryToRead_26[3] & input_3_bits_offset_0 | tryToRead_26[4] & input_4_bits_offset_0 | tryToRead_26[5]
    & input_5_bits_offset_0 | tryToRead_26[6] & input_6_bits_offset_0 | tryToRead_26[7] & input_7_bits_offset_0 | tryToRead_26[8] & input_8_bits_offset_0 | tryToRead_26[9] & input_9_bits_offset_0 | tryToRead_26[10] & input_10_bits_offset_0
    | tryToRead_26[11] & input_11_bits_offset_0 | tryToRead_26[12] & input_12_bits_offset_0 | tryToRead_26[13] & input_13_bits_offset_0 | tryToRead_26[14] & input_14_bits_offset_0 | tryToRead_26[15] & input_15_bits_offset_0
    | tryToRead_26[16] & input_16_bits_offset_0 | tryToRead_26[17] & input_17_bits_offset_0 | tryToRead_26[18] & input_18_bits_offset_0 | tryToRead_26[19] & input_19_bits_offset_0 | tryToRead_26[20] & input_20_bits_offset_0
    | tryToRead_26[21] & input_21_bits_offset_0 | tryToRead_26[22] & input_22_bits_offset_0 | tryToRead_26[23] & input_23_bits_offset_0 | tryToRead_26[24] & input_24_bits_offset_0 | tryToRead_26[25] & input_25_bits_offset_0
    | tryToRead_26[26] & input_26_bits_offset_0 | tryToRead_26[27] & input_27_bits_offset_0 | tryToRead_26[28] & input_28_bits_offset_0 | tryToRead_26[29] & input_29_bits_offset_0 | tryToRead_26[30] & input_30_bits_offset_0
    | tryToRead_26[31] & input_31_bits_offset_0;
  assign selectReq_26_bits_vs =
    (tryToRead_26[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_26[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_26[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_26[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_26[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_26[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_26[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_26[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_26[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_26[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_26[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_26[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_26[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_26[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_26[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_26[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_26[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_26[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_26[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_26[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_26[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_26[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_26[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_26[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_26[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_26[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_26[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_26[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_26[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_26[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_26[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_26[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_26_valid =
    tryToRead_26[0] & input_0_valid_0 | tryToRead_26[1] & input_1_valid_0 | tryToRead_26[2] & input_2_valid_0 | tryToRead_26[3] & input_3_valid_0 | tryToRead_26[4] & input_4_valid_0 | tryToRead_26[5] & input_5_valid_0 | tryToRead_26[6]
    & input_6_valid_0 | tryToRead_26[7] & input_7_valid_0 | tryToRead_26[8] & input_8_valid_0 | tryToRead_26[9] & input_9_valid_0 | tryToRead_26[10] & input_10_valid_0 | tryToRead_26[11] & input_11_valid_0 | tryToRead_26[12]
    & input_12_valid_0 | tryToRead_26[13] & input_13_valid_0 | tryToRead_26[14] & input_14_valid_0 | tryToRead_26[15] & input_15_valid_0 | tryToRead_26[16] & input_16_valid_0 | tryToRead_26[17] & input_17_valid_0 | tryToRead_26[18]
    & input_18_valid_0 | tryToRead_26[19] & input_19_valid_0 | tryToRead_26[20] & input_20_valid_0 | tryToRead_26[21] & input_21_valid_0 | tryToRead_26[22] & input_22_valid_0 | tryToRead_26[23] & input_23_valid_0 | tryToRead_26[24]
    & input_24_valid_0 | tryToRead_26[25] & input_25_valid_0 | tryToRead_26[26] & input_26_valid_0 | tryToRead_26[27] & input_27_valid_0 | tryToRead_26[28] & input_28_valid_0 | tryToRead_26[29] & input_29_valid_0 | tryToRead_26[30]
    & input_30_valid_0 | tryToRead_26[31] & input_31_valid_0;
  wire        selectReq_26_ready =
    tryToRead_26[0] & input_0_ready_0 | tryToRead_26[1] & input_1_ready_0 | tryToRead_26[2] & input_2_ready_0 | tryToRead_26[3] & input_3_ready_0 | tryToRead_26[4] & input_4_ready_0 | tryToRead_26[5] & input_5_ready_0 | tryToRead_26[6]
    & input_6_ready_0 | tryToRead_26[7] & input_7_ready_0 | tryToRead_26[8] & input_8_ready_0 | tryToRead_26[9] & input_9_ready_0 | tryToRead_26[10] & input_10_ready_0 | tryToRead_26[11] & input_11_ready_0 | tryToRead_26[12]
    & input_12_ready_0 | tryToRead_26[13] & input_13_ready_0 | tryToRead_26[14] & input_14_ready_0 | tryToRead_26[15] & input_15_ready_0 | tryToRead_26[16] & input_16_ready_0 | tryToRead_26[17] & input_17_ready_0 | tryToRead_26[18]
    & input_18_ready_0 | tryToRead_26[19] & input_19_ready_0 | tryToRead_26[20] & input_20_ready_0 | tryToRead_26[21] & input_21_ready_0 | tryToRead_26[22] & input_22_ready_0 | tryToRead_26[23] & input_23_ready_0 | tryToRead_26[24]
    & input_24_ready_0 | tryToRead_26[25] & input_25_ready_0 | tryToRead_26[26] & input_26_ready_0 | tryToRead_26[27] & input_27_ready_0 | tryToRead_26[28] & input_28_ready_0 | tryToRead_26[29] & input_29_ready_0 | tryToRead_26[30]
    & input_30_ready_0 | tryToRead_26[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_27 = {inputSelect1H_1[27], inputSelect1H_0[27]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_27 = {inputSelect1H_3[27], inputSelect1H_2[27]};
  wire [3:0]  tryToRead_lo_lo_lo_27 = {tryToRead_lo_lo_lo_hi_27, tryToRead_lo_lo_lo_lo_27};
  wire [1:0]  tryToRead_lo_lo_hi_lo_27 = {inputSelect1H_5[27], inputSelect1H_4[27]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_27 = {inputSelect1H_7[27], inputSelect1H_6[27]};
  wire [3:0]  tryToRead_lo_lo_hi_27 = {tryToRead_lo_lo_hi_hi_27, tryToRead_lo_lo_hi_lo_27};
  wire [7:0]  tryToRead_lo_lo_27 = {tryToRead_lo_lo_hi_27, tryToRead_lo_lo_lo_27};
  wire [1:0]  tryToRead_lo_hi_lo_lo_27 = {inputSelect1H_9[27], inputSelect1H_8[27]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_27 = {inputSelect1H_11[27], inputSelect1H_10[27]};
  wire [3:0]  tryToRead_lo_hi_lo_27 = {tryToRead_lo_hi_lo_hi_27, tryToRead_lo_hi_lo_lo_27};
  wire [1:0]  tryToRead_lo_hi_hi_lo_27 = {inputSelect1H_13[27], inputSelect1H_12[27]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_27 = {inputSelect1H_15[27], inputSelect1H_14[27]};
  wire [3:0]  tryToRead_lo_hi_hi_27 = {tryToRead_lo_hi_hi_hi_27, tryToRead_lo_hi_hi_lo_27};
  wire [7:0]  tryToRead_lo_hi_27 = {tryToRead_lo_hi_hi_27, tryToRead_lo_hi_lo_27};
  wire [15:0] tryToRead_lo_27 = {tryToRead_lo_hi_27, tryToRead_lo_lo_27};
  wire [1:0]  tryToRead_hi_lo_lo_lo_27 = {inputSelect1H_17[27], inputSelect1H_16[27]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_27 = {inputSelect1H_19[27], inputSelect1H_18[27]};
  wire [3:0]  tryToRead_hi_lo_lo_27 = {tryToRead_hi_lo_lo_hi_27, tryToRead_hi_lo_lo_lo_27};
  wire [1:0]  tryToRead_hi_lo_hi_lo_27 = {inputSelect1H_21[27], inputSelect1H_20[27]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_27 = {inputSelect1H_23[27], inputSelect1H_22[27]};
  wire [3:0]  tryToRead_hi_lo_hi_27 = {tryToRead_hi_lo_hi_hi_27, tryToRead_hi_lo_hi_lo_27};
  wire [7:0]  tryToRead_hi_lo_27 = {tryToRead_hi_lo_hi_27, tryToRead_hi_lo_lo_27};
  wire [1:0]  tryToRead_hi_hi_lo_lo_27 = {inputSelect1H_25[27], inputSelect1H_24[27]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_27 = {inputSelect1H_27[27], inputSelect1H_26[27]};
  wire [3:0]  tryToRead_hi_hi_lo_27 = {tryToRead_hi_hi_lo_hi_27, tryToRead_hi_hi_lo_lo_27};
  wire [1:0]  tryToRead_hi_hi_hi_lo_27 = {inputSelect1H_29[27], inputSelect1H_28[27]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_27 = {inputSelect1H_31[27], inputSelect1H_30[27]};
  wire [3:0]  tryToRead_hi_hi_hi_27 = {tryToRead_hi_hi_hi_hi_27, tryToRead_hi_hi_hi_lo_27};
  wire [7:0]  tryToRead_hi_hi_27 = {tryToRead_hi_hi_hi_27, tryToRead_hi_hi_lo_27};
  wire [15:0] tryToRead_hi_27 = {tryToRead_hi_hi_27, tryToRead_hi_lo_27};
  wire [31:0] tryToRead_27 = {tryToRead_hi_27, tryToRead_lo_27};
  wire        output_27_valid_0 = |tryToRead_27;
  wire [4:0]  output_27_bits_vs_0 = selectReq_27_bits_vs;
  wire        output_27_bits_offset_0 = selectReq_27_bits_offset;
  wire [4:0]  output_27_bits_writeIndex_0 = selectReq_27_bits_requestIndex;
  wire [1:0]  output_27_bits_dataOffset_0 = selectReq_27_bits_dataOffset;
  assign selectReq_27_bits_dataOffset =
    (tryToRead_27[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_27[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_27[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_27[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_27[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_27[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_27[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_27[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_27[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_27[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_27[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_27[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_27[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_27[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_27[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_27[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_27[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_27[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_27[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_27[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_27[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_27[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_27[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_27[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_27[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_27[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_27_bits_requestIndex =
    {4'h0, tryToRead_27[1]} | {3'h0, tryToRead_27[2], 1'h0} | (tryToRead_27[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_27[4], 2'h0} | (tryToRead_27[5] ? 5'h5 : 5'h0) | (tryToRead_27[6] ? 5'h6 : 5'h0) | (tryToRead_27[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_27[8], 3'h0} | (tryToRead_27[9] ? 5'h9 : 5'h0) | (tryToRead_27[10] ? 5'hA : 5'h0) | (tryToRead_27[11] ? 5'hB : 5'h0) | (tryToRead_27[12] ? 5'hC : 5'h0) | (tryToRead_27[13] ? 5'hD : 5'h0)
    | (tryToRead_27[14] ? 5'hE : 5'h0) | (tryToRead_27[15] ? 5'hF : 5'h0) | {tryToRead_27[16], 4'h0} | (tryToRead_27[17] ? 5'h11 : 5'h0) | (tryToRead_27[18] ? 5'h12 : 5'h0) | (tryToRead_27[19] ? 5'h13 : 5'h0)
    | (tryToRead_27[20] ? 5'h14 : 5'h0) | (tryToRead_27[21] ? 5'h15 : 5'h0) | (tryToRead_27[22] ? 5'h16 : 5'h0) | (tryToRead_27[23] ? 5'h17 : 5'h0) | (tryToRead_27[24] ? 5'h18 : 5'h0) | (tryToRead_27[25] ? 5'h19 : 5'h0)
    | (tryToRead_27[26] ? 5'h1A : 5'h0) | (tryToRead_27[27] ? 5'h1B : 5'h0) | (tryToRead_27[28] ? 5'h1C : 5'h0) | (tryToRead_27[29] ? 5'h1D : 5'h0) | (tryToRead_27[30] ? 5'h1E : 5'h0) | {5{tryToRead_27[31]}};
  wire [4:0]  selectReq_27_bits_readLane =
    (tryToRead_27[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_27[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_27[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_27[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_27[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_27[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_27[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_27[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_27[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_27[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_27[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_27[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_27[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_27[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_27[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_27[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_27[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_27[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_27[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_27[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_27[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_27[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_27[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_27[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_27[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_27[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_27[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_27[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_27[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_27[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_27[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_27[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_27_bits_offset =
    tryToRead_27[0] & input_0_bits_offset_0 | tryToRead_27[1] & input_1_bits_offset_0 | tryToRead_27[2] & input_2_bits_offset_0 | tryToRead_27[3] & input_3_bits_offset_0 | tryToRead_27[4] & input_4_bits_offset_0 | tryToRead_27[5]
    & input_5_bits_offset_0 | tryToRead_27[6] & input_6_bits_offset_0 | tryToRead_27[7] & input_7_bits_offset_0 | tryToRead_27[8] & input_8_bits_offset_0 | tryToRead_27[9] & input_9_bits_offset_0 | tryToRead_27[10] & input_10_bits_offset_0
    | tryToRead_27[11] & input_11_bits_offset_0 | tryToRead_27[12] & input_12_bits_offset_0 | tryToRead_27[13] & input_13_bits_offset_0 | tryToRead_27[14] & input_14_bits_offset_0 | tryToRead_27[15] & input_15_bits_offset_0
    | tryToRead_27[16] & input_16_bits_offset_0 | tryToRead_27[17] & input_17_bits_offset_0 | tryToRead_27[18] & input_18_bits_offset_0 | tryToRead_27[19] & input_19_bits_offset_0 | tryToRead_27[20] & input_20_bits_offset_0
    | tryToRead_27[21] & input_21_bits_offset_0 | tryToRead_27[22] & input_22_bits_offset_0 | tryToRead_27[23] & input_23_bits_offset_0 | tryToRead_27[24] & input_24_bits_offset_0 | tryToRead_27[25] & input_25_bits_offset_0
    | tryToRead_27[26] & input_26_bits_offset_0 | tryToRead_27[27] & input_27_bits_offset_0 | tryToRead_27[28] & input_28_bits_offset_0 | tryToRead_27[29] & input_29_bits_offset_0 | tryToRead_27[30] & input_30_bits_offset_0
    | tryToRead_27[31] & input_31_bits_offset_0;
  assign selectReq_27_bits_vs =
    (tryToRead_27[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_27[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_27[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_27[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_27[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_27[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_27[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_27[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_27[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_27[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_27[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_27[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_27[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_27[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_27[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_27[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_27[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_27[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_27[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_27[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_27[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_27[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_27[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_27[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_27[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_27[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_27[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_27[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_27[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_27[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_27[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_27[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_27_valid =
    tryToRead_27[0] & input_0_valid_0 | tryToRead_27[1] & input_1_valid_0 | tryToRead_27[2] & input_2_valid_0 | tryToRead_27[3] & input_3_valid_0 | tryToRead_27[4] & input_4_valid_0 | tryToRead_27[5] & input_5_valid_0 | tryToRead_27[6]
    & input_6_valid_0 | tryToRead_27[7] & input_7_valid_0 | tryToRead_27[8] & input_8_valid_0 | tryToRead_27[9] & input_9_valid_0 | tryToRead_27[10] & input_10_valid_0 | tryToRead_27[11] & input_11_valid_0 | tryToRead_27[12]
    & input_12_valid_0 | tryToRead_27[13] & input_13_valid_0 | tryToRead_27[14] & input_14_valid_0 | tryToRead_27[15] & input_15_valid_0 | tryToRead_27[16] & input_16_valid_0 | tryToRead_27[17] & input_17_valid_0 | tryToRead_27[18]
    & input_18_valid_0 | tryToRead_27[19] & input_19_valid_0 | tryToRead_27[20] & input_20_valid_0 | tryToRead_27[21] & input_21_valid_0 | tryToRead_27[22] & input_22_valid_0 | tryToRead_27[23] & input_23_valid_0 | tryToRead_27[24]
    & input_24_valid_0 | tryToRead_27[25] & input_25_valid_0 | tryToRead_27[26] & input_26_valid_0 | tryToRead_27[27] & input_27_valid_0 | tryToRead_27[28] & input_28_valid_0 | tryToRead_27[29] & input_29_valid_0 | tryToRead_27[30]
    & input_30_valid_0 | tryToRead_27[31] & input_31_valid_0;
  wire        selectReq_27_ready =
    tryToRead_27[0] & input_0_ready_0 | tryToRead_27[1] & input_1_ready_0 | tryToRead_27[2] & input_2_ready_0 | tryToRead_27[3] & input_3_ready_0 | tryToRead_27[4] & input_4_ready_0 | tryToRead_27[5] & input_5_ready_0 | tryToRead_27[6]
    & input_6_ready_0 | tryToRead_27[7] & input_7_ready_0 | tryToRead_27[8] & input_8_ready_0 | tryToRead_27[9] & input_9_ready_0 | tryToRead_27[10] & input_10_ready_0 | tryToRead_27[11] & input_11_ready_0 | tryToRead_27[12]
    & input_12_ready_0 | tryToRead_27[13] & input_13_ready_0 | tryToRead_27[14] & input_14_ready_0 | tryToRead_27[15] & input_15_ready_0 | tryToRead_27[16] & input_16_ready_0 | tryToRead_27[17] & input_17_ready_0 | tryToRead_27[18]
    & input_18_ready_0 | tryToRead_27[19] & input_19_ready_0 | tryToRead_27[20] & input_20_ready_0 | tryToRead_27[21] & input_21_ready_0 | tryToRead_27[22] & input_22_ready_0 | tryToRead_27[23] & input_23_ready_0 | tryToRead_27[24]
    & input_24_ready_0 | tryToRead_27[25] & input_25_ready_0 | tryToRead_27[26] & input_26_ready_0 | tryToRead_27[27] & input_27_ready_0 | tryToRead_27[28] & input_28_ready_0 | tryToRead_27[29] & input_29_ready_0 | tryToRead_27[30]
    & input_30_ready_0 | tryToRead_27[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_28 = {inputSelect1H_1[28], inputSelect1H_0[28]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_28 = {inputSelect1H_3[28], inputSelect1H_2[28]};
  wire [3:0]  tryToRead_lo_lo_lo_28 = {tryToRead_lo_lo_lo_hi_28, tryToRead_lo_lo_lo_lo_28};
  wire [1:0]  tryToRead_lo_lo_hi_lo_28 = {inputSelect1H_5[28], inputSelect1H_4[28]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_28 = {inputSelect1H_7[28], inputSelect1H_6[28]};
  wire [3:0]  tryToRead_lo_lo_hi_28 = {tryToRead_lo_lo_hi_hi_28, tryToRead_lo_lo_hi_lo_28};
  wire [7:0]  tryToRead_lo_lo_28 = {tryToRead_lo_lo_hi_28, tryToRead_lo_lo_lo_28};
  wire [1:0]  tryToRead_lo_hi_lo_lo_28 = {inputSelect1H_9[28], inputSelect1H_8[28]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_28 = {inputSelect1H_11[28], inputSelect1H_10[28]};
  wire [3:0]  tryToRead_lo_hi_lo_28 = {tryToRead_lo_hi_lo_hi_28, tryToRead_lo_hi_lo_lo_28};
  wire [1:0]  tryToRead_lo_hi_hi_lo_28 = {inputSelect1H_13[28], inputSelect1H_12[28]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_28 = {inputSelect1H_15[28], inputSelect1H_14[28]};
  wire [3:0]  tryToRead_lo_hi_hi_28 = {tryToRead_lo_hi_hi_hi_28, tryToRead_lo_hi_hi_lo_28};
  wire [7:0]  tryToRead_lo_hi_28 = {tryToRead_lo_hi_hi_28, tryToRead_lo_hi_lo_28};
  wire [15:0] tryToRead_lo_28 = {tryToRead_lo_hi_28, tryToRead_lo_lo_28};
  wire [1:0]  tryToRead_hi_lo_lo_lo_28 = {inputSelect1H_17[28], inputSelect1H_16[28]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_28 = {inputSelect1H_19[28], inputSelect1H_18[28]};
  wire [3:0]  tryToRead_hi_lo_lo_28 = {tryToRead_hi_lo_lo_hi_28, tryToRead_hi_lo_lo_lo_28};
  wire [1:0]  tryToRead_hi_lo_hi_lo_28 = {inputSelect1H_21[28], inputSelect1H_20[28]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_28 = {inputSelect1H_23[28], inputSelect1H_22[28]};
  wire [3:0]  tryToRead_hi_lo_hi_28 = {tryToRead_hi_lo_hi_hi_28, tryToRead_hi_lo_hi_lo_28};
  wire [7:0]  tryToRead_hi_lo_28 = {tryToRead_hi_lo_hi_28, tryToRead_hi_lo_lo_28};
  wire [1:0]  tryToRead_hi_hi_lo_lo_28 = {inputSelect1H_25[28], inputSelect1H_24[28]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_28 = {inputSelect1H_27[28], inputSelect1H_26[28]};
  wire [3:0]  tryToRead_hi_hi_lo_28 = {tryToRead_hi_hi_lo_hi_28, tryToRead_hi_hi_lo_lo_28};
  wire [1:0]  tryToRead_hi_hi_hi_lo_28 = {inputSelect1H_29[28], inputSelect1H_28[28]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_28 = {inputSelect1H_31[28], inputSelect1H_30[28]};
  wire [3:0]  tryToRead_hi_hi_hi_28 = {tryToRead_hi_hi_hi_hi_28, tryToRead_hi_hi_hi_lo_28};
  wire [7:0]  tryToRead_hi_hi_28 = {tryToRead_hi_hi_hi_28, tryToRead_hi_hi_lo_28};
  wire [15:0] tryToRead_hi_28 = {tryToRead_hi_hi_28, tryToRead_hi_lo_28};
  wire [31:0] tryToRead_28 = {tryToRead_hi_28, tryToRead_lo_28};
  wire        output_28_valid_0 = |tryToRead_28;
  wire [4:0]  output_28_bits_vs_0 = selectReq_28_bits_vs;
  wire        output_28_bits_offset_0 = selectReq_28_bits_offset;
  wire [4:0]  output_28_bits_writeIndex_0 = selectReq_28_bits_requestIndex;
  wire [1:0]  output_28_bits_dataOffset_0 = selectReq_28_bits_dataOffset;
  assign selectReq_28_bits_dataOffset =
    (tryToRead_28[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_28[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_28[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_28[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_28[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_28[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_28[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_28[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_28[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_28[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_28[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_28[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_28[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_28[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_28[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_28[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_28[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_28[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_28[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_28[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_28[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_28[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_28[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_28[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_28[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_28[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_28_bits_requestIndex =
    {4'h0, tryToRead_28[1]} | {3'h0, tryToRead_28[2], 1'h0} | (tryToRead_28[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_28[4], 2'h0} | (tryToRead_28[5] ? 5'h5 : 5'h0) | (tryToRead_28[6] ? 5'h6 : 5'h0) | (tryToRead_28[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_28[8], 3'h0} | (tryToRead_28[9] ? 5'h9 : 5'h0) | (tryToRead_28[10] ? 5'hA : 5'h0) | (tryToRead_28[11] ? 5'hB : 5'h0) | (tryToRead_28[12] ? 5'hC : 5'h0) | (tryToRead_28[13] ? 5'hD : 5'h0)
    | (tryToRead_28[14] ? 5'hE : 5'h0) | (tryToRead_28[15] ? 5'hF : 5'h0) | {tryToRead_28[16], 4'h0} | (tryToRead_28[17] ? 5'h11 : 5'h0) | (tryToRead_28[18] ? 5'h12 : 5'h0) | (tryToRead_28[19] ? 5'h13 : 5'h0)
    | (tryToRead_28[20] ? 5'h14 : 5'h0) | (tryToRead_28[21] ? 5'h15 : 5'h0) | (tryToRead_28[22] ? 5'h16 : 5'h0) | (tryToRead_28[23] ? 5'h17 : 5'h0) | (tryToRead_28[24] ? 5'h18 : 5'h0) | (tryToRead_28[25] ? 5'h19 : 5'h0)
    | (tryToRead_28[26] ? 5'h1A : 5'h0) | (tryToRead_28[27] ? 5'h1B : 5'h0) | (tryToRead_28[28] ? 5'h1C : 5'h0) | (tryToRead_28[29] ? 5'h1D : 5'h0) | (tryToRead_28[30] ? 5'h1E : 5'h0) | {5{tryToRead_28[31]}};
  wire [4:0]  selectReq_28_bits_readLane =
    (tryToRead_28[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_28[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_28[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_28[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_28[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_28[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_28[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_28[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_28[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_28[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_28[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_28[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_28[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_28[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_28[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_28[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_28[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_28[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_28[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_28[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_28[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_28[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_28[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_28[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_28[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_28[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_28[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_28[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_28[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_28[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_28[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_28[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_28_bits_offset =
    tryToRead_28[0] & input_0_bits_offset_0 | tryToRead_28[1] & input_1_bits_offset_0 | tryToRead_28[2] & input_2_bits_offset_0 | tryToRead_28[3] & input_3_bits_offset_0 | tryToRead_28[4] & input_4_bits_offset_0 | tryToRead_28[5]
    & input_5_bits_offset_0 | tryToRead_28[6] & input_6_bits_offset_0 | tryToRead_28[7] & input_7_bits_offset_0 | tryToRead_28[8] & input_8_bits_offset_0 | tryToRead_28[9] & input_9_bits_offset_0 | tryToRead_28[10] & input_10_bits_offset_0
    | tryToRead_28[11] & input_11_bits_offset_0 | tryToRead_28[12] & input_12_bits_offset_0 | tryToRead_28[13] & input_13_bits_offset_0 | tryToRead_28[14] & input_14_bits_offset_0 | tryToRead_28[15] & input_15_bits_offset_0
    | tryToRead_28[16] & input_16_bits_offset_0 | tryToRead_28[17] & input_17_bits_offset_0 | tryToRead_28[18] & input_18_bits_offset_0 | tryToRead_28[19] & input_19_bits_offset_0 | tryToRead_28[20] & input_20_bits_offset_0
    | tryToRead_28[21] & input_21_bits_offset_0 | tryToRead_28[22] & input_22_bits_offset_0 | tryToRead_28[23] & input_23_bits_offset_0 | tryToRead_28[24] & input_24_bits_offset_0 | tryToRead_28[25] & input_25_bits_offset_0
    | tryToRead_28[26] & input_26_bits_offset_0 | tryToRead_28[27] & input_27_bits_offset_0 | tryToRead_28[28] & input_28_bits_offset_0 | tryToRead_28[29] & input_29_bits_offset_0 | tryToRead_28[30] & input_30_bits_offset_0
    | tryToRead_28[31] & input_31_bits_offset_0;
  assign selectReq_28_bits_vs =
    (tryToRead_28[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_28[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_28[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_28[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_28[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_28[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_28[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_28[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_28[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_28[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_28[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_28[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_28[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_28[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_28[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_28[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_28[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_28[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_28[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_28[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_28[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_28[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_28[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_28[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_28[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_28[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_28[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_28[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_28[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_28[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_28[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_28[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_28_valid =
    tryToRead_28[0] & input_0_valid_0 | tryToRead_28[1] & input_1_valid_0 | tryToRead_28[2] & input_2_valid_0 | tryToRead_28[3] & input_3_valid_0 | tryToRead_28[4] & input_4_valid_0 | tryToRead_28[5] & input_5_valid_0 | tryToRead_28[6]
    & input_6_valid_0 | tryToRead_28[7] & input_7_valid_0 | tryToRead_28[8] & input_8_valid_0 | tryToRead_28[9] & input_9_valid_0 | tryToRead_28[10] & input_10_valid_0 | tryToRead_28[11] & input_11_valid_0 | tryToRead_28[12]
    & input_12_valid_0 | tryToRead_28[13] & input_13_valid_0 | tryToRead_28[14] & input_14_valid_0 | tryToRead_28[15] & input_15_valid_0 | tryToRead_28[16] & input_16_valid_0 | tryToRead_28[17] & input_17_valid_0 | tryToRead_28[18]
    & input_18_valid_0 | tryToRead_28[19] & input_19_valid_0 | tryToRead_28[20] & input_20_valid_0 | tryToRead_28[21] & input_21_valid_0 | tryToRead_28[22] & input_22_valid_0 | tryToRead_28[23] & input_23_valid_0 | tryToRead_28[24]
    & input_24_valid_0 | tryToRead_28[25] & input_25_valid_0 | tryToRead_28[26] & input_26_valid_0 | tryToRead_28[27] & input_27_valid_0 | tryToRead_28[28] & input_28_valid_0 | tryToRead_28[29] & input_29_valid_0 | tryToRead_28[30]
    & input_30_valid_0 | tryToRead_28[31] & input_31_valid_0;
  wire        selectReq_28_ready =
    tryToRead_28[0] & input_0_ready_0 | tryToRead_28[1] & input_1_ready_0 | tryToRead_28[2] & input_2_ready_0 | tryToRead_28[3] & input_3_ready_0 | tryToRead_28[4] & input_4_ready_0 | tryToRead_28[5] & input_5_ready_0 | tryToRead_28[6]
    & input_6_ready_0 | tryToRead_28[7] & input_7_ready_0 | tryToRead_28[8] & input_8_ready_0 | tryToRead_28[9] & input_9_ready_0 | tryToRead_28[10] & input_10_ready_0 | tryToRead_28[11] & input_11_ready_0 | tryToRead_28[12]
    & input_12_ready_0 | tryToRead_28[13] & input_13_ready_0 | tryToRead_28[14] & input_14_ready_0 | tryToRead_28[15] & input_15_ready_0 | tryToRead_28[16] & input_16_ready_0 | tryToRead_28[17] & input_17_ready_0 | tryToRead_28[18]
    & input_18_ready_0 | tryToRead_28[19] & input_19_ready_0 | tryToRead_28[20] & input_20_ready_0 | tryToRead_28[21] & input_21_ready_0 | tryToRead_28[22] & input_22_ready_0 | tryToRead_28[23] & input_23_ready_0 | tryToRead_28[24]
    & input_24_ready_0 | tryToRead_28[25] & input_25_ready_0 | tryToRead_28[26] & input_26_ready_0 | tryToRead_28[27] & input_27_ready_0 | tryToRead_28[28] & input_28_ready_0 | tryToRead_28[29] & input_29_ready_0 | tryToRead_28[30]
    & input_30_ready_0 | tryToRead_28[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_29 = {inputSelect1H_1[29], inputSelect1H_0[29]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_29 = {inputSelect1H_3[29], inputSelect1H_2[29]};
  wire [3:0]  tryToRead_lo_lo_lo_29 = {tryToRead_lo_lo_lo_hi_29, tryToRead_lo_lo_lo_lo_29};
  wire [1:0]  tryToRead_lo_lo_hi_lo_29 = {inputSelect1H_5[29], inputSelect1H_4[29]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_29 = {inputSelect1H_7[29], inputSelect1H_6[29]};
  wire [3:0]  tryToRead_lo_lo_hi_29 = {tryToRead_lo_lo_hi_hi_29, tryToRead_lo_lo_hi_lo_29};
  wire [7:0]  tryToRead_lo_lo_29 = {tryToRead_lo_lo_hi_29, tryToRead_lo_lo_lo_29};
  wire [1:0]  tryToRead_lo_hi_lo_lo_29 = {inputSelect1H_9[29], inputSelect1H_8[29]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_29 = {inputSelect1H_11[29], inputSelect1H_10[29]};
  wire [3:0]  tryToRead_lo_hi_lo_29 = {tryToRead_lo_hi_lo_hi_29, tryToRead_lo_hi_lo_lo_29};
  wire [1:0]  tryToRead_lo_hi_hi_lo_29 = {inputSelect1H_13[29], inputSelect1H_12[29]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_29 = {inputSelect1H_15[29], inputSelect1H_14[29]};
  wire [3:0]  tryToRead_lo_hi_hi_29 = {tryToRead_lo_hi_hi_hi_29, tryToRead_lo_hi_hi_lo_29};
  wire [7:0]  tryToRead_lo_hi_29 = {tryToRead_lo_hi_hi_29, tryToRead_lo_hi_lo_29};
  wire [15:0] tryToRead_lo_29 = {tryToRead_lo_hi_29, tryToRead_lo_lo_29};
  wire [1:0]  tryToRead_hi_lo_lo_lo_29 = {inputSelect1H_17[29], inputSelect1H_16[29]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_29 = {inputSelect1H_19[29], inputSelect1H_18[29]};
  wire [3:0]  tryToRead_hi_lo_lo_29 = {tryToRead_hi_lo_lo_hi_29, tryToRead_hi_lo_lo_lo_29};
  wire [1:0]  tryToRead_hi_lo_hi_lo_29 = {inputSelect1H_21[29], inputSelect1H_20[29]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_29 = {inputSelect1H_23[29], inputSelect1H_22[29]};
  wire [3:0]  tryToRead_hi_lo_hi_29 = {tryToRead_hi_lo_hi_hi_29, tryToRead_hi_lo_hi_lo_29};
  wire [7:0]  tryToRead_hi_lo_29 = {tryToRead_hi_lo_hi_29, tryToRead_hi_lo_lo_29};
  wire [1:0]  tryToRead_hi_hi_lo_lo_29 = {inputSelect1H_25[29], inputSelect1H_24[29]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_29 = {inputSelect1H_27[29], inputSelect1H_26[29]};
  wire [3:0]  tryToRead_hi_hi_lo_29 = {tryToRead_hi_hi_lo_hi_29, tryToRead_hi_hi_lo_lo_29};
  wire [1:0]  tryToRead_hi_hi_hi_lo_29 = {inputSelect1H_29[29], inputSelect1H_28[29]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_29 = {inputSelect1H_31[29], inputSelect1H_30[29]};
  wire [3:0]  tryToRead_hi_hi_hi_29 = {tryToRead_hi_hi_hi_hi_29, tryToRead_hi_hi_hi_lo_29};
  wire [7:0]  tryToRead_hi_hi_29 = {tryToRead_hi_hi_hi_29, tryToRead_hi_hi_lo_29};
  wire [15:0] tryToRead_hi_29 = {tryToRead_hi_hi_29, tryToRead_hi_lo_29};
  wire [31:0] tryToRead_29 = {tryToRead_hi_29, tryToRead_lo_29};
  wire        output_29_valid_0 = |tryToRead_29;
  wire [4:0]  output_29_bits_vs_0 = selectReq_29_bits_vs;
  wire        output_29_bits_offset_0 = selectReq_29_bits_offset;
  wire [4:0]  output_29_bits_writeIndex_0 = selectReq_29_bits_requestIndex;
  wire [1:0]  output_29_bits_dataOffset_0 = selectReq_29_bits_dataOffset;
  assign selectReq_29_bits_dataOffset =
    (tryToRead_29[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_29[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_29[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_29[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_29[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_29[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_29[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_29[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_29[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_29[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_29[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_29[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_29[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_29[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_29[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_29[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_29[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_29[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_29[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_29[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_29[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_29[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_29[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_29[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_29[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_29[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_29_bits_requestIndex =
    {4'h0, tryToRead_29[1]} | {3'h0, tryToRead_29[2], 1'h0} | (tryToRead_29[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_29[4], 2'h0} | (tryToRead_29[5] ? 5'h5 : 5'h0) | (tryToRead_29[6] ? 5'h6 : 5'h0) | (tryToRead_29[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_29[8], 3'h0} | (tryToRead_29[9] ? 5'h9 : 5'h0) | (tryToRead_29[10] ? 5'hA : 5'h0) | (tryToRead_29[11] ? 5'hB : 5'h0) | (tryToRead_29[12] ? 5'hC : 5'h0) | (tryToRead_29[13] ? 5'hD : 5'h0)
    | (tryToRead_29[14] ? 5'hE : 5'h0) | (tryToRead_29[15] ? 5'hF : 5'h0) | {tryToRead_29[16], 4'h0} | (tryToRead_29[17] ? 5'h11 : 5'h0) | (tryToRead_29[18] ? 5'h12 : 5'h0) | (tryToRead_29[19] ? 5'h13 : 5'h0)
    | (tryToRead_29[20] ? 5'h14 : 5'h0) | (tryToRead_29[21] ? 5'h15 : 5'h0) | (tryToRead_29[22] ? 5'h16 : 5'h0) | (tryToRead_29[23] ? 5'h17 : 5'h0) | (tryToRead_29[24] ? 5'h18 : 5'h0) | (tryToRead_29[25] ? 5'h19 : 5'h0)
    | (tryToRead_29[26] ? 5'h1A : 5'h0) | (tryToRead_29[27] ? 5'h1B : 5'h0) | (tryToRead_29[28] ? 5'h1C : 5'h0) | (tryToRead_29[29] ? 5'h1D : 5'h0) | (tryToRead_29[30] ? 5'h1E : 5'h0) | {5{tryToRead_29[31]}};
  wire [4:0]  selectReq_29_bits_readLane =
    (tryToRead_29[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_29[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_29[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_29[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_29[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_29[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_29[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_29[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_29[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_29[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_29[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_29[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_29[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_29[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_29[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_29[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_29[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_29[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_29[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_29[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_29[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_29[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_29[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_29[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_29[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_29[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_29[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_29[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_29[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_29[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_29[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_29[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_29_bits_offset =
    tryToRead_29[0] & input_0_bits_offset_0 | tryToRead_29[1] & input_1_bits_offset_0 | tryToRead_29[2] & input_2_bits_offset_0 | tryToRead_29[3] & input_3_bits_offset_0 | tryToRead_29[4] & input_4_bits_offset_0 | tryToRead_29[5]
    & input_5_bits_offset_0 | tryToRead_29[6] & input_6_bits_offset_0 | tryToRead_29[7] & input_7_bits_offset_0 | tryToRead_29[8] & input_8_bits_offset_0 | tryToRead_29[9] & input_9_bits_offset_0 | tryToRead_29[10] & input_10_bits_offset_0
    | tryToRead_29[11] & input_11_bits_offset_0 | tryToRead_29[12] & input_12_bits_offset_0 | tryToRead_29[13] & input_13_bits_offset_0 | tryToRead_29[14] & input_14_bits_offset_0 | tryToRead_29[15] & input_15_bits_offset_0
    | tryToRead_29[16] & input_16_bits_offset_0 | tryToRead_29[17] & input_17_bits_offset_0 | tryToRead_29[18] & input_18_bits_offset_0 | tryToRead_29[19] & input_19_bits_offset_0 | tryToRead_29[20] & input_20_bits_offset_0
    | tryToRead_29[21] & input_21_bits_offset_0 | tryToRead_29[22] & input_22_bits_offset_0 | tryToRead_29[23] & input_23_bits_offset_0 | tryToRead_29[24] & input_24_bits_offset_0 | tryToRead_29[25] & input_25_bits_offset_0
    | tryToRead_29[26] & input_26_bits_offset_0 | tryToRead_29[27] & input_27_bits_offset_0 | tryToRead_29[28] & input_28_bits_offset_0 | tryToRead_29[29] & input_29_bits_offset_0 | tryToRead_29[30] & input_30_bits_offset_0
    | tryToRead_29[31] & input_31_bits_offset_0;
  assign selectReq_29_bits_vs =
    (tryToRead_29[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_29[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_29[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_29[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_29[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_29[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_29[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_29[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_29[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_29[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_29[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_29[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_29[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_29[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_29[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_29[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_29[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_29[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_29[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_29[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_29[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_29[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_29[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_29[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_29[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_29[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_29[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_29[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_29[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_29[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_29[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_29[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_29_valid =
    tryToRead_29[0] & input_0_valid_0 | tryToRead_29[1] & input_1_valid_0 | tryToRead_29[2] & input_2_valid_0 | tryToRead_29[3] & input_3_valid_0 | tryToRead_29[4] & input_4_valid_0 | tryToRead_29[5] & input_5_valid_0 | tryToRead_29[6]
    & input_6_valid_0 | tryToRead_29[7] & input_7_valid_0 | tryToRead_29[8] & input_8_valid_0 | tryToRead_29[9] & input_9_valid_0 | tryToRead_29[10] & input_10_valid_0 | tryToRead_29[11] & input_11_valid_0 | tryToRead_29[12]
    & input_12_valid_0 | tryToRead_29[13] & input_13_valid_0 | tryToRead_29[14] & input_14_valid_0 | tryToRead_29[15] & input_15_valid_0 | tryToRead_29[16] & input_16_valid_0 | tryToRead_29[17] & input_17_valid_0 | tryToRead_29[18]
    & input_18_valid_0 | tryToRead_29[19] & input_19_valid_0 | tryToRead_29[20] & input_20_valid_0 | tryToRead_29[21] & input_21_valid_0 | tryToRead_29[22] & input_22_valid_0 | tryToRead_29[23] & input_23_valid_0 | tryToRead_29[24]
    & input_24_valid_0 | tryToRead_29[25] & input_25_valid_0 | tryToRead_29[26] & input_26_valid_0 | tryToRead_29[27] & input_27_valid_0 | tryToRead_29[28] & input_28_valid_0 | tryToRead_29[29] & input_29_valid_0 | tryToRead_29[30]
    & input_30_valid_0 | tryToRead_29[31] & input_31_valid_0;
  wire        selectReq_29_ready =
    tryToRead_29[0] & input_0_ready_0 | tryToRead_29[1] & input_1_ready_0 | tryToRead_29[2] & input_2_ready_0 | tryToRead_29[3] & input_3_ready_0 | tryToRead_29[4] & input_4_ready_0 | tryToRead_29[5] & input_5_ready_0 | tryToRead_29[6]
    & input_6_ready_0 | tryToRead_29[7] & input_7_ready_0 | tryToRead_29[8] & input_8_ready_0 | tryToRead_29[9] & input_9_ready_0 | tryToRead_29[10] & input_10_ready_0 | tryToRead_29[11] & input_11_ready_0 | tryToRead_29[12]
    & input_12_ready_0 | tryToRead_29[13] & input_13_ready_0 | tryToRead_29[14] & input_14_ready_0 | tryToRead_29[15] & input_15_ready_0 | tryToRead_29[16] & input_16_ready_0 | tryToRead_29[17] & input_17_ready_0 | tryToRead_29[18]
    & input_18_ready_0 | tryToRead_29[19] & input_19_ready_0 | tryToRead_29[20] & input_20_ready_0 | tryToRead_29[21] & input_21_ready_0 | tryToRead_29[22] & input_22_ready_0 | tryToRead_29[23] & input_23_ready_0 | tryToRead_29[24]
    & input_24_ready_0 | tryToRead_29[25] & input_25_ready_0 | tryToRead_29[26] & input_26_ready_0 | tryToRead_29[27] & input_27_ready_0 | tryToRead_29[28] & input_28_ready_0 | tryToRead_29[29] & input_29_ready_0 | tryToRead_29[30]
    & input_30_ready_0 | tryToRead_29[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_30 = {inputSelect1H_1[30], inputSelect1H_0[30]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_30 = {inputSelect1H_3[30], inputSelect1H_2[30]};
  wire [3:0]  tryToRead_lo_lo_lo_30 = {tryToRead_lo_lo_lo_hi_30, tryToRead_lo_lo_lo_lo_30};
  wire [1:0]  tryToRead_lo_lo_hi_lo_30 = {inputSelect1H_5[30], inputSelect1H_4[30]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_30 = {inputSelect1H_7[30], inputSelect1H_6[30]};
  wire [3:0]  tryToRead_lo_lo_hi_30 = {tryToRead_lo_lo_hi_hi_30, tryToRead_lo_lo_hi_lo_30};
  wire [7:0]  tryToRead_lo_lo_30 = {tryToRead_lo_lo_hi_30, tryToRead_lo_lo_lo_30};
  wire [1:0]  tryToRead_lo_hi_lo_lo_30 = {inputSelect1H_9[30], inputSelect1H_8[30]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_30 = {inputSelect1H_11[30], inputSelect1H_10[30]};
  wire [3:0]  tryToRead_lo_hi_lo_30 = {tryToRead_lo_hi_lo_hi_30, tryToRead_lo_hi_lo_lo_30};
  wire [1:0]  tryToRead_lo_hi_hi_lo_30 = {inputSelect1H_13[30], inputSelect1H_12[30]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_30 = {inputSelect1H_15[30], inputSelect1H_14[30]};
  wire [3:0]  tryToRead_lo_hi_hi_30 = {tryToRead_lo_hi_hi_hi_30, tryToRead_lo_hi_hi_lo_30};
  wire [7:0]  tryToRead_lo_hi_30 = {tryToRead_lo_hi_hi_30, tryToRead_lo_hi_lo_30};
  wire [15:0] tryToRead_lo_30 = {tryToRead_lo_hi_30, tryToRead_lo_lo_30};
  wire [1:0]  tryToRead_hi_lo_lo_lo_30 = {inputSelect1H_17[30], inputSelect1H_16[30]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_30 = {inputSelect1H_19[30], inputSelect1H_18[30]};
  wire [3:0]  tryToRead_hi_lo_lo_30 = {tryToRead_hi_lo_lo_hi_30, tryToRead_hi_lo_lo_lo_30};
  wire [1:0]  tryToRead_hi_lo_hi_lo_30 = {inputSelect1H_21[30], inputSelect1H_20[30]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_30 = {inputSelect1H_23[30], inputSelect1H_22[30]};
  wire [3:0]  tryToRead_hi_lo_hi_30 = {tryToRead_hi_lo_hi_hi_30, tryToRead_hi_lo_hi_lo_30};
  wire [7:0]  tryToRead_hi_lo_30 = {tryToRead_hi_lo_hi_30, tryToRead_hi_lo_lo_30};
  wire [1:0]  tryToRead_hi_hi_lo_lo_30 = {inputSelect1H_25[30], inputSelect1H_24[30]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_30 = {inputSelect1H_27[30], inputSelect1H_26[30]};
  wire [3:0]  tryToRead_hi_hi_lo_30 = {tryToRead_hi_hi_lo_hi_30, tryToRead_hi_hi_lo_lo_30};
  wire [1:0]  tryToRead_hi_hi_hi_lo_30 = {inputSelect1H_29[30], inputSelect1H_28[30]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_30 = {inputSelect1H_31[30], inputSelect1H_30[30]};
  wire [3:0]  tryToRead_hi_hi_hi_30 = {tryToRead_hi_hi_hi_hi_30, tryToRead_hi_hi_hi_lo_30};
  wire [7:0]  tryToRead_hi_hi_30 = {tryToRead_hi_hi_hi_30, tryToRead_hi_hi_lo_30};
  wire [15:0] tryToRead_hi_30 = {tryToRead_hi_hi_30, tryToRead_hi_lo_30};
  wire [31:0] tryToRead_30 = {tryToRead_hi_30, tryToRead_lo_30};
  wire        output_30_valid_0 = |tryToRead_30;
  wire [4:0]  output_30_bits_vs_0 = selectReq_30_bits_vs;
  wire        output_30_bits_offset_0 = selectReq_30_bits_offset;
  wire [4:0]  output_30_bits_writeIndex_0 = selectReq_30_bits_requestIndex;
  wire [1:0]  output_30_bits_dataOffset_0 = selectReq_30_bits_dataOffset;
  assign selectReq_30_bits_dataOffset =
    (tryToRead_30[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_30[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_30[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_30[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_30[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_30[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_30[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_30[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_30[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_30[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_30[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_30[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_30[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_30[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_30[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_30[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_30[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_30[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_30[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_30[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_30[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_30[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_30[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_30[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_30[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_30[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_30_bits_requestIndex =
    {4'h0, tryToRead_30[1]} | {3'h0, tryToRead_30[2], 1'h0} | (tryToRead_30[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_30[4], 2'h0} | (tryToRead_30[5] ? 5'h5 : 5'h0) | (tryToRead_30[6] ? 5'h6 : 5'h0) | (tryToRead_30[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_30[8], 3'h0} | (tryToRead_30[9] ? 5'h9 : 5'h0) | (tryToRead_30[10] ? 5'hA : 5'h0) | (tryToRead_30[11] ? 5'hB : 5'h0) | (tryToRead_30[12] ? 5'hC : 5'h0) | (tryToRead_30[13] ? 5'hD : 5'h0)
    | (tryToRead_30[14] ? 5'hE : 5'h0) | (tryToRead_30[15] ? 5'hF : 5'h0) | {tryToRead_30[16], 4'h0} | (tryToRead_30[17] ? 5'h11 : 5'h0) | (tryToRead_30[18] ? 5'h12 : 5'h0) | (tryToRead_30[19] ? 5'h13 : 5'h0)
    | (tryToRead_30[20] ? 5'h14 : 5'h0) | (tryToRead_30[21] ? 5'h15 : 5'h0) | (tryToRead_30[22] ? 5'h16 : 5'h0) | (tryToRead_30[23] ? 5'h17 : 5'h0) | (tryToRead_30[24] ? 5'h18 : 5'h0) | (tryToRead_30[25] ? 5'h19 : 5'h0)
    | (tryToRead_30[26] ? 5'h1A : 5'h0) | (tryToRead_30[27] ? 5'h1B : 5'h0) | (tryToRead_30[28] ? 5'h1C : 5'h0) | (tryToRead_30[29] ? 5'h1D : 5'h0) | (tryToRead_30[30] ? 5'h1E : 5'h0) | {5{tryToRead_30[31]}};
  wire [4:0]  selectReq_30_bits_readLane =
    (tryToRead_30[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_30[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_30[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_30[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_30[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_30[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_30[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_30[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_30[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_30[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_30[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_30[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_30[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_30[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_30[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_30[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_30[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_30[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_30[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_30[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_30[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_30[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_30[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_30[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_30[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_30[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_30[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_30[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_30[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_30[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_30[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_30[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_30_bits_offset =
    tryToRead_30[0] & input_0_bits_offset_0 | tryToRead_30[1] & input_1_bits_offset_0 | tryToRead_30[2] & input_2_bits_offset_0 | tryToRead_30[3] & input_3_bits_offset_0 | tryToRead_30[4] & input_4_bits_offset_0 | tryToRead_30[5]
    & input_5_bits_offset_0 | tryToRead_30[6] & input_6_bits_offset_0 | tryToRead_30[7] & input_7_bits_offset_0 | tryToRead_30[8] & input_8_bits_offset_0 | tryToRead_30[9] & input_9_bits_offset_0 | tryToRead_30[10] & input_10_bits_offset_0
    | tryToRead_30[11] & input_11_bits_offset_0 | tryToRead_30[12] & input_12_bits_offset_0 | tryToRead_30[13] & input_13_bits_offset_0 | tryToRead_30[14] & input_14_bits_offset_0 | tryToRead_30[15] & input_15_bits_offset_0
    | tryToRead_30[16] & input_16_bits_offset_0 | tryToRead_30[17] & input_17_bits_offset_0 | tryToRead_30[18] & input_18_bits_offset_0 | tryToRead_30[19] & input_19_bits_offset_0 | tryToRead_30[20] & input_20_bits_offset_0
    | tryToRead_30[21] & input_21_bits_offset_0 | tryToRead_30[22] & input_22_bits_offset_0 | tryToRead_30[23] & input_23_bits_offset_0 | tryToRead_30[24] & input_24_bits_offset_0 | tryToRead_30[25] & input_25_bits_offset_0
    | tryToRead_30[26] & input_26_bits_offset_0 | tryToRead_30[27] & input_27_bits_offset_0 | tryToRead_30[28] & input_28_bits_offset_0 | tryToRead_30[29] & input_29_bits_offset_0 | tryToRead_30[30] & input_30_bits_offset_0
    | tryToRead_30[31] & input_31_bits_offset_0;
  assign selectReq_30_bits_vs =
    (tryToRead_30[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_30[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_30[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_30[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_30[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_30[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_30[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_30[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_30[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_30[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_30[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_30[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_30[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_30[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_30[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_30[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_30[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_30[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_30[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_30[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_30[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_30[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_30[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_30[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_30[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_30[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_30[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_30[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_30[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_30[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_30[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_30[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_30_valid =
    tryToRead_30[0] & input_0_valid_0 | tryToRead_30[1] & input_1_valid_0 | tryToRead_30[2] & input_2_valid_0 | tryToRead_30[3] & input_3_valid_0 | tryToRead_30[4] & input_4_valid_0 | tryToRead_30[5] & input_5_valid_0 | tryToRead_30[6]
    & input_6_valid_0 | tryToRead_30[7] & input_7_valid_0 | tryToRead_30[8] & input_8_valid_0 | tryToRead_30[9] & input_9_valid_0 | tryToRead_30[10] & input_10_valid_0 | tryToRead_30[11] & input_11_valid_0 | tryToRead_30[12]
    & input_12_valid_0 | tryToRead_30[13] & input_13_valid_0 | tryToRead_30[14] & input_14_valid_0 | tryToRead_30[15] & input_15_valid_0 | tryToRead_30[16] & input_16_valid_0 | tryToRead_30[17] & input_17_valid_0 | tryToRead_30[18]
    & input_18_valid_0 | tryToRead_30[19] & input_19_valid_0 | tryToRead_30[20] & input_20_valid_0 | tryToRead_30[21] & input_21_valid_0 | tryToRead_30[22] & input_22_valid_0 | tryToRead_30[23] & input_23_valid_0 | tryToRead_30[24]
    & input_24_valid_0 | tryToRead_30[25] & input_25_valid_0 | tryToRead_30[26] & input_26_valid_0 | tryToRead_30[27] & input_27_valid_0 | tryToRead_30[28] & input_28_valid_0 | tryToRead_30[29] & input_29_valid_0 | tryToRead_30[30]
    & input_30_valid_0 | tryToRead_30[31] & input_31_valid_0;
  wire        selectReq_30_ready =
    tryToRead_30[0] & input_0_ready_0 | tryToRead_30[1] & input_1_ready_0 | tryToRead_30[2] & input_2_ready_0 | tryToRead_30[3] & input_3_ready_0 | tryToRead_30[4] & input_4_ready_0 | tryToRead_30[5] & input_5_ready_0 | tryToRead_30[6]
    & input_6_ready_0 | tryToRead_30[7] & input_7_ready_0 | tryToRead_30[8] & input_8_ready_0 | tryToRead_30[9] & input_9_ready_0 | tryToRead_30[10] & input_10_ready_0 | tryToRead_30[11] & input_11_ready_0 | tryToRead_30[12]
    & input_12_ready_0 | tryToRead_30[13] & input_13_ready_0 | tryToRead_30[14] & input_14_ready_0 | tryToRead_30[15] & input_15_ready_0 | tryToRead_30[16] & input_16_ready_0 | tryToRead_30[17] & input_17_ready_0 | tryToRead_30[18]
    & input_18_ready_0 | tryToRead_30[19] & input_19_ready_0 | tryToRead_30[20] & input_20_ready_0 | tryToRead_30[21] & input_21_ready_0 | tryToRead_30[22] & input_22_ready_0 | tryToRead_30[23] & input_23_ready_0 | tryToRead_30[24]
    & input_24_ready_0 | tryToRead_30[25] & input_25_ready_0 | tryToRead_30[26] & input_26_ready_0 | tryToRead_30[27] & input_27_ready_0 | tryToRead_30[28] & input_28_ready_0 | tryToRead_30[29] & input_29_ready_0 | tryToRead_30[30]
    & input_30_ready_0 | tryToRead_30[31] & input_31_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_lo_31 = {inputSelect1H_1[31], inputSelect1H_0[31]};
  wire [1:0]  tryToRead_lo_lo_lo_hi_31 = {inputSelect1H_3[31], inputSelect1H_2[31]};
  wire [3:0]  tryToRead_lo_lo_lo_31 = {tryToRead_lo_lo_lo_hi_31, tryToRead_lo_lo_lo_lo_31};
  wire [1:0]  tryToRead_lo_lo_hi_lo_31 = {inputSelect1H_5[31], inputSelect1H_4[31]};
  wire [1:0]  tryToRead_lo_lo_hi_hi_31 = {inputSelect1H_7[31], inputSelect1H_6[31]};
  wire [3:0]  tryToRead_lo_lo_hi_31 = {tryToRead_lo_lo_hi_hi_31, tryToRead_lo_lo_hi_lo_31};
  wire [7:0]  tryToRead_lo_lo_31 = {tryToRead_lo_lo_hi_31, tryToRead_lo_lo_lo_31};
  wire [1:0]  tryToRead_lo_hi_lo_lo_31 = {inputSelect1H_9[31], inputSelect1H_8[31]};
  wire [1:0]  tryToRead_lo_hi_lo_hi_31 = {inputSelect1H_11[31], inputSelect1H_10[31]};
  wire [3:0]  tryToRead_lo_hi_lo_31 = {tryToRead_lo_hi_lo_hi_31, tryToRead_lo_hi_lo_lo_31};
  wire [1:0]  tryToRead_lo_hi_hi_lo_31 = {inputSelect1H_13[31], inputSelect1H_12[31]};
  wire [1:0]  tryToRead_lo_hi_hi_hi_31 = {inputSelect1H_15[31], inputSelect1H_14[31]};
  wire [3:0]  tryToRead_lo_hi_hi_31 = {tryToRead_lo_hi_hi_hi_31, tryToRead_lo_hi_hi_lo_31};
  wire [7:0]  tryToRead_lo_hi_31 = {tryToRead_lo_hi_hi_31, tryToRead_lo_hi_lo_31};
  wire [15:0] tryToRead_lo_31 = {tryToRead_lo_hi_31, tryToRead_lo_lo_31};
  wire [1:0]  tryToRead_hi_lo_lo_lo_31 = {inputSelect1H_17[31], inputSelect1H_16[31]};
  wire [1:0]  tryToRead_hi_lo_lo_hi_31 = {inputSelect1H_19[31], inputSelect1H_18[31]};
  wire [3:0]  tryToRead_hi_lo_lo_31 = {tryToRead_hi_lo_lo_hi_31, tryToRead_hi_lo_lo_lo_31};
  wire [1:0]  tryToRead_hi_lo_hi_lo_31 = {inputSelect1H_21[31], inputSelect1H_20[31]};
  wire [1:0]  tryToRead_hi_lo_hi_hi_31 = {inputSelect1H_23[31], inputSelect1H_22[31]};
  wire [3:0]  tryToRead_hi_lo_hi_31 = {tryToRead_hi_lo_hi_hi_31, tryToRead_hi_lo_hi_lo_31};
  wire [7:0]  tryToRead_hi_lo_31 = {tryToRead_hi_lo_hi_31, tryToRead_hi_lo_lo_31};
  wire [1:0]  tryToRead_hi_hi_lo_lo_31 = {inputSelect1H_25[31], inputSelect1H_24[31]};
  wire [1:0]  tryToRead_hi_hi_lo_hi_31 = {inputSelect1H_27[31], inputSelect1H_26[31]};
  wire [3:0]  tryToRead_hi_hi_lo_31 = {tryToRead_hi_hi_lo_hi_31, tryToRead_hi_hi_lo_lo_31};
  wire [1:0]  tryToRead_hi_hi_hi_lo_31 = {inputSelect1H_29[31], inputSelect1H_28[31]};
  wire [1:0]  tryToRead_hi_hi_hi_hi_31 = {inputSelect1H_31[31], inputSelect1H_30[31]};
  wire [3:0]  tryToRead_hi_hi_hi_31 = {tryToRead_hi_hi_hi_hi_31, tryToRead_hi_hi_hi_lo_31};
  wire [7:0]  tryToRead_hi_hi_31 = {tryToRead_hi_hi_hi_31, tryToRead_hi_hi_lo_31};
  wire [15:0] tryToRead_hi_31 = {tryToRead_hi_hi_31, tryToRead_hi_lo_31};
  wire [31:0] tryToRead_31 = {tryToRead_hi_31, tryToRead_lo_31};
  wire        output_31_valid_0 = |tryToRead_31;
  wire [4:0]  output_31_bits_vs_0 = selectReq_31_bits_vs;
  wire        output_31_bits_offset_0 = selectReq_31_bits_offset;
  wire [4:0]  output_31_bits_writeIndex_0 = selectReq_31_bits_requestIndex;
  wire [1:0]  output_31_bits_dataOffset_0 = selectReq_31_bits_dataOffset;
  assign selectReq_31_bits_dataOffset =
    (tryToRead_31[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_31[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_31[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_31[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_31[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_31[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_31[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_31[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_31[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_31[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_31[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_31[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_31[15] ? input_15_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[16] ? input_16_bits_dataOffset_0 : 2'h0) | (tryToRead_31[17] ? input_17_bits_dataOffset_0 : 2'h0) | (tryToRead_31[18] ? input_18_bits_dataOffset_0 : 2'h0) | (tryToRead_31[19] ? input_19_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[20] ? input_20_bits_dataOffset_0 : 2'h0) | (tryToRead_31[21] ? input_21_bits_dataOffset_0 : 2'h0) | (tryToRead_31[22] ? input_22_bits_dataOffset_0 : 2'h0) | (tryToRead_31[23] ? input_23_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[24] ? input_24_bits_dataOffset_0 : 2'h0) | (tryToRead_31[25] ? input_25_bits_dataOffset_0 : 2'h0) | (tryToRead_31[26] ? input_26_bits_dataOffset_0 : 2'h0) | (tryToRead_31[27] ? input_27_bits_dataOffset_0 : 2'h0)
    | (tryToRead_31[28] ? input_28_bits_dataOffset_0 : 2'h0) | (tryToRead_31[29] ? input_29_bits_dataOffset_0 : 2'h0) | (tryToRead_31[30] ? input_30_bits_dataOffset_0 : 2'h0) | (tryToRead_31[31] ? input_31_bits_dataOffset_0 : 2'h0);
  assign selectReq_31_bits_requestIndex =
    {4'h0, tryToRead_31[1]} | {3'h0, tryToRead_31[2], 1'h0} | (tryToRead_31[3] ? 5'h3 : 5'h0) | {2'h0, tryToRead_31[4], 2'h0} | (tryToRead_31[5] ? 5'h5 : 5'h0) | (tryToRead_31[6] ? 5'h6 : 5'h0) | (tryToRead_31[7] ? 5'h7 : 5'h0)
    | {1'h0, tryToRead_31[8], 3'h0} | (tryToRead_31[9] ? 5'h9 : 5'h0) | (tryToRead_31[10] ? 5'hA : 5'h0) | (tryToRead_31[11] ? 5'hB : 5'h0) | (tryToRead_31[12] ? 5'hC : 5'h0) | (tryToRead_31[13] ? 5'hD : 5'h0)
    | (tryToRead_31[14] ? 5'hE : 5'h0) | (tryToRead_31[15] ? 5'hF : 5'h0) | {tryToRead_31[16], 4'h0} | (tryToRead_31[17] ? 5'h11 : 5'h0) | (tryToRead_31[18] ? 5'h12 : 5'h0) | (tryToRead_31[19] ? 5'h13 : 5'h0)
    | (tryToRead_31[20] ? 5'h14 : 5'h0) | (tryToRead_31[21] ? 5'h15 : 5'h0) | (tryToRead_31[22] ? 5'h16 : 5'h0) | (tryToRead_31[23] ? 5'h17 : 5'h0) | (tryToRead_31[24] ? 5'h18 : 5'h0) | (tryToRead_31[25] ? 5'h19 : 5'h0)
    | (tryToRead_31[26] ? 5'h1A : 5'h0) | (tryToRead_31[27] ? 5'h1B : 5'h0) | (tryToRead_31[28] ? 5'h1C : 5'h0) | (tryToRead_31[29] ? 5'h1D : 5'h0) | (tryToRead_31[30] ? 5'h1E : 5'h0) | {5{tryToRead_31[31]}};
  wire [4:0]  selectReq_31_bits_readLane =
    (tryToRead_31[0] ? input_0_bits_readLane_0 : 5'h0) | (tryToRead_31[1] ? input_1_bits_readLane_0 : 5'h0) | (tryToRead_31[2] ? input_2_bits_readLane_0 : 5'h0) | (tryToRead_31[3] ? input_3_bits_readLane_0 : 5'h0)
    | (tryToRead_31[4] ? input_4_bits_readLane_0 : 5'h0) | (tryToRead_31[5] ? input_5_bits_readLane_0 : 5'h0) | (tryToRead_31[6] ? input_6_bits_readLane_0 : 5'h0) | (tryToRead_31[7] ? input_7_bits_readLane_0 : 5'h0)
    | (tryToRead_31[8] ? input_8_bits_readLane_0 : 5'h0) | (tryToRead_31[9] ? input_9_bits_readLane_0 : 5'h0) | (tryToRead_31[10] ? input_10_bits_readLane_0 : 5'h0) | (tryToRead_31[11] ? input_11_bits_readLane_0 : 5'h0)
    | (tryToRead_31[12] ? input_12_bits_readLane_0 : 5'h0) | (tryToRead_31[13] ? input_13_bits_readLane_0 : 5'h0) | (tryToRead_31[14] ? input_14_bits_readLane_0 : 5'h0) | (tryToRead_31[15] ? input_15_bits_readLane_0 : 5'h0)
    | (tryToRead_31[16] ? input_16_bits_readLane_0 : 5'h0) | (tryToRead_31[17] ? input_17_bits_readLane_0 : 5'h0) | (tryToRead_31[18] ? input_18_bits_readLane_0 : 5'h0) | (tryToRead_31[19] ? input_19_bits_readLane_0 : 5'h0)
    | (tryToRead_31[20] ? input_20_bits_readLane_0 : 5'h0) | (tryToRead_31[21] ? input_21_bits_readLane_0 : 5'h0) | (tryToRead_31[22] ? input_22_bits_readLane_0 : 5'h0) | (tryToRead_31[23] ? input_23_bits_readLane_0 : 5'h0)
    | (tryToRead_31[24] ? input_24_bits_readLane_0 : 5'h0) | (tryToRead_31[25] ? input_25_bits_readLane_0 : 5'h0) | (tryToRead_31[26] ? input_26_bits_readLane_0 : 5'h0) | (tryToRead_31[27] ? input_27_bits_readLane_0 : 5'h0)
    | (tryToRead_31[28] ? input_28_bits_readLane_0 : 5'h0) | (tryToRead_31[29] ? input_29_bits_readLane_0 : 5'h0) | (tryToRead_31[30] ? input_30_bits_readLane_0 : 5'h0) | (tryToRead_31[31] ? input_31_bits_readLane_0 : 5'h0);
  assign selectReq_31_bits_offset =
    tryToRead_31[0] & input_0_bits_offset_0 | tryToRead_31[1] & input_1_bits_offset_0 | tryToRead_31[2] & input_2_bits_offset_0 | tryToRead_31[3] & input_3_bits_offset_0 | tryToRead_31[4] & input_4_bits_offset_0 | tryToRead_31[5]
    & input_5_bits_offset_0 | tryToRead_31[6] & input_6_bits_offset_0 | tryToRead_31[7] & input_7_bits_offset_0 | tryToRead_31[8] & input_8_bits_offset_0 | tryToRead_31[9] & input_9_bits_offset_0 | tryToRead_31[10] & input_10_bits_offset_0
    | tryToRead_31[11] & input_11_bits_offset_0 | tryToRead_31[12] & input_12_bits_offset_0 | tryToRead_31[13] & input_13_bits_offset_0 | tryToRead_31[14] & input_14_bits_offset_0 | tryToRead_31[15] & input_15_bits_offset_0
    | tryToRead_31[16] & input_16_bits_offset_0 | tryToRead_31[17] & input_17_bits_offset_0 | tryToRead_31[18] & input_18_bits_offset_0 | tryToRead_31[19] & input_19_bits_offset_0 | tryToRead_31[20] & input_20_bits_offset_0
    | tryToRead_31[21] & input_21_bits_offset_0 | tryToRead_31[22] & input_22_bits_offset_0 | tryToRead_31[23] & input_23_bits_offset_0 | tryToRead_31[24] & input_24_bits_offset_0 | tryToRead_31[25] & input_25_bits_offset_0
    | tryToRead_31[26] & input_26_bits_offset_0 | tryToRead_31[27] & input_27_bits_offset_0 | tryToRead_31[28] & input_28_bits_offset_0 | tryToRead_31[29] & input_29_bits_offset_0 | tryToRead_31[30] & input_30_bits_offset_0
    | tryToRead_31[31] & input_31_bits_offset_0;
  assign selectReq_31_bits_vs =
    (tryToRead_31[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_31[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_31[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_31[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_31[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_31[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_31[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_31[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_31[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_31[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_31[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_31[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_31[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_31[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_31[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_31[15] ? input_15_bits_vs_0 : 5'h0) | (tryToRead_31[16] ? input_16_bits_vs_0 : 5'h0) | (tryToRead_31[17] ? input_17_bits_vs_0 : 5'h0)
    | (tryToRead_31[18] ? input_18_bits_vs_0 : 5'h0) | (tryToRead_31[19] ? input_19_bits_vs_0 : 5'h0) | (tryToRead_31[20] ? input_20_bits_vs_0 : 5'h0) | (tryToRead_31[21] ? input_21_bits_vs_0 : 5'h0)
    | (tryToRead_31[22] ? input_22_bits_vs_0 : 5'h0) | (tryToRead_31[23] ? input_23_bits_vs_0 : 5'h0) | (tryToRead_31[24] ? input_24_bits_vs_0 : 5'h0) | (tryToRead_31[25] ? input_25_bits_vs_0 : 5'h0)
    | (tryToRead_31[26] ? input_26_bits_vs_0 : 5'h0) | (tryToRead_31[27] ? input_27_bits_vs_0 : 5'h0) | (tryToRead_31[28] ? input_28_bits_vs_0 : 5'h0) | (tryToRead_31[29] ? input_29_bits_vs_0 : 5'h0)
    | (tryToRead_31[30] ? input_30_bits_vs_0 : 5'h0) | (tryToRead_31[31] ? input_31_bits_vs_0 : 5'h0);
  wire        selectReq_31_valid =
    tryToRead_31[0] & input_0_valid_0 | tryToRead_31[1] & input_1_valid_0 | tryToRead_31[2] & input_2_valid_0 | tryToRead_31[3] & input_3_valid_0 | tryToRead_31[4] & input_4_valid_0 | tryToRead_31[5] & input_5_valid_0 | tryToRead_31[6]
    & input_6_valid_0 | tryToRead_31[7] & input_7_valid_0 | tryToRead_31[8] & input_8_valid_0 | tryToRead_31[9] & input_9_valid_0 | tryToRead_31[10] & input_10_valid_0 | tryToRead_31[11] & input_11_valid_0 | tryToRead_31[12]
    & input_12_valid_0 | tryToRead_31[13] & input_13_valid_0 | tryToRead_31[14] & input_14_valid_0 | tryToRead_31[15] & input_15_valid_0 | tryToRead_31[16] & input_16_valid_0 | tryToRead_31[17] & input_17_valid_0 | tryToRead_31[18]
    & input_18_valid_0 | tryToRead_31[19] & input_19_valid_0 | tryToRead_31[20] & input_20_valid_0 | tryToRead_31[21] & input_21_valid_0 | tryToRead_31[22] & input_22_valid_0 | tryToRead_31[23] & input_23_valid_0 | tryToRead_31[24]
    & input_24_valid_0 | tryToRead_31[25] & input_25_valid_0 | tryToRead_31[26] & input_26_valid_0 | tryToRead_31[27] & input_27_valid_0 | tryToRead_31[28] & input_28_valid_0 | tryToRead_31[29] & input_29_valid_0 | tryToRead_31[30]
    & input_30_valid_0 | tryToRead_31[31] & input_31_valid_0;
  wire        selectReq_31_ready =
    tryToRead_31[0] & input_0_ready_0 | tryToRead_31[1] & input_1_ready_0 | tryToRead_31[2] & input_2_ready_0 | tryToRead_31[3] & input_3_ready_0 | tryToRead_31[4] & input_4_ready_0 | tryToRead_31[5] & input_5_ready_0 | tryToRead_31[6]
    & input_6_ready_0 | tryToRead_31[7] & input_7_ready_0 | tryToRead_31[8] & input_8_ready_0 | tryToRead_31[9] & input_9_ready_0 | tryToRead_31[10] & input_10_ready_0 | tryToRead_31[11] & input_11_ready_0 | tryToRead_31[12]
    & input_12_ready_0 | tryToRead_31[13] & input_13_ready_0 | tryToRead_31[14] & input_14_ready_0 | tryToRead_31[15] & input_15_ready_0 | tryToRead_31[16] & input_16_ready_0 | tryToRead_31[17] & input_17_ready_0 | tryToRead_31[18]
    & input_18_ready_0 | tryToRead_31[19] & input_19_ready_0 | tryToRead_31[20] & input_20_ready_0 | tryToRead_31[21] & input_21_ready_0 | tryToRead_31[22] & input_22_ready_0 | tryToRead_31[23] & input_23_ready_0 | tryToRead_31[24]
    & input_24_ready_0 | tryToRead_31[25] & input_25_ready_0 | tryToRead_31[26] & input_26_ready_0 | tryToRead_31[27] & input_27_ready_0 | tryToRead_31[28] & input_28_ready_0 | tryToRead_31[29] & input_29_ready_0 | tryToRead_31[30]
    & input_30_ready_0 | tryToRead_31[31] & input_31_ready_0;
  assign input_0_ready = input_0_ready_0;
  assign input_1_ready = input_1_ready_0;
  assign input_2_ready = input_2_ready_0;
  assign input_3_ready = input_3_ready_0;
  assign input_4_ready = input_4_ready_0;
  assign input_5_ready = input_5_ready_0;
  assign input_6_ready = input_6_ready_0;
  assign input_7_ready = input_7_ready_0;
  assign input_8_ready = input_8_ready_0;
  assign input_9_ready = input_9_ready_0;
  assign input_10_ready = input_10_ready_0;
  assign input_11_ready = input_11_ready_0;
  assign input_12_ready = input_12_ready_0;
  assign input_13_ready = input_13_ready_0;
  assign input_14_ready = input_14_ready_0;
  assign input_15_ready = input_15_ready_0;
  assign input_16_ready = input_16_ready_0;
  assign input_17_ready = input_17_ready_0;
  assign input_18_ready = input_18_ready_0;
  assign input_19_ready = input_19_ready_0;
  assign input_20_ready = input_20_ready_0;
  assign input_21_ready = input_21_ready_0;
  assign input_22_ready = input_22_ready_0;
  assign input_23_ready = input_23_ready_0;
  assign input_24_ready = input_24_ready_0;
  assign input_25_ready = input_25_ready_0;
  assign input_26_ready = input_26_ready_0;
  assign input_27_ready = input_27_ready_0;
  assign input_28_ready = input_28_ready_0;
  assign input_29_ready = input_29_ready_0;
  assign input_30_ready = input_30_ready_0;
  assign input_31_ready = input_31_ready_0;
  assign output_0_valid = output_0_valid_0;
  assign output_0_bits_vs = output_0_bits_vs_0;
  assign output_0_bits_offset = output_0_bits_offset_0;
  assign output_0_bits_writeIndex = output_0_bits_writeIndex_0;
  assign output_0_bits_dataOffset = output_0_bits_dataOffset_0;
  assign output_1_valid = output_1_valid_0;
  assign output_1_bits_vs = output_1_bits_vs_0;
  assign output_1_bits_offset = output_1_bits_offset_0;
  assign output_1_bits_writeIndex = output_1_bits_writeIndex_0;
  assign output_1_bits_dataOffset = output_1_bits_dataOffset_0;
  assign output_2_valid = output_2_valid_0;
  assign output_2_bits_vs = output_2_bits_vs_0;
  assign output_2_bits_offset = output_2_bits_offset_0;
  assign output_2_bits_writeIndex = output_2_bits_writeIndex_0;
  assign output_2_bits_dataOffset = output_2_bits_dataOffset_0;
  assign output_3_valid = output_3_valid_0;
  assign output_3_bits_vs = output_3_bits_vs_0;
  assign output_3_bits_offset = output_3_bits_offset_0;
  assign output_3_bits_writeIndex = output_3_bits_writeIndex_0;
  assign output_3_bits_dataOffset = output_3_bits_dataOffset_0;
  assign output_4_valid = output_4_valid_0;
  assign output_4_bits_vs = output_4_bits_vs_0;
  assign output_4_bits_offset = output_4_bits_offset_0;
  assign output_4_bits_writeIndex = output_4_bits_writeIndex_0;
  assign output_4_bits_dataOffset = output_4_bits_dataOffset_0;
  assign output_5_valid = output_5_valid_0;
  assign output_5_bits_vs = output_5_bits_vs_0;
  assign output_5_bits_offset = output_5_bits_offset_0;
  assign output_5_bits_writeIndex = output_5_bits_writeIndex_0;
  assign output_5_bits_dataOffset = output_5_bits_dataOffset_0;
  assign output_6_valid = output_6_valid_0;
  assign output_6_bits_vs = output_6_bits_vs_0;
  assign output_6_bits_offset = output_6_bits_offset_0;
  assign output_6_bits_writeIndex = output_6_bits_writeIndex_0;
  assign output_6_bits_dataOffset = output_6_bits_dataOffset_0;
  assign output_7_valid = output_7_valid_0;
  assign output_7_bits_vs = output_7_bits_vs_0;
  assign output_7_bits_offset = output_7_bits_offset_0;
  assign output_7_bits_writeIndex = output_7_bits_writeIndex_0;
  assign output_7_bits_dataOffset = output_7_bits_dataOffset_0;
  assign output_8_valid = output_8_valid_0;
  assign output_8_bits_vs = output_8_bits_vs_0;
  assign output_8_bits_offset = output_8_bits_offset_0;
  assign output_8_bits_writeIndex = output_8_bits_writeIndex_0;
  assign output_8_bits_dataOffset = output_8_bits_dataOffset_0;
  assign output_9_valid = output_9_valid_0;
  assign output_9_bits_vs = output_9_bits_vs_0;
  assign output_9_bits_offset = output_9_bits_offset_0;
  assign output_9_bits_writeIndex = output_9_bits_writeIndex_0;
  assign output_9_bits_dataOffset = output_9_bits_dataOffset_0;
  assign output_10_valid = output_10_valid_0;
  assign output_10_bits_vs = output_10_bits_vs_0;
  assign output_10_bits_offset = output_10_bits_offset_0;
  assign output_10_bits_writeIndex = output_10_bits_writeIndex_0;
  assign output_10_bits_dataOffset = output_10_bits_dataOffset_0;
  assign output_11_valid = output_11_valid_0;
  assign output_11_bits_vs = output_11_bits_vs_0;
  assign output_11_bits_offset = output_11_bits_offset_0;
  assign output_11_bits_writeIndex = output_11_bits_writeIndex_0;
  assign output_11_bits_dataOffset = output_11_bits_dataOffset_0;
  assign output_12_valid = output_12_valid_0;
  assign output_12_bits_vs = output_12_bits_vs_0;
  assign output_12_bits_offset = output_12_bits_offset_0;
  assign output_12_bits_writeIndex = output_12_bits_writeIndex_0;
  assign output_12_bits_dataOffset = output_12_bits_dataOffset_0;
  assign output_13_valid = output_13_valid_0;
  assign output_13_bits_vs = output_13_bits_vs_0;
  assign output_13_bits_offset = output_13_bits_offset_0;
  assign output_13_bits_writeIndex = output_13_bits_writeIndex_0;
  assign output_13_bits_dataOffset = output_13_bits_dataOffset_0;
  assign output_14_valid = output_14_valid_0;
  assign output_14_bits_vs = output_14_bits_vs_0;
  assign output_14_bits_offset = output_14_bits_offset_0;
  assign output_14_bits_writeIndex = output_14_bits_writeIndex_0;
  assign output_14_bits_dataOffset = output_14_bits_dataOffset_0;
  assign output_15_valid = output_15_valid_0;
  assign output_15_bits_vs = output_15_bits_vs_0;
  assign output_15_bits_offset = output_15_bits_offset_0;
  assign output_15_bits_writeIndex = output_15_bits_writeIndex_0;
  assign output_15_bits_dataOffset = output_15_bits_dataOffset_0;
  assign output_16_valid = output_16_valid_0;
  assign output_16_bits_vs = output_16_bits_vs_0;
  assign output_16_bits_offset = output_16_bits_offset_0;
  assign output_16_bits_writeIndex = output_16_bits_writeIndex_0;
  assign output_16_bits_dataOffset = output_16_bits_dataOffset_0;
  assign output_17_valid = output_17_valid_0;
  assign output_17_bits_vs = output_17_bits_vs_0;
  assign output_17_bits_offset = output_17_bits_offset_0;
  assign output_17_bits_writeIndex = output_17_bits_writeIndex_0;
  assign output_17_bits_dataOffset = output_17_bits_dataOffset_0;
  assign output_18_valid = output_18_valid_0;
  assign output_18_bits_vs = output_18_bits_vs_0;
  assign output_18_bits_offset = output_18_bits_offset_0;
  assign output_18_bits_writeIndex = output_18_bits_writeIndex_0;
  assign output_18_bits_dataOffset = output_18_bits_dataOffset_0;
  assign output_19_valid = output_19_valid_0;
  assign output_19_bits_vs = output_19_bits_vs_0;
  assign output_19_bits_offset = output_19_bits_offset_0;
  assign output_19_bits_writeIndex = output_19_bits_writeIndex_0;
  assign output_19_bits_dataOffset = output_19_bits_dataOffset_0;
  assign output_20_valid = output_20_valid_0;
  assign output_20_bits_vs = output_20_bits_vs_0;
  assign output_20_bits_offset = output_20_bits_offset_0;
  assign output_20_bits_writeIndex = output_20_bits_writeIndex_0;
  assign output_20_bits_dataOffset = output_20_bits_dataOffset_0;
  assign output_21_valid = output_21_valid_0;
  assign output_21_bits_vs = output_21_bits_vs_0;
  assign output_21_bits_offset = output_21_bits_offset_0;
  assign output_21_bits_writeIndex = output_21_bits_writeIndex_0;
  assign output_21_bits_dataOffset = output_21_bits_dataOffset_0;
  assign output_22_valid = output_22_valid_0;
  assign output_22_bits_vs = output_22_bits_vs_0;
  assign output_22_bits_offset = output_22_bits_offset_0;
  assign output_22_bits_writeIndex = output_22_bits_writeIndex_0;
  assign output_22_bits_dataOffset = output_22_bits_dataOffset_0;
  assign output_23_valid = output_23_valid_0;
  assign output_23_bits_vs = output_23_bits_vs_0;
  assign output_23_bits_offset = output_23_bits_offset_0;
  assign output_23_bits_writeIndex = output_23_bits_writeIndex_0;
  assign output_23_bits_dataOffset = output_23_bits_dataOffset_0;
  assign output_24_valid = output_24_valid_0;
  assign output_24_bits_vs = output_24_bits_vs_0;
  assign output_24_bits_offset = output_24_bits_offset_0;
  assign output_24_bits_writeIndex = output_24_bits_writeIndex_0;
  assign output_24_bits_dataOffset = output_24_bits_dataOffset_0;
  assign output_25_valid = output_25_valid_0;
  assign output_25_bits_vs = output_25_bits_vs_0;
  assign output_25_bits_offset = output_25_bits_offset_0;
  assign output_25_bits_writeIndex = output_25_bits_writeIndex_0;
  assign output_25_bits_dataOffset = output_25_bits_dataOffset_0;
  assign output_26_valid = output_26_valid_0;
  assign output_26_bits_vs = output_26_bits_vs_0;
  assign output_26_bits_offset = output_26_bits_offset_0;
  assign output_26_bits_writeIndex = output_26_bits_writeIndex_0;
  assign output_26_bits_dataOffset = output_26_bits_dataOffset_0;
  assign output_27_valid = output_27_valid_0;
  assign output_27_bits_vs = output_27_bits_vs_0;
  assign output_27_bits_offset = output_27_bits_offset_0;
  assign output_27_bits_writeIndex = output_27_bits_writeIndex_0;
  assign output_27_bits_dataOffset = output_27_bits_dataOffset_0;
  assign output_28_valid = output_28_valid_0;
  assign output_28_bits_vs = output_28_bits_vs_0;
  assign output_28_bits_offset = output_28_bits_offset_0;
  assign output_28_bits_writeIndex = output_28_bits_writeIndex_0;
  assign output_28_bits_dataOffset = output_28_bits_dataOffset_0;
  assign output_29_valid = output_29_valid_0;
  assign output_29_bits_vs = output_29_bits_vs_0;
  assign output_29_bits_offset = output_29_bits_offset_0;
  assign output_29_bits_writeIndex = output_29_bits_writeIndex_0;
  assign output_29_bits_dataOffset = output_29_bits_dataOffset_0;
  assign output_30_valid = output_30_valid_0;
  assign output_30_bits_vs = output_30_bits_vs_0;
  assign output_30_bits_offset = output_30_bits_offset_0;
  assign output_30_bits_writeIndex = output_30_bits_writeIndex_0;
  assign output_30_bits_dataOffset = output_30_bits_dataOffset_0;
  assign output_31_valid = output_31_valid_0;
  assign output_31_bits_vs = output_31_bits_vs_0;
  assign output_31_bits_offset = output_31_bits_offset_0;
  assign output_31_bits_writeIndex = output_31_bits_writeIndex_0;
  assign output_31_bits_dataOffset = output_31_bits_dataOffset_0;
endmodule

