
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module StoreUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [63:0]  maskInput,
  output         maskSelect_valid,
  output [4:0]   maskSelect_bits,
  input          memRequest_ready,
  output         memRequest_valid,
  output [511:0] memRequest_bits_data,
  output [63:0]  memRequest_bits_mask,
  output [5:0]   memRequest_bits_index,
  output [31:0]  memRequest_bits_address,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [1:0]   vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [1:0]   vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [1:0]   vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [1:0]   vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadDataPorts_4_ready,
  output         vrfReadDataPorts_4_valid,
  output [4:0]   vrfReadDataPorts_4_bits_vs,
  output [1:0]   vrfReadDataPorts_4_bits_offset,
  output [2:0]   vrfReadDataPorts_4_bits_instructionIndex,
  input          vrfReadDataPorts_5_ready,
  output         vrfReadDataPorts_5_valid,
  output [4:0]   vrfReadDataPorts_5_bits_vs,
  output [1:0]   vrfReadDataPorts_5_bits_offset,
  output [2:0]   vrfReadDataPorts_5_bits_instructionIndex,
  input          vrfReadDataPorts_6_ready,
  output         vrfReadDataPorts_6_valid,
  output [4:0]   vrfReadDataPorts_6_bits_vs,
  output [1:0]   vrfReadDataPorts_6_bits_offset,
  output [2:0]   vrfReadDataPorts_6_bits_instructionIndex,
  input          vrfReadDataPorts_7_ready,
  output         vrfReadDataPorts_7_valid,
  output [4:0]   vrfReadDataPorts_7_bits_vs,
  output [1:0]   vrfReadDataPorts_7_bits_offset,
  output [2:0]   vrfReadDataPorts_7_bits_instructionIndex,
  input          vrfReadDataPorts_8_ready,
  output         vrfReadDataPorts_8_valid,
  output [4:0]   vrfReadDataPorts_8_bits_vs,
  output [1:0]   vrfReadDataPorts_8_bits_offset,
  output [2:0]   vrfReadDataPorts_8_bits_instructionIndex,
  input          vrfReadDataPorts_9_ready,
  output         vrfReadDataPorts_9_valid,
  output [4:0]   vrfReadDataPorts_9_bits_vs,
  output [1:0]   vrfReadDataPorts_9_bits_offset,
  output [2:0]   vrfReadDataPorts_9_bits_instructionIndex,
  input          vrfReadDataPorts_10_ready,
  output         vrfReadDataPorts_10_valid,
  output [4:0]   vrfReadDataPorts_10_bits_vs,
  output [1:0]   vrfReadDataPorts_10_bits_offset,
  output [2:0]   vrfReadDataPorts_10_bits_instructionIndex,
  input          vrfReadDataPorts_11_ready,
  output         vrfReadDataPorts_11_valid,
  output [4:0]   vrfReadDataPorts_11_bits_vs,
  output [1:0]   vrfReadDataPorts_11_bits_offset,
  output [2:0]   vrfReadDataPorts_11_bits_instructionIndex,
  input          vrfReadDataPorts_12_ready,
  output         vrfReadDataPorts_12_valid,
  output [4:0]   vrfReadDataPorts_12_bits_vs,
  output [1:0]   vrfReadDataPorts_12_bits_offset,
  output [2:0]   vrfReadDataPorts_12_bits_instructionIndex,
  input          vrfReadDataPorts_13_ready,
  output         vrfReadDataPorts_13_valid,
  output [4:0]   vrfReadDataPorts_13_bits_vs,
  output [1:0]   vrfReadDataPorts_13_bits_offset,
  output [2:0]   vrfReadDataPorts_13_bits_instructionIndex,
  input          vrfReadDataPorts_14_ready,
  output         vrfReadDataPorts_14_valid,
  output [4:0]   vrfReadDataPorts_14_bits_vs,
  output [1:0]   vrfReadDataPorts_14_bits_offset,
  output [2:0]   vrfReadDataPorts_14_bits_instructionIndex,
  input          vrfReadDataPorts_15_ready,
  output         vrfReadDataPorts_15_valid,
  output [4:0]   vrfReadDataPorts_15_bits_vs,
  output [1:0]   vrfReadDataPorts_15_bits_offset,
  output [2:0]   vrfReadDataPorts_15_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfReadResults_4_valid,
  input  [31:0]  vrfReadResults_4_bits,
  input          vrfReadResults_5_valid,
  input  [31:0]  vrfReadResults_5_bits,
  input          vrfReadResults_6_valid,
  input  [31:0]  vrfReadResults_6_bits,
  input          vrfReadResults_7_valid,
  input  [31:0]  vrfReadResults_7_bits,
  input          vrfReadResults_8_valid,
  input  [31:0]  vrfReadResults_8_bits,
  input          vrfReadResults_9_valid,
  input  [31:0]  vrfReadResults_9_bits,
  input          vrfReadResults_10_valid,
  input  [31:0]  vrfReadResults_10_bits,
  input          vrfReadResults_11_valid,
  input  [31:0]  vrfReadResults_11_bits,
  input          vrfReadResults_12_valid,
  input  [31:0]  vrfReadResults_12_bits,
  input          vrfReadResults_13_valid,
  input  [31:0]  vrfReadResults_13_bits,
  input          vrfReadResults_14_valid,
  input  [31:0]  vrfReadResults_14_bits,
  input          vrfReadResults_15_valid,
  input  [31:0]  vrfReadResults_15_bits,
  input          storeResponse
);

  wire             _addressQueue_fifo_empty;
  wire             _addressQueue_fifo_full;
  wire             _addressQueue_fifo_error;
  wire             _vrfReadQueueVec_fifo_15_empty;
  wire             _vrfReadQueueVec_fifo_15_full;
  wire             _vrfReadQueueVec_fifo_15_error;
  wire [31:0]      _vrfReadQueueVec_fifo_15_data_out;
  wire             _vrfReadQueueVec_fifo_14_empty;
  wire             _vrfReadQueueVec_fifo_14_full;
  wire             _vrfReadQueueVec_fifo_14_error;
  wire [31:0]      _vrfReadQueueVec_fifo_14_data_out;
  wire             _vrfReadQueueVec_fifo_13_empty;
  wire             _vrfReadQueueVec_fifo_13_full;
  wire             _vrfReadQueueVec_fifo_13_error;
  wire [31:0]      _vrfReadQueueVec_fifo_13_data_out;
  wire             _vrfReadQueueVec_fifo_12_empty;
  wire             _vrfReadQueueVec_fifo_12_full;
  wire             _vrfReadQueueVec_fifo_12_error;
  wire [31:0]      _vrfReadQueueVec_fifo_12_data_out;
  wire             _vrfReadQueueVec_fifo_11_empty;
  wire             _vrfReadQueueVec_fifo_11_full;
  wire             _vrfReadQueueVec_fifo_11_error;
  wire [31:0]      _vrfReadQueueVec_fifo_11_data_out;
  wire             _vrfReadQueueVec_fifo_10_empty;
  wire             _vrfReadQueueVec_fifo_10_full;
  wire             _vrfReadQueueVec_fifo_10_error;
  wire [31:0]      _vrfReadQueueVec_fifo_10_data_out;
  wire             _vrfReadQueueVec_fifo_9_empty;
  wire             _vrfReadQueueVec_fifo_9_full;
  wire             _vrfReadQueueVec_fifo_9_error;
  wire [31:0]      _vrfReadQueueVec_fifo_9_data_out;
  wire             _vrfReadQueueVec_fifo_8_empty;
  wire             _vrfReadQueueVec_fifo_8_full;
  wire             _vrfReadQueueVec_fifo_8_error;
  wire [31:0]      _vrfReadQueueVec_fifo_8_data_out;
  wire             _vrfReadQueueVec_fifo_7_empty;
  wire             _vrfReadQueueVec_fifo_7_full;
  wire             _vrfReadQueueVec_fifo_7_error;
  wire [31:0]      _vrfReadQueueVec_fifo_7_data_out;
  wire             _vrfReadQueueVec_fifo_6_empty;
  wire             _vrfReadQueueVec_fifo_6_full;
  wire             _vrfReadQueueVec_fifo_6_error;
  wire [31:0]      _vrfReadQueueVec_fifo_6_data_out;
  wire             _vrfReadQueueVec_fifo_5_empty;
  wire             _vrfReadQueueVec_fifo_5_full;
  wire             _vrfReadQueueVec_fifo_5_error;
  wire [31:0]      _vrfReadQueueVec_fifo_5_data_out;
  wire             _vrfReadQueueVec_fifo_4_empty;
  wire             _vrfReadQueueVec_fifo_4_full;
  wire             _vrfReadQueueVec_fifo_4_error;
  wire [31:0]      _vrfReadQueueVec_fifo_4_data_out;
  wire             _vrfReadQueueVec_fifo_3_empty;
  wire             _vrfReadQueueVec_fifo_3_full;
  wire             _vrfReadQueueVec_fifo_3_error;
  wire [31:0]      _vrfReadQueueVec_fifo_3_data_out;
  wire             _vrfReadQueueVec_fifo_2_empty;
  wire             _vrfReadQueueVec_fifo_2_full;
  wire             _vrfReadQueueVec_fifo_2_error;
  wire [31:0]      _vrfReadQueueVec_fifo_2_data_out;
  wire             _vrfReadQueueVec_fifo_1_empty;
  wire             _vrfReadQueueVec_fifo_1_full;
  wire             _vrfReadQueueVec_fifo_1_error;
  wire [31:0]      _vrfReadQueueVec_fifo_1_data_out;
  wire             _vrfReadQueueVec_fifo_empty;
  wire             _vrfReadQueueVec_fifo_full;
  wire             _vrfReadQueueVec_fifo_error;
  wire [31:0]      _vrfReadQueueVec_fifo_data_out;
  wire             addressQueue_almostFull;
  wire             addressQueue_almostEmpty;
  wire             vrfReadQueueVec_15_almostFull;
  wire             vrfReadQueueVec_15_almostEmpty;
  wire             vrfReadQueueVec_14_almostFull;
  wire             vrfReadQueueVec_14_almostEmpty;
  wire             vrfReadQueueVec_13_almostFull;
  wire             vrfReadQueueVec_13_almostEmpty;
  wire             vrfReadQueueVec_12_almostFull;
  wire             vrfReadQueueVec_12_almostEmpty;
  wire             vrfReadQueueVec_11_almostFull;
  wire             vrfReadQueueVec_11_almostEmpty;
  wire             vrfReadQueueVec_10_almostFull;
  wire             vrfReadQueueVec_10_almostEmpty;
  wire             vrfReadQueueVec_9_almostFull;
  wire             vrfReadQueueVec_9_almostEmpty;
  wire             vrfReadQueueVec_8_almostFull;
  wire             vrfReadQueueVec_8_almostEmpty;
  wire             vrfReadQueueVec_7_almostFull;
  wire             vrfReadQueueVec_7_almostEmpty;
  wire             vrfReadQueueVec_6_almostFull;
  wire             vrfReadQueueVec_6_almostEmpty;
  wire             vrfReadQueueVec_5_almostFull;
  wire             vrfReadQueueVec_5_almostEmpty;
  wire             vrfReadQueueVec_4_almostFull;
  wire             vrfReadQueueVec_4_almostEmpty;
  wire             vrfReadQueueVec_3_almostFull;
  wire             vrfReadQueueVec_3_almostEmpty;
  wire             vrfReadQueueVec_2_almostFull;
  wire             vrfReadQueueVec_2_almostEmpty;
  wire             vrfReadQueueVec_1_almostFull;
  wire             vrfReadQueueVec_1_almostEmpty;
  wire             vrfReadQueueVec_0_almostFull;
  wire             vrfReadQueueVec_0_almostEmpty;
  wire             memRequest_ready_0 = memRequest_ready;
  wire             vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire             vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire             vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire             vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire             vrfReadDataPorts_4_ready_0 = vrfReadDataPorts_4_ready;
  wire             vrfReadDataPorts_5_ready_0 = vrfReadDataPorts_5_ready;
  wire             vrfReadDataPorts_6_ready_0 = vrfReadDataPorts_6_ready;
  wire             vrfReadDataPorts_7_ready_0 = vrfReadDataPorts_7_ready;
  wire             vrfReadDataPorts_8_ready_0 = vrfReadDataPorts_8_ready;
  wire             vrfReadDataPorts_9_ready_0 = vrfReadDataPorts_9_ready;
  wire             vrfReadDataPorts_10_ready_0 = vrfReadDataPorts_10_ready;
  wire             vrfReadDataPorts_11_ready_0 = vrfReadDataPorts_11_ready;
  wire             vrfReadDataPorts_12_ready_0 = vrfReadDataPorts_12_ready;
  wire             vrfReadDataPorts_13_ready_0 = vrfReadDataPorts_13_ready;
  wire             vrfReadDataPorts_14_ready_0 = vrfReadDataPorts_14_ready;
  wire             vrfReadDataPorts_15_ready_0 = vrfReadDataPorts_15_ready;
  wire             vrfReadQueueVec_0_enq_valid = vrfReadResults_0_valid;
  wire [31:0]      vrfReadQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire             vrfReadQueueVec_1_enq_valid = vrfReadResults_1_valid;
  wire [31:0]      vrfReadQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire             vrfReadQueueVec_2_enq_valid = vrfReadResults_2_valid;
  wire [31:0]      vrfReadQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire             vrfReadQueueVec_3_enq_valid = vrfReadResults_3_valid;
  wire [31:0]      vrfReadQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire             vrfReadQueueVec_4_enq_valid = vrfReadResults_4_valid;
  wire [31:0]      vrfReadQueueVec_4_enq_bits = vrfReadResults_4_bits;
  wire             vrfReadQueueVec_5_enq_valid = vrfReadResults_5_valid;
  wire [31:0]      vrfReadQueueVec_5_enq_bits = vrfReadResults_5_bits;
  wire             vrfReadQueueVec_6_enq_valid = vrfReadResults_6_valid;
  wire [31:0]      vrfReadQueueVec_6_enq_bits = vrfReadResults_6_bits;
  wire             vrfReadQueueVec_7_enq_valid = vrfReadResults_7_valid;
  wire [31:0]      vrfReadQueueVec_7_enq_bits = vrfReadResults_7_bits;
  wire             vrfReadQueueVec_8_enq_valid = vrfReadResults_8_valid;
  wire [31:0]      vrfReadQueueVec_8_enq_bits = vrfReadResults_8_bits;
  wire             vrfReadQueueVec_9_enq_valid = vrfReadResults_9_valid;
  wire [31:0]      vrfReadQueueVec_9_enq_bits = vrfReadResults_9_bits;
  wire             vrfReadQueueVec_10_enq_valid = vrfReadResults_10_valid;
  wire [31:0]      vrfReadQueueVec_10_enq_bits = vrfReadResults_10_bits;
  wire             vrfReadQueueVec_11_enq_valid = vrfReadResults_11_valid;
  wire [31:0]      vrfReadQueueVec_11_enq_bits = vrfReadResults_11_bits;
  wire             vrfReadQueueVec_12_enq_valid = vrfReadResults_12_valid;
  wire [31:0]      vrfReadQueueVec_12_enq_bits = vrfReadResults_12_bits;
  wire             vrfReadQueueVec_13_enq_valid = vrfReadResults_13_valid;
  wire [31:0]      vrfReadQueueVec_13_enq_bits = vrfReadResults_13_bits;
  wire             vrfReadQueueVec_14_enq_valid = vrfReadResults_14_valid;
  wire [31:0]      vrfReadQueueVec_14_enq_bits = vrfReadResults_14_bits;
  wire             vrfReadQueueVec_15_enq_valid = vrfReadResults_15_valid;
  wire [31:0]      vrfReadQueueVec_15_enq_bits = vrfReadResults_15_bits;
  wire             addressQueue_deq_ready = storeResponse;
  wire [1:0]       accessStateCheck_lo_lo_lo = 2'h0;
  wire [1:0]       accessStateCheck_lo_lo_hi = 2'h0;
  wire [1:0]       accessStateCheck_lo_hi_lo = 2'h0;
  wire [1:0]       accessStateCheck_lo_hi_hi = 2'h0;
  wire [1:0]       accessStateCheck_hi_lo_lo = 2'h0;
  wire [1:0]       accessStateCheck_hi_lo_hi = 2'h0;
  wire [1:0]       accessStateCheck_hi_hi_lo = 2'h0;
  wire [1:0]       accessStateCheck_hi_hi_hi = 2'h0;
  wire [3:0]       accessStateCheck_lo_lo = 4'h0;
  wire [3:0]       accessStateCheck_lo_hi = 4'h0;
  wire [3:0]       accessStateCheck_hi_lo = 4'h0;
  wire [3:0]       accessStateCheck_hi_hi = 4'h0;
  wire [7:0]       accessStateCheck_lo = 8'h0;
  wire [7:0]       accessStateCheck_hi = 8'h0;
  wire             accessStateCheck = 1'h1;
  wire             accessStateUpdate_0 = 1'h0;
  wire             accessStateUpdate_1 = 1'h0;
  wire             accessStateUpdate_2 = 1'h0;
  wire             accessStateUpdate_3 = 1'h0;
  wire             accessStateUpdate_4 = 1'h0;
  wire             accessStateUpdate_5 = 1'h0;
  wire             accessStateUpdate_6 = 1'h0;
  wire             accessStateUpdate_7 = 1'h0;
  wire             accessStateUpdate_8 = 1'h0;
  wire             accessStateUpdate_9 = 1'h0;
  wire             accessStateUpdate_10 = 1'h0;
  wire             accessStateUpdate_11 = 1'h0;
  wire             accessStateUpdate_12 = 1'h0;
  wire             accessStateUpdate_13 = 1'h0;
  wire             accessStateUpdate_14 = 1'h0;
  wire             accessStateUpdate_15 = 1'h0;
  wire [2047:0]    hi = 2048'h0;
  wire [2047:0]    hi_1 = 2048'h0;
  wire [2047:0]    hi_2 = 2048'h0;
  wire [2047:0]    hi_3 = 2048'h0;
  wire [2047:0]    hi_8 = 2048'h0;
  wire [2047:0]    hi_9 = 2048'h0;
  wire [2047:0]    hi_10 = 2048'h0;
  wire [2047:0]    hi_11 = 2048'h0;
  wire [2047:0]    hi_16 = 2048'h0;
  wire [2047:0]    hi_17 = 2048'h0;
  wire [2047:0]    hi_18 = 2048'h0;
  wire [2047:0]    hi_19 = 2048'h0;
  wire [1023:0]    lo_hi = 1024'h0;
  wire [1023:0]    hi_lo = 1024'h0;
  wire [1023:0]    hi_hi = 1024'h0;
  wire [1023:0]    lo_hi_1 = 1024'h0;
  wire [1023:0]    hi_lo_1 = 1024'h0;
  wire [1023:0]    hi_hi_1 = 1024'h0;
  wire [1023:0]    hi_lo_2 = 1024'h0;
  wire [1023:0]    hi_hi_2 = 1024'h0;
  wire [1023:0]    hi_lo_3 = 1024'h0;
  wire [1023:0]    hi_hi_3 = 1024'h0;
  wire [1023:0]    hi_hi_4 = 1024'h0;
  wire [1023:0]    hi_hi_5 = 1024'h0;
  wire [1023:0]    lo_hi_8 = 1024'h0;
  wire [1023:0]    hi_lo_8 = 1024'h0;
  wire [1023:0]    hi_hi_8 = 1024'h0;
  wire [1023:0]    lo_hi_9 = 1024'h0;
  wire [1023:0]    hi_lo_9 = 1024'h0;
  wire [1023:0]    hi_hi_9 = 1024'h0;
  wire [1023:0]    hi_lo_10 = 1024'h0;
  wire [1023:0]    hi_hi_10 = 1024'h0;
  wire [1023:0]    hi_lo_11 = 1024'h0;
  wire [1023:0]    hi_hi_11 = 1024'h0;
  wire [1023:0]    hi_hi_12 = 1024'h0;
  wire [1023:0]    hi_hi_13 = 1024'h0;
  wire [1023:0]    lo_hi_16 = 1024'h0;
  wire [1023:0]    hi_lo_16 = 1024'h0;
  wire [1023:0]    hi_hi_16 = 1024'h0;
  wire [1023:0]    lo_hi_17 = 1024'h0;
  wire [1023:0]    hi_lo_17 = 1024'h0;
  wire [1023:0]    hi_hi_17 = 1024'h0;
  wire [1023:0]    hi_lo_18 = 1024'h0;
  wire [1023:0]    hi_hi_18 = 1024'h0;
  wire [1023:0]    hi_lo_19 = 1024'h0;
  wire [1023:0]    hi_hi_19 = 1024'h0;
  wire [1023:0]    hi_hi_20 = 1024'h0;
  wire [1023:0]    hi_hi_21 = 1024'h0;
  wire [511:0]     res_1 = 512'h0;
  wire [511:0]     res_2 = 512'h0;
  wire [511:0]     res_3 = 512'h0;
  wire [511:0]     res_4 = 512'h0;
  wire [511:0]     res_5 = 512'h0;
  wire [511:0]     res_6 = 512'h0;
  wire [511:0]     res_7 = 512'h0;
  wire [511:0]     res_10 = 512'h0;
  wire [511:0]     res_11 = 512'h0;
  wire [511:0]     res_12 = 512'h0;
  wire [511:0]     res_13 = 512'h0;
  wire [511:0]     res_14 = 512'h0;
  wire [511:0]     res_15 = 512'h0;
  wire [511:0]     res_19 = 512'h0;
  wire [511:0]     res_20 = 512'h0;
  wire [511:0]     res_21 = 512'h0;
  wire [511:0]     res_22 = 512'h0;
  wire [511:0]     res_23 = 512'h0;
  wire [511:0]     res_28 = 512'h0;
  wire [511:0]     res_29 = 512'h0;
  wire [511:0]     res_30 = 512'h0;
  wire [511:0]     res_31 = 512'h0;
  wire [511:0]     res_37 = 512'h0;
  wire [511:0]     res_38 = 512'h0;
  wire [511:0]     res_39 = 512'h0;
  wire [511:0]     res_46 = 512'h0;
  wire [511:0]     res_47 = 512'h0;
  wire [511:0]     res_55 = 512'h0;
  wire [511:0]     res_65 = 512'h0;
  wire [511:0]     res_66 = 512'h0;
  wire [511:0]     res_67 = 512'h0;
  wire [511:0]     res_68 = 512'h0;
  wire [511:0]     res_69 = 512'h0;
  wire [511:0]     res_70 = 512'h0;
  wire [511:0]     res_71 = 512'h0;
  wire [511:0]     res_74 = 512'h0;
  wire [511:0]     res_75 = 512'h0;
  wire [511:0]     res_76 = 512'h0;
  wire [511:0]     res_77 = 512'h0;
  wire [511:0]     res_78 = 512'h0;
  wire [511:0]     res_79 = 512'h0;
  wire [511:0]     res_83 = 512'h0;
  wire [511:0]     res_84 = 512'h0;
  wire [511:0]     res_85 = 512'h0;
  wire [511:0]     res_86 = 512'h0;
  wire [511:0]     res_87 = 512'h0;
  wire [511:0]     res_92 = 512'h0;
  wire [511:0]     res_93 = 512'h0;
  wire [511:0]     res_94 = 512'h0;
  wire [511:0]     res_95 = 512'h0;
  wire [511:0]     res_101 = 512'h0;
  wire [511:0]     res_102 = 512'h0;
  wire [511:0]     res_103 = 512'h0;
  wire [511:0]     res_110 = 512'h0;
  wire [511:0]     res_111 = 512'h0;
  wire [511:0]     res_119 = 512'h0;
  wire [511:0]     res_129 = 512'h0;
  wire [511:0]     res_130 = 512'h0;
  wire [511:0]     res_131 = 512'h0;
  wire [511:0]     res_132 = 512'h0;
  wire [511:0]     res_133 = 512'h0;
  wire [511:0]     res_134 = 512'h0;
  wire [511:0]     res_135 = 512'h0;
  wire [511:0]     res_138 = 512'h0;
  wire [511:0]     res_139 = 512'h0;
  wire [511:0]     res_140 = 512'h0;
  wire [511:0]     res_141 = 512'h0;
  wire [511:0]     res_142 = 512'h0;
  wire [511:0]     res_143 = 512'h0;
  wire [511:0]     res_147 = 512'h0;
  wire [511:0]     res_148 = 512'h0;
  wire [511:0]     res_149 = 512'h0;
  wire [511:0]     res_150 = 512'h0;
  wire [511:0]     res_151 = 512'h0;
  wire [511:0]     res_156 = 512'h0;
  wire [511:0]     res_157 = 512'h0;
  wire [511:0]     res_158 = 512'h0;
  wire [511:0]     res_159 = 512'h0;
  wire [511:0]     res_165 = 512'h0;
  wire [511:0]     res_166 = 512'h0;
  wire [511:0]     res_167 = 512'h0;
  wire [511:0]     res_174 = 512'h0;
  wire [511:0]     res_175 = 512'h0;
  wire [511:0]     res_183 = 512'h0;
  wire [1:0]       vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_4_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_5_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_6_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_7_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_8_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_9_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_10_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_11_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_12_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_13_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_14_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_15_bits_readSource = 2'h2;
  wire [31:0]      alignedDequeueAddress;
  reg  [2:0]       lsuRequestReg_instructionInformation_nf;
  reg              lsuRequestReg_instructionInformation_mew;
  reg  [1:0]       lsuRequestReg_instructionInformation_mop;
  reg  [4:0]       lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]       lsuRequestReg_instructionInformation_eew;
  reg  [4:0]       lsuRequestReg_instructionInformation_vs3;
  reg              lsuRequestReg_instructionInformation_isStore;
  reg              lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]      lsuRequestReg_rs1Data;
  reg  [31:0]      lsuRequestReg_rs2Data;
  reg  [2:0]       lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_4_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_5_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_6_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_7_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_8_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_9_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_10_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_11_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_12_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_13_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_14_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_15_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [11:0]      csrInterfaceReg_vl;
  reg  [11:0]      csrInterfaceReg_vStart;
  reg  [2:0]       csrInterfaceReg_vlmul;
  reg  [1:0]       csrInterfaceReg_vSew;
  reg  [1:0]       csrInterfaceReg_vxrm;
  reg              csrInterfaceReg_vta;
  reg              csrInterfaceReg_vma;
  reg              requestFireNext;
  reg  [1:0]       dataEEW;
  wire [3:0]       _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]       dataEEWOH = _dataEEWOH_T[2:0];
  wire             isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [63:0]      maskAmend = isMaskType ? maskInput : 64'hFFFFFFFFFFFFFFFF;
  reg  [63:0]      maskReg;
  wire [63:0]      _lastMaskAmend_T_1 = 64'h1 << csrInterface_vl[5:0];
  wire [61:0]      _GEN = _lastMaskAmend_T_1[62:1] | _lastMaskAmend_T_1[63:2];
  wire [60:0]      _GEN_0 = _GEN[60:0] | {_lastMaskAmend_T_1[63], _GEN[61:2]};
  wire [58:0]      _GEN_1 = _GEN_0[58:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:4]};
  wire [54:0]      _GEN_2 = _GEN_1[54:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:8]};
  wire [46:0]      _GEN_3 = _GEN_2[46:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:16]};
  wire [62:0]      lastMaskAmend =
    {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:47], _GEN_3[46:31], _GEN_3[30:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:47], _GEN_3[46:32]}};
  reg              needAmend;
  reg  [62:0]      lastMaskAmendReg;
  wire [1:0]       countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [4:0]       maskGroupCounter;
  wire [4:0]       nextMaskGroup = maskGroupCounter + 5'h1;
  reg  [1:0]       maskCounterInGroup;
  wire [1:0]       nextMaskCount = maskCounterInGroup + 2'h1;
  wire             isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [4:0]       _maskSelect_bits_output = lsuRequest_valid ? 5'h0 : nextMaskGroup;
  reg              isLastMaskGroup;
  wire [63:0]      maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 64'hFFFFFFFFFFFFFFFF);
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo = {maskForGroupWire_lo_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi = {maskForGroupWire_lo_lo_lo_hi_hi, maskForGroupWire_lo_lo_lo_hi_lo};
  wire [15:0]      maskForGroupWire_lo_lo_lo = {maskForGroupWire_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo = {maskForGroupWire_lo_lo_hi_lo_hi, maskForGroupWire_lo_lo_hi_lo_lo};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi = {maskForGroupWire_lo_lo_hi_hi_hi, maskForGroupWire_lo_lo_hi_hi_lo};
  wire [15:0]      maskForGroupWire_lo_lo_hi = {maskForGroupWire_lo_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo};
  wire [31:0]      maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo_lo = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo_hi = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo = {maskForGroupWire_lo_hi_lo_lo_hi, maskForGroupWire_lo_hi_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi_lo = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi_hi = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi = {maskForGroupWire_lo_hi_lo_hi_hi, maskForGroupWire_lo_hi_lo_hi_lo};
  wire [15:0]      maskForGroupWire_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo_lo = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo_hi = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo = {maskForGroupWire_lo_hi_hi_lo_hi, maskForGroupWire_lo_hi_hi_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi_lo = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi_hi = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi = {maskForGroupWire_lo_hi_hi_hi_hi, maskForGroupWire_lo_hi_hi_hi_lo};
  wire [15:0]      maskForGroupWire_lo_hi_hi = {maskForGroupWire_lo_hi_hi_hi, maskForGroupWire_lo_hi_hi_lo};
  wire [31:0]      maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [63:0]      maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo_lo = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo_hi = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo = {maskForGroupWire_hi_lo_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi_lo = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi_hi = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi = {maskForGroupWire_hi_lo_lo_hi_hi, maskForGroupWire_hi_lo_lo_hi_lo};
  wire [15:0]      maskForGroupWire_hi_lo_lo = {maskForGroupWire_hi_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo_lo = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo_hi = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo = {maskForGroupWire_hi_lo_hi_lo_hi, maskForGroupWire_hi_lo_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi_lo = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi_hi = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi = {maskForGroupWire_hi_lo_hi_hi_hi, maskForGroupWire_hi_lo_hi_hi_lo};
  wire [15:0]      maskForGroupWire_hi_lo_hi = {maskForGroupWire_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo};
  wire [31:0]      maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo_lo = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo_hi = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo = {maskForGroupWire_hi_hi_lo_lo_hi, maskForGroupWire_hi_hi_lo_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi_lo = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi_hi = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi = {maskForGroupWire_hi_hi_lo_hi_hi, maskForGroupWire_hi_hi_lo_hi_lo};
  wire [15:0]      maskForGroupWire_hi_hi_lo = {maskForGroupWire_hi_hi_lo_hi, maskForGroupWire_hi_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo_lo = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo_hi = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo = {maskForGroupWire_hi_hi_hi_lo_hi, maskForGroupWire_hi_hi_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi_lo = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi_hi = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_hi_lo};
  wire [15:0]      maskForGroupWire_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_lo};
  wire [31:0]      maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [63:0]      maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_1 = {maskForGroupWire_lo_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_1 = {maskForGroupWire_lo_lo_hi_lo_hi_1, maskForGroupWire_lo_lo_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_1 = {maskForGroupWire_lo_lo_hi_hi_hi_1, maskForGroupWire_lo_lo_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_lo_hi_1 = {maskForGroupWire_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_1};
  wire [31:0]      maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo_lo_1 = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo_hi_1 = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_1 = {maskForGroupWire_lo_hi_lo_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi_lo_1 = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi_hi_1 = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_1 = {maskForGroupWire_lo_hi_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo_lo_1 = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo_hi_1 = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_1 = {maskForGroupWire_lo_hi_hi_lo_hi_1, maskForGroupWire_lo_hi_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi_lo_1 = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi_hi_1 = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_1};
  wire [31:0]      maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [63:0]      maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo_lo_1 = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo_hi_1 = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_1 = {maskForGroupWire_hi_lo_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi_lo_1 = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi_hi_1 = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_1 = {maskForGroupWire_hi_lo_lo_hi_hi_1, maskForGroupWire_hi_lo_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_lo_lo_1 = {maskForGroupWire_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo_lo_1 = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo_hi_1 = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_1 = {maskForGroupWire_hi_lo_hi_lo_hi_1, maskForGroupWire_hi_lo_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi_lo_1 = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi_hi_1 = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_1 = {maskForGroupWire_hi_lo_hi_hi_hi_1, maskForGroupWire_hi_lo_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_1};
  wire [31:0]      maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo_lo_1 = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo_hi_1 = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_1 = {maskForGroupWire_hi_hi_lo_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi_lo_1 = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi_hi_1 = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_1 = {maskForGroupWire_hi_hi_lo_hi_hi_1, maskForGroupWire_hi_hi_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo_lo_1 = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo_hi_1 = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_1 = {maskForGroupWire_hi_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi_lo_1 = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi_hi_1 = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_1};
  wire [31:0]      maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [63:0]      maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]       _maskForGroupWire_T_261 = 4'h1 << maskCounterInGroup;
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_hi_2 = {maskForGroupWire_lo_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_lo_2 = {maskForGroupWire_lo_lo_hi_lo_hi_2, maskForGroupWire_lo_lo_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_hi_2 = {maskForGroupWire_lo_lo_hi_hi_hi_2, maskForGroupWire_lo_lo_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_lo_hi_2 = {maskForGroupWire_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_2};
  wire [63:0]      maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_lo_2 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_hi_2 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_lo_2 = {maskForGroupWire_lo_hi_lo_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_lo_2 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_hi_2 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_hi_2 = {maskForGroupWire_lo_hi_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_lo_2 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_hi_2 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_lo_2 = {maskForGroupWire_lo_hi_hi_lo_hi_2, maskForGroupWire_lo_hi_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_lo_2 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_hi_2 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_2};
  wire [63:0]      maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [127:0]     maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_lo_2 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_hi_2 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_lo_2 = {maskForGroupWire_hi_lo_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_lo_2 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_hi_2 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_hi_2 = {maskForGroupWire_hi_lo_lo_hi_hi_2, maskForGroupWire_hi_lo_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_lo_lo_2 = {maskForGroupWire_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_lo_2 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_hi_2 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_lo_2 = {maskForGroupWire_hi_lo_hi_lo_hi_2, maskForGroupWire_hi_lo_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_lo_2 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_hi_2 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_hi_2 = {maskForGroupWire_hi_lo_hi_hi_hi_2, maskForGroupWire_hi_lo_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_2};
  wire [63:0]      maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_lo_2 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_hi_2 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_lo_2 = {maskForGroupWire_hi_hi_lo_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_lo_2 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_hi_2 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_hi_2 = {maskForGroupWire_hi_hi_lo_hi_hi_2, maskForGroupWire_hi_hi_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_lo_2 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_hi_2 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_lo_2 = {maskForGroupWire_hi_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_lo_2 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_hi_2 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_2};
  wire [63:0]      maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [127:0]     maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_hi_3 = {maskForGroupWire_lo_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_lo_3 = {maskForGroupWire_lo_lo_hi_lo_hi_3, maskForGroupWire_lo_lo_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_hi_3 = {maskForGroupWire_lo_lo_hi_hi_hi_3, maskForGroupWire_lo_lo_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_lo_hi_3 = {maskForGroupWire_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_3};
  wire [63:0]      maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_lo_3 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_hi_3 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_lo_3 = {maskForGroupWire_lo_hi_lo_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_lo_3 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_hi_3 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_hi_3 = {maskForGroupWire_lo_hi_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_lo_3 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_hi_3 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_lo_3 = {maskForGroupWire_lo_hi_hi_lo_hi_3, maskForGroupWire_lo_hi_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_lo_3 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_hi_3 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_3};
  wire [63:0]      maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [127:0]     maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_lo_3 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_hi_3 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_lo_3 = {maskForGroupWire_hi_lo_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_lo_3 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_hi_3 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_hi_3 = {maskForGroupWire_hi_lo_lo_hi_hi_3, maskForGroupWire_hi_lo_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_lo_lo_3 = {maskForGroupWire_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_lo_3 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_hi_3 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_lo_3 = {maskForGroupWire_hi_lo_hi_lo_hi_3, maskForGroupWire_hi_lo_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_lo_3 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_hi_3 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_hi_3 = {maskForGroupWire_hi_lo_hi_hi_hi_3, maskForGroupWire_hi_lo_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_3};
  wire [63:0]      maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_lo_3 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_hi_3 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_lo_3 = {maskForGroupWire_hi_hi_lo_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_lo_3 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_hi_3 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_hi_3 = {maskForGroupWire_hi_hi_lo_hi_hi_3, maskForGroupWire_hi_hi_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_lo_3 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_hi_3 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_lo_3 = {maskForGroupWire_hi_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_lo_3 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_hi_3 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_3};
  wire [63:0]      maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [127:0]     maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_hi_4 = {maskForGroupWire_lo_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_lo_4 = {maskForGroupWire_lo_lo_hi_lo_hi_4, maskForGroupWire_lo_lo_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_hi_4 = {maskForGroupWire_lo_lo_hi_hi_hi_4, maskForGroupWire_lo_lo_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_lo_hi_4 = {maskForGroupWire_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_4};
  wire [63:0]      maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_lo_4 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_hi_4 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_lo_4 = {maskForGroupWire_lo_hi_lo_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_lo_4 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_hi_4 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_hi_4 = {maskForGroupWire_lo_hi_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_lo_4 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_hi_4 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_lo_4 = {maskForGroupWire_lo_hi_hi_lo_hi_4, maskForGroupWire_lo_hi_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_lo_4 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_hi_4 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_4};
  wire [63:0]      maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [127:0]     maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_lo_4 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_hi_4 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_lo_4 = {maskForGroupWire_hi_lo_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_lo_4 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_hi_4 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_hi_4 = {maskForGroupWire_hi_lo_lo_hi_hi_4, maskForGroupWire_hi_lo_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_lo_lo_4 = {maskForGroupWire_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_lo_4 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_hi_4 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_lo_4 = {maskForGroupWire_hi_lo_hi_lo_hi_4, maskForGroupWire_hi_lo_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_lo_4 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_hi_4 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_hi_4 = {maskForGroupWire_hi_lo_hi_hi_hi_4, maskForGroupWire_hi_lo_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_4};
  wire [63:0]      maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_lo_4 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_hi_4 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_lo_4 = {maskForGroupWire_hi_hi_lo_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_lo_4 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_hi_4 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_hi_4 = {maskForGroupWire_hi_hi_lo_hi_hi_4, maskForGroupWire_hi_hi_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_lo_4 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_hi_4 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_lo_4 = {maskForGroupWire_hi_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_lo_4 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_hi_4 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_4};
  wire [63:0]      maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [127:0]     maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_hi_5 = {maskForGroupWire_lo_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_lo_5 = {maskForGroupWire_lo_lo_hi_lo_hi_5, maskForGroupWire_lo_lo_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_hi_5 = {maskForGroupWire_lo_lo_hi_hi_hi_5, maskForGroupWire_lo_lo_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_lo_hi_5 = {maskForGroupWire_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_5};
  wire [63:0]      maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_lo_5 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_hi_5 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_lo_5 = {maskForGroupWire_lo_hi_lo_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_lo_5 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_hi_5 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_hi_5 = {maskForGroupWire_lo_hi_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_lo_5 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_hi_5 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_lo_5 = {maskForGroupWire_lo_hi_hi_lo_hi_5, maskForGroupWire_lo_hi_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_lo_5 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_hi_5 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_5};
  wire [63:0]      maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [127:0]     maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_lo_5 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_hi_5 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_lo_5 = {maskForGroupWire_hi_lo_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_lo_5 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_hi_5 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_hi_5 = {maskForGroupWire_hi_lo_lo_hi_hi_5, maskForGroupWire_hi_lo_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_lo_lo_5 = {maskForGroupWire_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_lo_5 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_hi_5 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_lo_5 = {maskForGroupWire_hi_lo_hi_lo_hi_5, maskForGroupWire_hi_lo_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_lo_5 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_hi_5 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_hi_5 = {maskForGroupWire_hi_lo_hi_hi_hi_5, maskForGroupWire_hi_lo_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_5};
  wire [63:0]      maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_lo_5 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_hi_5 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_lo_5 = {maskForGroupWire_hi_hi_lo_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_lo_5 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_hi_5 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_hi_5 = {maskForGroupWire_hi_hi_lo_hi_hi_5, maskForGroupWire_hi_hi_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_lo_5 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_hi_5 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_lo_5 = {maskForGroupWire_hi_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_lo_5 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_hi_5 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_5};
  wire [63:0]      maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [127:0]     maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [63:0]      maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 64'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 64'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_261[0] ? maskForGroupWire_lo_2[63:0] : 64'h0) | (_maskForGroupWire_T_261[1] ? maskForGroupWire_lo_3[127:64] : 64'h0) | (_maskForGroupWire_T_261[2] ? maskForGroupWire_hi_4[63:0] : 64'h0)
           | (_maskForGroupWire_T_261[3] ? maskForGroupWire_hi_5[127:64] : 64'h0)
         : 64'h0);
  wire [1:0]       initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]       fillBySeg_lo_lo_lo_lo_lo = maskForGroupWire[1:0];
  wire [1:0]       initSendState_hi = maskForGroupWire[3:2];
  wire [1:0]       fillBySeg_lo_lo_lo_lo_hi = maskForGroupWire[3:2];
  wire             initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]       initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]       fillBySeg_lo_lo_lo_hi_lo = maskForGroupWire[5:4];
  wire [1:0]       initSendState_hi_1 = maskForGroupWire[7:6];
  wire [1:0]       fillBySeg_lo_lo_lo_hi_hi = maskForGroupWire[7:6];
  wire             initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]       initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]       fillBySeg_lo_lo_hi_lo_lo = maskForGroupWire[9:8];
  wire [1:0]       initSendState_hi_2 = maskForGroupWire[11:10];
  wire [1:0]       fillBySeg_lo_lo_hi_lo_hi = maskForGroupWire[11:10];
  wire             initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]       initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]       fillBySeg_lo_lo_hi_hi_lo = maskForGroupWire[13:12];
  wire [1:0]       initSendState_hi_3 = maskForGroupWire[15:14];
  wire [1:0]       fillBySeg_lo_lo_hi_hi_hi = maskForGroupWire[15:14];
  wire             initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  wire [1:0]       initSendState_lo_4 = maskForGroupWire[17:16];
  wire [1:0]       fillBySeg_lo_hi_lo_lo_lo = maskForGroupWire[17:16];
  wire [1:0]       initSendState_hi_4 = maskForGroupWire[19:18];
  wire [1:0]       fillBySeg_lo_hi_lo_lo_hi = maskForGroupWire[19:18];
  wire             initSendState_4 = |{initSendState_hi_4, initSendState_lo_4};
  wire [1:0]       initSendState_lo_5 = maskForGroupWire[21:20];
  wire [1:0]       fillBySeg_lo_hi_lo_hi_lo = maskForGroupWire[21:20];
  wire [1:0]       initSendState_hi_5 = maskForGroupWire[23:22];
  wire [1:0]       fillBySeg_lo_hi_lo_hi_hi = maskForGroupWire[23:22];
  wire             initSendState_5 = |{initSendState_hi_5, initSendState_lo_5};
  wire [1:0]       initSendState_lo_6 = maskForGroupWire[25:24];
  wire [1:0]       fillBySeg_lo_hi_hi_lo_lo = maskForGroupWire[25:24];
  wire [1:0]       initSendState_hi_6 = maskForGroupWire[27:26];
  wire [1:0]       fillBySeg_lo_hi_hi_lo_hi = maskForGroupWire[27:26];
  wire             initSendState_6 = |{initSendState_hi_6, initSendState_lo_6};
  wire [1:0]       initSendState_lo_7 = maskForGroupWire[29:28];
  wire [1:0]       fillBySeg_lo_hi_hi_hi_lo = maskForGroupWire[29:28];
  wire [1:0]       initSendState_hi_7 = maskForGroupWire[31:30];
  wire [1:0]       fillBySeg_lo_hi_hi_hi_hi = maskForGroupWire[31:30];
  wire             initSendState_7 = |{initSendState_hi_7, initSendState_lo_7};
  wire [1:0]       initSendState_lo_8 = maskForGroupWire[33:32];
  wire [1:0]       fillBySeg_hi_lo_lo_lo_lo = maskForGroupWire[33:32];
  wire [1:0]       initSendState_hi_8 = maskForGroupWire[35:34];
  wire [1:0]       fillBySeg_hi_lo_lo_lo_hi = maskForGroupWire[35:34];
  wire             initSendState_8 = |{initSendState_hi_8, initSendState_lo_8};
  wire [1:0]       initSendState_lo_9 = maskForGroupWire[37:36];
  wire [1:0]       fillBySeg_hi_lo_lo_hi_lo = maskForGroupWire[37:36];
  wire [1:0]       initSendState_hi_9 = maskForGroupWire[39:38];
  wire [1:0]       fillBySeg_hi_lo_lo_hi_hi = maskForGroupWire[39:38];
  wire             initSendState_9 = |{initSendState_hi_9, initSendState_lo_9};
  wire [1:0]       initSendState_lo_10 = maskForGroupWire[41:40];
  wire [1:0]       fillBySeg_hi_lo_hi_lo_lo = maskForGroupWire[41:40];
  wire [1:0]       initSendState_hi_10 = maskForGroupWire[43:42];
  wire [1:0]       fillBySeg_hi_lo_hi_lo_hi = maskForGroupWire[43:42];
  wire             initSendState_10 = |{initSendState_hi_10, initSendState_lo_10};
  wire [1:0]       initSendState_lo_11 = maskForGroupWire[45:44];
  wire [1:0]       fillBySeg_hi_lo_hi_hi_lo = maskForGroupWire[45:44];
  wire [1:0]       initSendState_hi_11 = maskForGroupWire[47:46];
  wire [1:0]       fillBySeg_hi_lo_hi_hi_hi = maskForGroupWire[47:46];
  wire             initSendState_11 = |{initSendState_hi_11, initSendState_lo_11};
  wire [1:0]       initSendState_lo_12 = maskForGroupWire[49:48];
  wire [1:0]       fillBySeg_hi_hi_lo_lo_lo = maskForGroupWire[49:48];
  wire [1:0]       initSendState_hi_12 = maskForGroupWire[51:50];
  wire [1:0]       fillBySeg_hi_hi_lo_lo_hi = maskForGroupWire[51:50];
  wire             initSendState_12 = |{initSendState_hi_12, initSendState_lo_12};
  wire [1:0]       initSendState_lo_13 = maskForGroupWire[53:52];
  wire [1:0]       fillBySeg_hi_hi_lo_hi_lo = maskForGroupWire[53:52];
  wire [1:0]       initSendState_hi_13 = maskForGroupWire[55:54];
  wire [1:0]       fillBySeg_hi_hi_lo_hi_hi = maskForGroupWire[55:54];
  wire             initSendState_13 = |{initSendState_hi_13, initSendState_lo_13};
  wire [1:0]       initSendState_lo_14 = maskForGroupWire[57:56];
  wire [1:0]       fillBySeg_hi_hi_hi_lo_lo = maskForGroupWire[57:56];
  wire [1:0]       initSendState_hi_14 = maskForGroupWire[59:58];
  wire [1:0]       fillBySeg_hi_hi_hi_lo_hi = maskForGroupWire[59:58];
  wire             initSendState_14 = |{initSendState_hi_14, initSendState_lo_14};
  wire [1:0]       initSendState_lo_15 = maskForGroupWire[61:60];
  wire [1:0]       fillBySeg_hi_hi_hi_hi_lo = maskForGroupWire[61:60];
  wire [1:0]       initSendState_hi_15 = maskForGroupWire[63:62];
  wire [1:0]       fillBySeg_hi_hi_hi_hi_hi = maskForGroupWire[63:62];
  wire             initSendState_15 = |{initSendState_hi_15, initSendState_lo_15};
  reg  [511:0]     accessData_0;
  wire [511:0]     accessDataUpdate_1 = accessData_0;
  reg  [511:0]     accessData_1;
  wire [511:0]     accessDataUpdate_2 = accessData_1;
  reg  [511:0]     accessData_2;
  wire [511:0]     accessDataUpdate_3 = accessData_2;
  reg  [511:0]     accessData_3;
  wire [511:0]     accessDataUpdate_4 = accessData_3;
  reg  [511:0]     accessData_4;
  wire [511:0]     accessDataUpdate_5 = accessData_4;
  reg  [511:0]     accessData_5;
  wire [511:0]     accessDataUpdate_6 = accessData_5;
  reg  [511:0]     accessData_6;
  wire [511:0]     accessDataUpdate_7 = accessData_6;
  reg  [511:0]     accessData_7;
  reg  [2:0]       accessPtr;
  reg  [4:0]       dataGroup;
  reg  [511:0]     dataBuffer_0;
  reg  [511:0]     dataBuffer_1;
  reg  [511:0]     dataBuffer_2;
  reg  [511:0]     dataBuffer_3;
  reg  [511:0]     dataBuffer_4;
  reg  [511:0]     dataBuffer_5;
  reg  [511:0]     dataBuffer_6;
  reg  [511:0]     dataBuffer_7;
  reg  [5:0]       bufferBaseCacheLineIndex;
  wire [5:0]       memRequest_bits_index_0 = bufferBaseCacheLineIndex;
  reg  [2:0]       cacheLineIndexInBuffer;
  wire [5:0]       initOffset = lsuRequestReg_rs1Data[5:0];
  wire             invalidInstruction = csrInterface_vl == 12'h0;
  reg              invalidInstructionNext;
  wire             wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]       nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]       segmentInstructionIndexInterval;
  wire [18:0]      bytePerInstruction = {3'h0, {12'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [18:0]      accessMemSize = bytePerInstruction + {13'h0, lsuRequest_bits_rs1Data[5:0]};
  wire [12:0]      lastCacheLineIndex = accessMemSize[18:6] - {12'h0, accessMemSize[5:0] == 6'h0};
  wire [12:0]      lastWriteVrfIndex = bytePerInstruction[18:6] - {12'h0, bytePerInstruction[5:0] == 6'h0};
  reg  [12:0]      lastWriteVrfIndexReg;
  reg              lastCacheNeedPush;
  reg  [12:0]      cacheLineNumberReg;
  wire [14:0]      dataByteSize = {3'h0, csrInterface_vl} << lsuRequest_bits_instructionInformation_eew;
  wire [8:0]       lastDataGroupForInstruction = dataByteSize[14:6] - {8'h0, dataByteSize[5:0] == 6'h0};
  reg  [8:0]       lastDataGroupReg;
  wire [4:0]       nextDataGroup = lsuRequest_valid ? 5'h0 : dataGroup + 5'h1;
  wire             isLastRead = {4'h0, dataGroup} == lastDataGroupReg;
  reg              hazardCheck;
  wire             accessBufferEnqueueFire;
  wire             vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_enq_ready = ~_vrfReadQueueVec_fifo_full | vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_deq_valid = ~_vrfReadQueueVec_fifo_empty | vrfReadQueueVec_0_enq_valid;
  wire [31:0]      vrfReadQueueVec_0_deq_bits = _vrfReadQueueVec_fifo_empty ? vrfReadQueueVec_0_enq_bits : _vrfReadQueueVec_fifo_data_out;
  wire             vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_enq_ready = ~_vrfReadQueueVec_fifo_1_full | vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_deq_valid = ~_vrfReadQueueVec_fifo_1_empty | vrfReadQueueVec_1_enq_valid;
  wire [31:0]      vrfReadQueueVec_1_deq_bits = _vrfReadQueueVec_fifo_1_empty ? vrfReadQueueVec_1_enq_bits : _vrfReadQueueVec_fifo_1_data_out;
  wire             vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_enq_ready = ~_vrfReadQueueVec_fifo_2_full | vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_deq_valid = ~_vrfReadQueueVec_fifo_2_empty | vrfReadQueueVec_2_enq_valid;
  wire [31:0]      vrfReadQueueVec_2_deq_bits = _vrfReadQueueVec_fifo_2_empty ? vrfReadQueueVec_2_enq_bits : _vrfReadQueueVec_fifo_2_data_out;
  wire             vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_enq_ready = ~_vrfReadQueueVec_fifo_3_full | vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_deq_valid = ~_vrfReadQueueVec_fifo_3_empty | vrfReadQueueVec_3_enq_valid;
  wire [31:0]      vrfReadQueueVec_3_deq_bits = _vrfReadQueueVec_fifo_3_empty ? vrfReadQueueVec_3_enq_bits : _vrfReadQueueVec_fifo_3_data_out;
  wire             vrfReadQueueVec_4_deq_ready;
  wire             vrfReadQueueVec_4_enq_ready = ~_vrfReadQueueVec_fifo_4_full | vrfReadQueueVec_4_deq_ready;
  wire             vrfReadQueueVec_4_deq_valid = ~_vrfReadQueueVec_fifo_4_empty | vrfReadQueueVec_4_enq_valid;
  wire [31:0]      vrfReadQueueVec_4_deq_bits = _vrfReadQueueVec_fifo_4_empty ? vrfReadQueueVec_4_enq_bits : _vrfReadQueueVec_fifo_4_data_out;
  wire             vrfReadQueueVec_5_deq_ready;
  wire             vrfReadQueueVec_5_enq_ready = ~_vrfReadQueueVec_fifo_5_full | vrfReadQueueVec_5_deq_ready;
  wire             vrfReadQueueVec_5_deq_valid = ~_vrfReadQueueVec_fifo_5_empty | vrfReadQueueVec_5_enq_valid;
  wire [31:0]      vrfReadQueueVec_5_deq_bits = _vrfReadQueueVec_fifo_5_empty ? vrfReadQueueVec_5_enq_bits : _vrfReadQueueVec_fifo_5_data_out;
  wire             vrfReadQueueVec_6_deq_ready;
  wire             vrfReadQueueVec_6_enq_ready = ~_vrfReadQueueVec_fifo_6_full | vrfReadQueueVec_6_deq_ready;
  wire             vrfReadQueueVec_6_deq_valid = ~_vrfReadQueueVec_fifo_6_empty | vrfReadQueueVec_6_enq_valid;
  wire [31:0]      vrfReadQueueVec_6_deq_bits = _vrfReadQueueVec_fifo_6_empty ? vrfReadQueueVec_6_enq_bits : _vrfReadQueueVec_fifo_6_data_out;
  wire             vrfReadQueueVec_7_deq_ready;
  wire             vrfReadQueueVec_7_enq_ready = ~_vrfReadQueueVec_fifo_7_full | vrfReadQueueVec_7_deq_ready;
  wire             vrfReadQueueVec_7_deq_valid = ~_vrfReadQueueVec_fifo_7_empty | vrfReadQueueVec_7_enq_valid;
  wire [31:0]      vrfReadQueueVec_7_deq_bits = _vrfReadQueueVec_fifo_7_empty ? vrfReadQueueVec_7_enq_bits : _vrfReadQueueVec_fifo_7_data_out;
  wire             vrfReadQueueVec_8_deq_ready;
  wire             vrfReadQueueVec_8_enq_ready = ~_vrfReadQueueVec_fifo_8_full | vrfReadQueueVec_8_deq_ready;
  wire             vrfReadQueueVec_8_deq_valid = ~_vrfReadQueueVec_fifo_8_empty | vrfReadQueueVec_8_enq_valid;
  wire [31:0]      vrfReadQueueVec_8_deq_bits = _vrfReadQueueVec_fifo_8_empty ? vrfReadQueueVec_8_enq_bits : _vrfReadQueueVec_fifo_8_data_out;
  wire             vrfReadQueueVec_9_deq_ready;
  wire             vrfReadQueueVec_9_enq_ready = ~_vrfReadQueueVec_fifo_9_full | vrfReadQueueVec_9_deq_ready;
  wire             vrfReadQueueVec_9_deq_valid = ~_vrfReadQueueVec_fifo_9_empty | vrfReadQueueVec_9_enq_valid;
  wire [31:0]      vrfReadQueueVec_9_deq_bits = _vrfReadQueueVec_fifo_9_empty ? vrfReadQueueVec_9_enq_bits : _vrfReadQueueVec_fifo_9_data_out;
  wire             vrfReadQueueVec_10_deq_ready;
  wire             vrfReadQueueVec_10_enq_ready = ~_vrfReadQueueVec_fifo_10_full | vrfReadQueueVec_10_deq_ready;
  wire             vrfReadQueueVec_10_deq_valid = ~_vrfReadQueueVec_fifo_10_empty | vrfReadQueueVec_10_enq_valid;
  wire [31:0]      vrfReadQueueVec_10_deq_bits = _vrfReadQueueVec_fifo_10_empty ? vrfReadQueueVec_10_enq_bits : _vrfReadQueueVec_fifo_10_data_out;
  wire             vrfReadQueueVec_11_deq_ready;
  wire             vrfReadQueueVec_11_enq_ready = ~_vrfReadQueueVec_fifo_11_full | vrfReadQueueVec_11_deq_ready;
  wire             vrfReadQueueVec_11_deq_valid = ~_vrfReadQueueVec_fifo_11_empty | vrfReadQueueVec_11_enq_valid;
  wire [31:0]      vrfReadQueueVec_11_deq_bits = _vrfReadQueueVec_fifo_11_empty ? vrfReadQueueVec_11_enq_bits : _vrfReadQueueVec_fifo_11_data_out;
  wire             vrfReadQueueVec_12_deq_ready;
  wire             vrfReadQueueVec_12_enq_ready = ~_vrfReadQueueVec_fifo_12_full | vrfReadQueueVec_12_deq_ready;
  wire             vrfReadQueueVec_12_deq_valid = ~_vrfReadQueueVec_fifo_12_empty | vrfReadQueueVec_12_enq_valid;
  wire [31:0]      vrfReadQueueVec_12_deq_bits = _vrfReadQueueVec_fifo_12_empty ? vrfReadQueueVec_12_enq_bits : _vrfReadQueueVec_fifo_12_data_out;
  wire             vrfReadQueueVec_13_deq_ready;
  wire             vrfReadQueueVec_13_enq_ready = ~_vrfReadQueueVec_fifo_13_full | vrfReadQueueVec_13_deq_ready;
  wire             vrfReadQueueVec_13_deq_valid = ~_vrfReadQueueVec_fifo_13_empty | vrfReadQueueVec_13_enq_valid;
  wire [31:0]      vrfReadQueueVec_13_deq_bits = _vrfReadQueueVec_fifo_13_empty ? vrfReadQueueVec_13_enq_bits : _vrfReadQueueVec_fifo_13_data_out;
  wire             vrfReadQueueVec_14_deq_ready;
  wire             vrfReadQueueVec_14_enq_ready = ~_vrfReadQueueVec_fifo_14_full | vrfReadQueueVec_14_deq_ready;
  wire             vrfReadQueueVec_14_deq_valid = ~_vrfReadQueueVec_fifo_14_empty | vrfReadQueueVec_14_enq_valid;
  wire [31:0]      vrfReadQueueVec_14_deq_bits = _vrfReadQueueVec_fifo_14_empty ? vrfReadQueueVec_14_enq_bits : _vrfReadQueueVec_fifo_14_data_out;
  wire             vrfReadQueueVec_15_deq_ready;
  wire             vrfReadQueueVec_15_enq_ready = ~_vrfReadQueueVec_fifo_15_full | vrfReadQueueVec_15_deq_ready;
  wire             vrfReadQueueVec_15_deq_valid = ~_vrfReadQueueVec_fifo_15_empty | vrfReadQueueVec_15_enq_valid;
  wire [31:0]      vrfReadQueueVec_15_deq_bits = _vrfReadQueueVec_fifo_15_empty ? vrfReadQueueVec_15_enq_bits : _vrfReadQueueVec_fifo_15_data_out;
  reg  [2:0]       readStageValid_segPtr;
  reg  [4:0]       readStageValid_readCount;
  reg              readStageValid_stageValid;
  wire             readStageValid_lastReadPtr = readStageValid_segPtr == 3'h0;
  wire [4:0]       readStageValid_nextReadCount = lsuRequest_valid ? 5'h0 : readStageValid_readCount + 5'h1;
  wire             readStageValid_lastReadGroup = {4'h0, readStageValid_readCount} == lastDataGroupReg;
  wire             vrfReadDataPorts_0_valid_0;
  wire             _readStageValid_T_11 = vrfReadDataPorts_0_ready_0 & vrfReadDataPorts_0_valid_0;
  reg  [3:0]       readStageValid_readCounter;
  wire [3:0]       readStageValid_counterChange = _readStageValid_T_11 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_0_valid_0 = readStageValid_stageValid & ~(readStageValid_readCounter[3]);
  wire [4:0]       _GEN_4 = {1'h0, segmentInstructionIndexInterval};
  wire [4:0]       vrfReadDataPorts_0_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr} * _GEN_4 + {2'h0, readStageValid_readCount[4:2]};
  wire [1:0]       vrfReadDataPorts_0_bits_offset_0 = readStageValid_readCount[1:0];
  reg  [2:0]       readStageValid_segPtr_1;
  reg  [4:0]       readStageValid_readCount_1;
  reg              readStageValid_stageValid_1;
  wire             readStageValid_lastReadPtr_1 = readStageValid_segPtr_1 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_1 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_1 + 5'h1;
  wire             readStageValid_lastReadGroup_1 = {4'h0, readStageValid_readCount_1} == lastDataGroupReg;
  wire             vrfReadDataPorts_1_valid_0;
  wire             _readStageValid_T_30 = vrfReadDataPorts_1_ready_0 & vrfReadDataPorts_1_valid_0;
  reg  [3:0]       readStageValid_readCounter_1;
  wire [3:0]       readStageValid_counterChange_1 = _readStageValid_T_30 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_1_valid_0 = readStageValid_stageValid_1 & ~(readStageValid_readCounter_1[3]);
  wire [4:0]       vrfReadDataPorts_1_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_1} * _GEN_4 + {2'h0, readStageValid_readCount_1[4:2]};
  wire [1:0]       vrfReadDataPorts_1_bits_offset_0 = readStageValid_readCount_1[1:0];
  reg  [2:0]       readStageValid_segPtr_2;
  reg  [4:0]       readStageValid_readCount_2;
  reg              readStageValid_stageValid_2;
  wire             readStageValid_lastReadPtr_2 = readStageValid_segPtr_2 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_2 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_2 + 5'h1;
  wire             readStageValid_lastReadGroup_2 = {4'h0, readStageValid_readCount_2} == lastDataGroupReg;
  wire             vrfReadDataPorts_2_valid_0;
  wire             _readStageValid_T_49 = vrfReadDataPorts_2_ready_0 & vrfReadDataPorts_2_valid_0;
  reg  [3:0]       readStageValid_readCounter_2;
  wire [3:0]       readStageValid_counterChange_2 = _readStageValid_T_49 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_2_valid_0 = readStageValid_stageValid_2 & ~(readStageValid_readCounter_2[3]);
  wire [4:0]       vrfReadDataPorts_2_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_2} * _GEN_4 + {2'h0, readStageValid_readCount_2[4:2]};
  wire [1:0]       vrfReadDataPorts_2_bits_offset_0 = readStageValid_readCount_2[1:0];
  reg  [2:0]       readStageValid_segPtr_3;
  reg  [4:0]       readStageValid_readCount_3;
  reg              readStageValid_stageValid_3;
  wire             readStageValid_lastReadPtr_3 = readStageValid_segPtr_3 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_3 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_3 + 5'h1;
  wire             readStageValid_lastReadGroup_3 = {4'h0, readStageValid_readCount_3} == lastDataGroupReg;
  wire             vrfReadDataPorts_3_valid_0;
  wire             _readStageValid_T_68 = vrfReadDataPorts_3_ready_0 & vrfReadDataPorts_3_valid_0;
  reg  [3:0]       readStageValid_readCounter_3;
  wire [3:0]       readStageValid_counterChange_3 = _readStageValid_T_68 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_3_valid_0 = readStageValid_stageValid_3 & ~(readStageValid_readCounter_3[3]);
  wire [4:0]       vrfReadDataPorts_3_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_3} * _GEN_4 + {2'h0, readStageValid_readCount_3[4:2]};
  wire [1:0]       vrfReadDataPorts_3_bits_offset_0 = readStageValid_readCount_3[1:0];
  reg  [2:0]       readStageValid_segPtr_4;
  reg  [4:0]       readStageValid_readCount_4;
  reg              readStageValid_stageValid_4;
  wire             readStageValid_lastReadPtr_4 = readStageValid_segPtr_4 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_4 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_4 + 5'h1;
  wire             readStageValid_lastReadGroup_4 = {4'h0, readStageValid_readCount_4} == lastDataGroupReg;
  wire             vrfReadDataPorts_4_valid_0;
  wire             _readStageValid_T_87 = vrfReadDataPorts_4_ready_0 & vrfReadDataPorts_4_valid_0;
  reg  [3:0]       readStageValid_readCounter_4;
  wire [3:0]       readStageValid_counterChange_4 = _readStageValid_T_87 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_4_valid_0 = readStageValid_stageValid_4 & ~(readStageValid_readCounter_4[3]);
  wire [4:0]       vrfReadDataPorts_4_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_4} * _GEN_4 + {2'h0, readStageValid_readCount_4[4:2]};
  wire [1:0]       vrfReadDataPorts_4_bits_offset_0 = readStageValid_readCount_4[1:0];
  reg  [2:0]       readStageValid_segPtr_5;
  reg  [4:0]       readStageValid_readCount_5;
  reg              readStageValid_stageValid_5;
  wire             readStageValid_lastReadPtr_5 = readStageValid_segPtr_5 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_5 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_5 + 5'h1;
  wire             readStageValid_lastReadGroup_5 = {4'h0, readStageValid_readCount_5} == lastDataGroupReg;
  wire             vrfReadDataPorts_5_valid_0;
  wire             _readStageValid_T_106 = vrfReadDataPorts_5_ready_0 & vrfReadDataPorts_5_valid_0;
  reg  [3:0]       readStageValid_readCounter_5;
  wire [3:0]       readStageValid_counterChange_5 = _readStageValid_T_106 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_5_valid_0 = readStageValid_stageValid_5 & ~(readStageValid_readCounter_5[3]);
  wire [4:0]       vrfReadDataPorts_5_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_5} * _GEN_4 + {2'h0, readStageValid_readCount_5[4:2]};
  wire [1:0]       vrfReadDataPorts_5_bits_offset_0 = readStageValid_readCount_5[1:0];
  reg  [2:0]       readStageValid_segPtr_6;
  reg  [4:0]       readStageValid_readCount_6;
  reg              readStageValid_stageValid_6;
  wire             readStageValid_lastReadPtr_6 = readStageValid_segPtr_6 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_6 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_6 + 5'h1;
  wire             readStageValid_lastReadGroup_6 = {4'h0, readStageValid_readCount_6} == lastDataGroupReg;
  wire             vrfReadDataPorts_6_valid_0;
  wire             _readStageValid_T_125 = vrfReadDataPorts_6_ready_0 & vrfReadDataPorts_6_valid_0;
  reg  [3:0]       readStageValid_readCounter_6;
  wire [3:0]       readStageValid_counterChange_6 = _readStageValid_T_125 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_6_valid_0 = readStageValid_stageValid_6 & ~(readStageValid_readCounter_6[3]);
  wire [4:0]       vrfReadDataPorts_6_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_6} * _GEN_4 + {2'h0, readStageValid_readCount_6[4:2]};
  wire [1:0]       vrfReadDataPorts_6_bits_offset_0 = readStageValid_readCount_6[1:0];
  reg  [2:0]       readStageValid_segPtr_7;
  reg  [4:0]       readStageValid_readCount_7;
  reg              readStageValid_stageValid_7;
  wire             readStageValid_lastReadPtr_7 = readStageValid_segPtr_7 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_7 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_7 + 5'h1;
  wire             readStageValid_lastReadGroup_7 = {4'h0, readStageValid_readCount_7} == lastDataGroupReg;
  wire             vrfReadDataPorts_7_valid_0;
  wire             _readStageValid_T_144 = vrfReadDataPorts_7_ready_0 & vrfReadDataPorts_7_valid_0;
  reg  [3:0]       readStageValid_readCounter_7;
  wire [3:0]       readStageValid_counterChange_7 = _readStageValid_T_144 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_7_valid_0 = readStageValid_stageValid_7 & ~(readStageValid_readCounter_7[3]);
  wire [4:0]       vrfReadDataPorts_7_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_7} * _GEN_4 + {2'h0, readStageValid_readCount_7[4:2]};
  wire [1:0]       vrfReadDataPorts_7_bits_offset_0 = readStageValid_readCount_7[1:0];
  reg  [2:0]       readStageValid_segPtr_8;
  reg  [4:0]       readStageValid_readCount_8;
  reg              readStageValid_stageValid_8;
  wire             readStageValid_lastReadPtr_8 = readStageValid_segPtr_8 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_8 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_8 + 5'h1;
  wire             readStageValid_lastReadGroup_8 = {4'h0, readStageValid_readCount_8} == lastDataGroupReg;
  wire             vrfReadDataPorts_8_valid_0;
  wire             _readStageValid_T_163 = vrfReadDataPorts_8_ready_0 & vrfReadDataPorts_8_valid_0;
  reg  [3:0]       readStageValid_readCounter_8;
  wire [3:0]       readStageValid_counterChange_8 = _readStageValid_T_163 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_8_valid_0 = readStageValid_stageValid_8 & ~(readStageValid_readCounter_8[3]);
  wire [4:0]       vrfReadDataPorts_8_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_8} * _GEN_4 + {2'h0, readStageValid_readCount_8[4:2]};
  wire [1:0]       vrfReadDataPorts_8_bits_offset_0 = readStageValid_readCount_8[1:0];
  reg  [2:0]       readStageValid_segPtr_9;
  reg  [4:0]       readStageValid_readCount_9;
  reg              readStageValid_stageValid_9;
  wire             readStageValid_lastReadPtr_9 = readStageValid_segPtr_9 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_9 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_9 + 5'h1;
  wire             readStageValid_lastReadGroup_9 = {4'h0, readStageValid_readCount_9} == lastDataGroupReg;
  wire             vrfReadDataPorts_9_valid_0;
  wire             _readStageValid_T_182 = vrfReadDataPorts_9_ready_0 & vrfReadDataPorts_9_valid_0;
  reg  [3:0]       readStageValid_readCounter_9;
  wire [3:0]       readStageValid_counterChange_9 = _readStageValid_T_182 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_9_valid_0 = readStageValid_stageValid_9 & ~(readStageValid_readCounter_9[3]);
  wire [4:0]       vrfReadDataPorts_9_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_9} * _GEN_4 + {2'h0, readStageValid_readCount_9[4:2]};
  wire [1:0]       vrfReadDataPorts_9_bits_offset_0 = readStageValid_readCount_9[1:0];
  reg  [2:0]       readStageValid_segPtr_10;
  reg  [4:0]       readStageValid_readCount_10;
  reg              readStageValid_stageValid_10;
  wire             readStageValid_lastReadPtr_10 = readStageValid_segPtr_10 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_10 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_10 + 5'h1;
  wire             readStageValid_lastReadGroup_10 = {4'h0, readStageValid_readCount_10} == lastDataGroupReg;
  wire             vrfReadDataPorts_10_valid_0;
  wire             _readStageValid_T_201 = vrfReadDataPorts_10_ready_0 & vrfReadDataPorts_10_valid_0;
  reg  [3:0]       readStageValid_readCounter_10;
  wire [3:0]       readStageValid_counterChange_10 = _readStageValid_T_201 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_10_valid_0 = readStageValid_stageValid_10 & ~(readStageValid_readCounter_10[3]);
  wire [4:0]       vrfReadDataPorts_10_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_10} * _GEN_4 + {2'h0, readStageValid_readCount_10[4:2]};
  wire [1:0]       vrfReadDataPorts_10_bits_offset_0 = readStageValid_readCount_10[1:0];
  reg  [2:0]       readStageValid_segPtr_11;
  reg  [4:0]       readStageValid_readCount_11;
  reg              readStageValid_stageValid_11;
  wire             readStageValid_lastReadPtr_11 = readStageValid_segPtr_11 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_11 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_11 + 5'h1;
  wire             readStageValid_lastReadGroup_11 = {4'h0, readStageValid_readCount_11} == lastDataGroupReg;
  wire             vrfReadDataPorts_11_valid_0;
  wire             _readStageValid_T_220 = vrfReadDataPorts_11_ready_0 & vrfReadDataPorts_11_valid_0;
  reg  [3:0]       readStageValid_readCounter_11;
  wire [3:0]       readStageValid_counterChange_11 = _readStageValid_T_220 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_11_valid_0 = readStageValid_stageValid_11 & ~(readStageValid_readCounter_11[3]);
  wire [4:0]       vrfReadDataPorts_11_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_11} * _GEN_4 + {2'h0, readStageValid_readCount_11[4:2]};
  wire [1:0]       vrfReadDataPorts_11_bits_offset_0 = readStageValid_readCount_11[1:0];
  reg  [2:0]       readStageValid_segPtr_12;
  reg  [4:0]       readStageValid_readCount_12;
  reg              readStageValid_stageValid_12;
  wire             readStageValid_lastReadPtr_12 = readStageValid_segPtr_12 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_12 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_12 + 5'h1;
  wire             readStageValid_lastReadGroup_12 = {4'h0, readStageValid_readCount_12} == lastDataGroupReg;
  wire             vrfReadDataPorts_12_valid_0;
  wire             _readStageValid_T_239 = vrfReadDataPorts_12_ready_0 & vrfReadDataPorts_12_valid_0;
  reg  [3:0]       readStageValid_readCounter_12;
  wire [3:0]       readStageValid_counterChange_12 = _readStageValid_T_239 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_12_valid_0 = readStageValid_stageValid_12 & ~(readStageValid_readCounter_12[3]);
  wire [4:0]       vrfReadDataPorts_12_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_12} * _GEN_4 + {2'h0, readStageValid_readCount_12[4:2]};
  wire [1:0]       vrfReadDataPorts_12_bits_offset_0 = readStageValid_readCount_12[1:0];
  reg  [2:0]       readStageValid_segPtr_13;
  reg  [4:0]       readStageValid_readCount_13;
  reg              readStageValid_stageValid_13;
  wire             readStageValid_lastReadPtr_13 = readStageValid_segPtr_13 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_13 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_13 + 5'h1;
  wire             readStageValid_lastReadGroup_13 = {4'h0, readStageValid_readCount_13} == lastDataGroupReg;
  wire             vrfReadDataPorts_13_valid_0;
  wire             _readStageValid_T_258 = vrfReadDataPorts_13_ready_0 & vrfReadDataPorts_13_valid_0;
  reg  [3:0]       readStageValid_readCounter_13;
  wire [3:0]       readStageValid_counterChange_13 = _readStageValid_T_258 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_13_valid_0 = readStageValid_stageValid_13 & ~(readStageValid_readCounter_13[3]);
  wire [4:0]       vrfReadDataPorts_13_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_13} * _GEN_4 + {2'h0, readStageValid_readCount_13[4:2]};
  wire [1:0]       vrfReadDataPorts_13_bits_offset_0 = readStageValid_readCount_13[1:0];
  reg  [2:0]       readStageValid_segPtr_14;
  reg  [4:0]       readStageValid_readCount_14;
  reg              readStageValid_stageValid_14;
  wire             readStageValid_lastReadPtr_14 = readStageValid_segPtr_14 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_14 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_14 + 5'h1;
  wire             readStageValid_lastReadGroup_14 = {4'h0, readStageValid_readCount_14} == lastDataGroupReg;
  wire             vrfReadDataPorts_14_valid_0;
  wire             _readStageValid_T_277 = vrfReadDataPorts_14_ready_0 & vrfReadDataPorts_14_valid_0;
  reg  [3:0]       readStageValid_readCounter_14;
  wire [3:0]       readStageValid_counterChange_14 = _readStageValid_T_277 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_14_valid_0 = readStageValid_stageValid_14 & ~(readStageValid_readCounter_14[3]);
  wire [4:0]       vrfReadDataPorts_14_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_14} * _GEN_4 + {2'h0, readStageValid_readCount_14[4:2]};
  wire [1:0]       vrfReadDataPorts_14_bits_offset_0 = readStageValid_readCount_14[1:0];
  reg  [2:0]       readStageValid_segPtr_15;
  reg  [4:0]       readStageValid_readCount_15;
  reg              readStageValid_stageValid_15;
  wire             readStageValid_lastReadPtr_15 = readStageValid_segPtr_15 == 3'h0;
  wire [4:0]       readStageValid_nextReadCount_15 = lsuRequest_valid ? 5'h0 : readStageValid_readCount_15 + 5'h1;
  wire             readStageValid_lastReadGroup_15 = {4'h0, readStageValid_readCount_15} == lastDataGroupReg;
  wire             vrfReadDataPorts_15_valid_0;
  wire             _readStageValid_T_296 = vrfReadDataPorts_15_ready_0 & vrfReadDataPorts_15_valid_0;
  reg  [3:0]       readStageValid_readCounter_15;
  wire [3:0]       readStageValid_counterChange_15 = _readStageValid_T_296 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_15_valid_0 = readStageValid_stageValid_15 & ~(readStageValid_readCounter_15[3]);
  wire [4:0]       vrfReadDataPorts_15_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_15} * _GEN_4 + {2'h0, readStageValid_readCount_15[4:2]};
  wire [1:0]       vrfReadDataPorts_15_bits_offset_0 = readStageValid_readCount_15[1:0];
  wire             readStageValid =
    |{readStageValid_stageValid,
      readStageValid_readCounter,
      readStageValid_stageValid_1,
      readStageValid_readCounter_1,
      readStageValid_stageValid_2,
      readStageValid_readCounter_2,
      readStageValid_stageValid_3,
      readStageValid_readCounter_3,
      readStageValid_stageValid_4,
      readStageValid_readCounter_4,
      readStageValid_stageValid_5,
      readStageValid_readCounter_5,
      readStageValid_stageValid_6,
      readStageValid_readCounter_6,
      readStageValid_stageValid_7,
      readStageValid_readCounter_7,
      readStageValid_stageValid_8,
      readStageValid_readCounter_8,
      readStageValid_stageValid_9,
      readStageValid_readCounter_9,
      readStageValid_stageValid_10,
      readStageValid_readCounter_10,
      readStageValid_stageValid_11,
      readStageValid_readCounter_11,
      readStageValid_stageValid_12,
      readStageValid_readCounter_12,
      readStageValid_stageValid_13,
      readStageValid_readCounter_13,
      readStageValid_stageValid_14,
      readStageValid_readCounter_14,
      readStageValid_stageValid_15,
      readStageValid_readCounter_15};
  reg              bufferFull;
  wire             accessBufferDequeueReady;
  wire             accessBufferEnqueueReady = ~bufferFull | accessBufferDequeueReady;
  wire             accessBufferEnqueueValid =
    vrfReadQueueVec_0_deq_valid & vrfReadQueueVec_1_deq_valid & vrfReadQueueVec_2_deq_valid & vrfReadQueueVec_3_deq_valid & vrfReadQueueVec_4_deq_valid & vrfReadQueueVec_5_deq_valid & vrfReadQueueVec_6_deq_valid
    & vrfReadQueueVec_7_deq_valid & vrfReadQueueVec_8_deq_valid & vrfReadQueueVec_9_deq_valid & vrfReadQueueVec_10_deq_valid & vrfReadQueueVec_11_deq_valid & vrfReadQueueVec_12_deq_valid & vrfReadQueueVec_13_deq_valid
    & vrfReadQueueVec_14_deq_valid & vrfReadQueueVec_15_deq_valid;
  wire             readQueueClear =
    ~(vrfReadQueueVec_0_deq_valid | vrfReadQueueVec_1_deq_valid | vrfReadQueueVec_2_deq_valid | vrfReadQueueVec_3_deq_valid | vrfReadQueueVec_4_deq_valid | vrfReadQueueVec_5_deq_valid | vrfReadQueueVec_6_deq_valid
      | vrfReadQueueVec_7_deq_valid | vrfReadQueueVec_8_deq_valid | vrfReadQueueVec_9_deq_valid | vrfReadQueueVec_10_deq_valid | vrfReadQueueVec_11_deq_valid | vrfReadQueueVec_12_deq_valid | vrfReadQueueVec_13_deq_valid
      | vrfReadQueueVec_14_deq_valid | vrfReadQueueVec_15_deq_valid);
  assign accessBufferEnqueueFire = accessBufferEnqueueValid & accessBufferEnqueueReady;
  assign vrfReadQueueVec_0_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_1_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_2_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_3_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_4_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_5_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_6_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_7_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_8_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_9_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_10_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_11_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_12_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_13_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_14_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_15_deq_ready = accessBufferEnqueueFire;
  wire             lastPtr = accessPtr == 3'h0;
  wire             lastPtrEnq = lastPtr & accessBufferEnqueueFire;
  wire             accessBufferDequeueValid = bufferFull | lastPtrEnq;
  wire             accessBufferDequeueFire = accessBufferDequeueValid & accessBufferDequeueReady;
  wire [63:0]      accessDataUpdate_lo_lo_lo = {vrfReadQueueVec_1_deq_bits, vrfReadQueueVec_0_deq_bits};
  wire [63:0]      accessDataUpdate_lo_lo_hi = {vrfReadQueueVec_3_deq_bits, vrfReadQueueVec_2_deq_bits};
  wire [127:0]     accessDataUpdate_lo_lo = {accessDataUpdate_lo_lo_hi, accessDataUpdate_lo_lo_lo};
  wire [63:0]      accessDataUpdate_lo_hi_lo = {vrfReadQueueVec_5_deq_bits, vrfReadQueueVec_4_deq_bits};
  wire [63:0]      accessDataUpdate_lo_hi_hi = {vrfReadQueueVec_7_deq_bits, vrfReadQueueVec_6_deq_bits};
  wire [127:0]     accessDataUpdate_lo_hi = {accessDataUpdate_lo_hi_hi, accessDataUpdate_lo_hi_lo};
  wire [255:0]     accessDataUpdate_lo = {accessDataUpdate_lo_hi, accessDataUpdate_lo_lo};
  wire [63:0]      accessDataUpdate_hi_lo_lo = {vrfReadQueueVec_9_deq_bits, vrfReadQueueVec_8_deq_bits};
  wire [63:0]      accessDataUpdate_hi_lo_hi = {vrfReadQueueVec_11_deq_bits, vrfReadQueueVec_10_deq_bits};
  wire [127:0]     accessDataUpdate_hi_lo = {accessDataUpdate_hi_lo_hi, accessDataUpdate_hi_lo_lo};
  wire [63:0]      accessDataUpdate_hi_hi_lo = {vrfReadQueueVec_13_deq_bits, vrfReadQueueVec_12_deq_bits};
  wire [63:0]      accessDataUpdate_hi_hi_hi = {vrfReadQueueVec_15_deq_bits, vrfReadQueueVec_14_deq_bits};
  wire [127:0]     accessDataUpdate_hi_hi = {accessDataUpdate_hi_hi_hi, accessDataUpdate_hi_hi_lo};
  wire [255:0]     accessDataUpdate_hi = {accessDataUpdate_hi_hi, accessDataUpdate_hi_lo};
  wire [511:0]     accessDataUpdate_0 = {accessDataUpdate_hi, accessDataUpdate_lo};
  reg              bufferValid;
  reg  [63:0]      maskForBufferData_0;
  reg  [63:0]      maskForBufferData_1;
  reg  [63:0]      maskForBufferData_2;
  reg  [63:0]      maskForBufferData_3;
  reg  [63:0]      maskForBufferData_4;
  reg  [63:0]      maskForBufferData_5;
  reg  [63:0]      maskForBufferData_6;
  reg  [63:0]      maskForBufferData_7;
  reg              lastDataGroupInDataBuffer;
  wire             memRequest_valid_0;
  wire             _addressQueue_enq_valid_T = memRequest_ready_0 & memRequest_valid_0;
  wire             alignedDequeueFire;
  assign alignedDequeueFire = _addressQueue_enq_valid_T;
  wire             addressQueue_enq_valid;
  assign addressQueue_enq_valid = _addressQueue_enq_valid_T;
  reg  [511:0]     cacheLineTemp;
  reg  [63:0]      maskTemp;
  reg              canSendTail;
  wire             isLastCacheLineInBuffer = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire             bufferWillClear = alignedDequeueFire & isLastCacheLineInBuffer;
  wire             addressQueue_enq_ready;
  wire             addressQueueFree;
  assign accessBufferDequeueReady = ~bufferValid | memRequest_ready_0 & isLastCacheLineInBuffer & addressQueueFree;
  wire [511:0]     bufferStageEnqueueData_0 = bufferFull ? accessData_0 : accessDataUpdate_0;
  wire [511:0]     bufferStageEnqueueData_1 = bufferFull ? accessData_1 : accessDataUpdate_1;
  wire [511:0]     bufferStageEnqueueData_2 = bufferFull ? accessData_2 : accessDataUpdate_2;
  wire [511:0]     bufferStageEnqueueData_3 = bufferFull ? accessData_3 : accessDataUpdate_3;
  wire [511:0]     bufferStageEnqueueData_4 = bufferFull ? accessData_4 : accessDataUpdate_4;
  wire [511:0]     bufferStageEnqueueData_5 = bufferFull ? accessData_5 : accessDataUpdate_5;
  wire [511:0]     bufferStageEnqueueData_6 = bufferFull ? accessData_6 : accessDataUpdate_6;
  wire [511:0]     bufferStageEnqueueData_7 = bufferFull ? accessData_7 : accessDataUpdate_7;
  wire [7:0]       _fillBySeg_T = 8'h1 << lsuRequestReg_instructionInformation_nf;
  wire [3:0]       fillBySeg_lo_lo_lo_lo = {fillBySeg_lo_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_lo_lo_hi = {fillBySeg_lo_lo_lo_hi_hi, fillBySeg_lo_lo_lo_hi_lo};
  wire [7:0]       fillBySeg_lo_lo_lo = {fillBySeg_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_lo_hi_lo = {fillBySeg_lo_lo_hi_lo_hi, fillBySeg_lo_lo_hi_lo_lo};
  wire [3:0]       fillBySeg_lo_lo_hi_hi = {fillBySeg_lo_lo_hi_hi_hi, fillBySeg_lo_lo_hi_hi_lo};
  wire [7:0]       fillBySeg_lo_lo_hi = {fillBySeg_lo_lo_hi_hi, fillBySeg_lo_lo_hi_lo};
  wire [15:0]      fillBySeg_lo_lo = {fillBySeg_lo_lo_hi, fillBySeg_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_lo_lo = {fillBySeg_lo_hi_lo_lo_hi, fillBySeg_lo_hi_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_lo_hi = {fillBySeg_lo_hi_lo_hi_hi, fillBySeg_lo_hi_lo_hi_lo};
  wire [7:0]       fillBySeg_lo_hi_lo = {fillBySeg_lo_hi_lo_hi, fillBySeg_lo_hi_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_hi_lo = {fillBySeg_lo_hi_hi_lo_hi, fillBySeg_lo_hi_hi_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_hi_hi = {fillBySeg_lo_hi_hi_hi_hi, fillBySeg_lo_hi_hi_hi_lo};
  wire [7:0]       fillBySeg_lo_hi_hi = {fillBySeg_lo_hi_hi_hi, fillBySeg_lo_hi_hi_lo};
  wire [15:0]      fillBySeg_lo_hi = {fillBySeg_lo_hi_hi, fillBySeg_lo_hi_lo};
  wire [31:0]      fillBySeg_lo = {fillBySeg_lo_hi, fillBySeg_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_lo_lo = {fillBySeg_hi_lo_lo_lo_hi, fillBySeg_hi_lo_lo_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_lo_hi = {fillBySeg_hi_lo_lo_hi_hi, fillBySeg_hi_lo_lo_hi_lo};
  wire [7:0]       fillBySeg_hi_lo_lo = {fillBySeg_hi_lo_lo_hi, fillBySeg_hi_lo_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_hi_lo = {fillBySeg_hi_lo_hi_lo_hi, fillBySeg_hi_lo_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_hi_hi = {fillBySeg_hi_lo_hi_hi_hi, fillBySeg_hi_lo_hi_hi_lo};
  wire [7:0]       fillBySeg_hi_lo_hi = {fillBySeg_hi_lo_hi_hi, fillBySeg_hi_lo_hi_lo};
  wire [15:0]      fillBySeg_hi_lo = {fillBySeg_hi_lo_hi, fillBySeg_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_lo_lo = {fillBySeg_hi_hi_lo_lo_hi, fillBySeg_hi_hi_lo_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_lo_hi = {fillBySeg_hi_hi_lo_hi_hi, fillBySeg_hi_hi_lo_hi_lo};
  wire [7:0]       fillBySeg_hi_hi_lo = {fillBySeg_hi_hi_lo_hi, fillBySeg_hi_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_hi_lo = {fillBySeg_hi_hi_hi_lo_hi, fillBySeg_hi_hi_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_hi_hi = {fillBySeg_hi_hi_hi_hi_hi, fillBySeg_hi_hi_hi_hi_lo};
  wire [7:0]       fillBySeg_hi_hi_hi = {fillBySeg_hi_hi_hi_hi, fillBySeg_hi_hi_hi_lo};
  wire [15:0]      fillBySeg_hi_hi = {fillBySeg_hi_hi_hi, fillBySeg_hi_hi_lo};
  wire [31:0]      fillBySeg_hi = {fillBySeg_hi_hi, fillBySeg_hi_lo};
  wire [3:0]       fillBySeg_lo_lo_lo_lo_lo_1 = {{2{maskForGroupWire[1]}}, {2{maskForGroupWire[0]}}};
  wire [3:0]       fillBySeg_lo_lo_lo_lo_hi_1 = {{2{maskForGroupWire[3]}}, {2{maskForGroupWire[2]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_lo_lo_hi_lo_1 = {{2{maskForGroupWire[5]}}, {2{maskForGroupWire[4]}}};
  wire [3:0]       fillBySeg_lo_lo_lo_hi_hi_1 = {{2{maskForGroupWire[7]}}, {2{maskForGroupWire[6]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_hi_1 = {fillBySeg_lo_lo_lo_hi_hi_1, fillBySeg_lo_lo_lo_hi_lo_1};
  wire [15:0]      fillBySeg_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_lo_hi_lo_lo_1 = {{2{maskForGroupWire[9]}}, {2{maskForGroupWire[8]}}};
  wire [3:0]       fillBySeg_lo_lo_hi_lo_hi_1 = {{2{maskForGroupWire[11]}}, {2{maskForGroupWire[10]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_lo_1 = {fillBySeg_lo_lo_hi_lo_hi_1, fillBySeg_lo_lo_hi_lo_lo_1};
  wire [3:0]       fillBySeg_lo_lo_hi_hi_lo_1 = {{2{maskForGroupWire[13]}}, {2{maskForGroupWire[12]}}};
  wire [3:0]       fillBySeg_lo_lo_hi_hi_hi_1 = {{2{maskForGroupWire[15]}}, {2{maskForGroupWire[14]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_hi_1 = {fillBySeg_lo_lo_hi_hi_hi_1, fillBySeg_lo_lo_hi_hi_lo_1};
  wire [15:0]      fillBySeg_lo_lo_hi_1 = {fillBySeg_lo_lo_hi_hi_1, fillBySeg_lo_lo_hi_lo_1};
  wire [31:0]      fillBySeg_lo_lo_1 = {fillBySeg_lo_lo_hi_1, fillBySeg_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_lo_lo_lo_1 = {{2{maskForGroupWire[17]}}, {2{maskForGroupWire[16]}}};
  wire [3:0]       fillBySeg_lo_hi_lo_lo_hi_1 = {{2{maskForGroupWire[19]}}, {2{maskForGroupWire[18]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_lo_1 = {fillBySeg_lo_hi_lo_lo_hi_1, fillBySeg_lo_hi_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_lo_hi_lo_1 = {{2{maskForGroupWire[21]}}, {2{maskForGroupWire[20]}}};
  wire [3:0]       fillBySeg_lo_hi_lo_hi_hi_1 = {{2{maskForGroupWire[23]}}, {2{maskForGroupWire[22]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_hi_1 = {fillBySeg_lo_hi_lo_hi_hi_1, fillBySeg_lo_hi_lo_hi_lo_1};
  wire [15:0]      fillBySeg_lo_hi_lo_1 = {fillBySeg_lo_hi_lo_hi_1, fillBySeg_lo_hi_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_hi_lo_lo_1 = {{2{maskForGroupWire[25]}}, {2{maskForGroupWire[24]}}};
  wire [3:0]       fillBySeg_lo_hi_hi_lo_hi_1 = {{2{maskForGroupWire[27]}}, {2{maskForGroupWire[26]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_lo_1 = {fillBySeg_lo_hi_hi_lo_hi_1, fillBySeg_lo_hi_hi_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_hi_hi_lo_1 = {{2{maskForGroupWire[29]}}, {2{maskForGroupWire[28]}}};
  wire [3:0]       fillBySeg_lo_hi_hi_hi_hi_1 = {{2{maskForGroupWire[31]}}, {2{maskForGroupWire[30]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_hi_1, fillBySeg_lo_hi_hi_hi_lo_1};
  wire [15:0]      fillBySeg_lo_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_1, fillBySeg_lo_hi_hi_lo_1};
  wire [31:0]      fillBySeg_lo_hi_1 = {fillBySeg_lo_hi_hi_1, fillBySeg_lo_hi_lo_1};
  wire [63:0]      fillBySeg_lo_1 = {fillBySeg_lo_hi_1, fillBySeg_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_lo_lo_lo_1 = {{2{maskForGroupWire[33]}}, {2{maskForGroupWire[32]}}};
  wire [3:0]       fillBySeg_hi_lo_lo_lo_hi_1 = {{2{maskForGroupWire[35]}}, {2{maskForGroupWire[34]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_lo_1 = {fillBySeg_hi_lo_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_lo_hi_lo_1 = {{2{maskForGroupWire[37]}}, {2{maskForGroupWire[36]}}};
  wire [3:0]       fillBySeg_hi_lo_lo_hi_hi_1 = {{2{maskForGroupWire[39]}}, {2{maskForGroupWire[38]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_hi_1 = {fillBySeg_hi_lo_lo_hi_hi_1, fillBySeg_hi_lo_lo_hi_lo_1};
  wire [15:0]      fillBySeg_hi_lo_lo_1 = {fillBySeg_hi_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_hi_lo_lo_1 = {{2{maskForGroupWire[41]}}, {2{maskForGroupWire[40]}}};
  wire [3:0]       fillBySeg_hi_lo_hi_lo_hi_1 = {{2{maskForGroupWire[43]}}, {2{maskForGroupWire[42]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_lo_1 = {fillBySeg_hi_lo_hi_lo_hi_1, fillBySeg_hi_lo_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_hi_hi_lo_1 = {{2{maskForGroupWire[45]}}, {2{maskForGroupWire[44]}}};
  wire [3:0]       fillBySeg_hi_lo_hi_hi_hi_1 = {{2{maskForGroupWire[47]}}, {2{maskForGroupWire[46]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_hi_1 = {fillBySeg_hi_lo_hi_hi_hi_1, fillBySeg_hi_lo_hi_hi_lo_1};
  wire [15:0]      fillBySeg_hi_lo_hi_1 = {fillBySeg_hi_lo_hi_hi_1, fillBySeg_hi_lo_hi_lo_1};
  wire [31:0]      fillBySeg_hi_lo_1 = {fillBySeg_hi_lo_hi_1, fillBySeg_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_lo_lo_lo_1 = {{2{maskForGroupWire[49]}}, {2{maskForGroupWire[48]}}};
  wire [3:0]       fillBySeg_hi_hi_lo_lo_hi_1 = {{2{maskForGroupWire[51]}}, {2{maskForGroupWire[50]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_lo_1 = {fillBySeg_hi_hi_lo_lo_hi_1, fillBySeg_hi_hi_lo_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_lo_hi_lo_1 = {{2{maskForGroupWire[53]}}, {2{maskForGroupWire[52]}}};
  wire [3:0]       fillBySeg_hi_hi_lo_hi_hi_1 = {{2{maskForGroupWire[55]}}, {2{maskForGroupWire[54]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_hi_1 = {fillBySeg_hi_hi_lo_hi_hi_1, fillBySeg_hi_hi_lo_hi_lo_1};
  wire [15:0]      fillBySeg_hi_hi_lo_1 = {fillBySeg_hi_hi_lo_hi_1, fillBySeg_hi_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_hi_lo_lo_1 = {{2{maskForGroupWire[57]}}, {2{maskForGroupWire[56]}}};
  wire [3:0]       fillBySeg_hi_hi_hi_lo_hi_1 = {{2{maskForGroupWire[59]}}, {2{maskForGroupWire[58]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_lo_1 = {fillBySeg_hi_hi_hi_lo_hi_1, fillBySeg_hi_hi_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_hi_hi_lo_1 = {{2{maskForGroupWire[61]}}, {2{maskForGroupWire[60]}}};
  wire [3:0]       fillBySeg_hi_hi_hi_hi_hi_1 = {{2{maskForGroupWire[63]}}, {2{maskForGroupWire[62]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_hi_lo_1};
  wire [15:0]      fillBySeg_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_lo_1};
  wire [31:0]      fillBySeg_hi_hi_1 = {fillBySeg_hi_hi_hi_1, fillBySeg_hi_hi_lo_1};
  wire [63:0]      fillBySeg_hi_1 = {fillBySeg_hi_hi_1, fillBySeg_hi_lo_1};
  wire [5:0]       fillBySeg_lo_lo_lo_lo_lo_2 = {{3{maskForGroupWire[1]}}, {3{maskForGroupWire[0]}}};
  wire [5:0]       fillBySeg_lo_lo_lo_lo_hi_2 = {{3{maskForGroupWire[3]}}, {3{maskForGroupWire[2]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_lo_lo_hi_lo_2 = {{3{maskForGroupWire[5]}}, {3{maskForGroupWire[4]}}};
  wire [5:0]       fillBySeg_lo_lo_lo_hi_hi_2 = {{3{maskForGroupWire[7]}}, {3{maskForGroupWire[6]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_hi_2 = {fillBySeg_lo_lo_lo_hi_hi_2, fillBySeg_lo_lo_lo_hi_lo_2};
  wire [23:0]      fillBySeg_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_lo_hi_lo_lo_2 = {{3{maskForGroupWire[9]}}, {3{maskForGroupWire[8]}}};
  wire [5:0]       fillBySeg_lo_lo_hi_lo_hi_2 = {{3{maskForGroupWire[11]}}, {3{maskForGroupWire[10]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_lo_2 = {fillBySeg_lo_lo_hi_lo_hi_2, fillBySeg_lo_lo_hi_lo_lo_2};
  wire [5:0]       fillBySeg_lo_lo_hi_hi_lo_2 = {{3{maskForGroupWire[13]}}, {3{maskForGroupWire[12]}}};
  wire [5:0]       fillBySeg_lo_lo_hi_hi_hi_2 = {{3{maskForGroupWire[15]}}, {3{maskForGroupWire[14]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_hi_2 = {fillBySeg_lo_lo_hi_hi_hi_2, fillBySeg_lo_lo_hi_hi_lo_2};
  wire [23:0]      fillBySeg_lo_lo_hi_2 = {fillBySeg_lo_lo_hi_hi_2, fillBySeg_lo_lo_hi_lo_2};
  wire [47:0]      fillBySeg_lo_lo_2 = {fillBySeg_lo_lo_hi_2, fillBySeg_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_lo_lo_lo_2 = {{3{maskForGroupWire[17]}}, {3{maskForGroupWire[16]}}};
  wire [5:0]       fillBySeg_lo_hi_lo_lo_hi_2 = {{3{maskForGroupWire[19]}}, {3{maskForGroupWire[18]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_lo_2 = {fillBySeg_lo_hi_lo_lo_hi_2, fillBySeg_lo_hi_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_lo_hi_lo_2 = {{3{maskForGroupWire[21]}}, {3{maskForGroupWire[20]}}};
  wire [5:0]       fillBySeg_lo_hi_lo_hi_hi_2 = {{3{maskForGroupWire[23]}}, {3{maskForGroupWire[22]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_hi_2 = {fillBySeg_lo_hi_lo_hi_hi_2, fillBySeg_lo_hi_lo_hi_lo_2};
  wire [23:0]      fillBySeg_lo_hi_lo_2 = {fillBySeg_lo_hi_lo_hi_2, fillBySeg_lo_hi_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_hi_lo_lo_2 = {{3{maskForGroupWire[25]}}, {3{maskForGroupWire[24]}}};
  wire [5:0]       fillBySeg_lo_hi_hi_lo_hi_2 = {{3{maskForGroupWire[27]}}, {3{maskForGroupWire[26]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_lo_2 = {fillBySeg_lo_hi_hi_lo_hi_2, fillBySeg_lo_hi_hi_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_hi_hi_lo_2 = {{3{maskForGroupWire[29]}}, {3{maskForGroupWire[28]}}};
  wire [5:0]       fillBySeg_lo_hi_hi_hi_hi_2 = {{3{maskForGroupWire[31]}}, {3{maskForGroupWire[30]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_hi_2, fillBySeg_lo_hi_hi_hi_lo_2};
  wire [23:0]      fillBySeg_lo_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_2, fillBySeg_lo_hi_hi_lo_2};
  wire [47:0]      fillBySeg_lo_hi_2 = {fillBySeg_lo_hi_hi_2, fillBySeg_lo_hi_lo_2};
  wire [95:0]      fillBySeg_lo_2 = {fillBySeg_lo_hi_2, fillBySeg_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_lo_lo_lo_2 = {{3{maskForGroupWire[33]}}, {3{maskForGroupWire[32]}}};
  wire [5:0]       fillBySeg_hi_lo_lo_lo_hi_2 = {{3{maskForGroupWire[35]}}, {3{maskForGroupWire[34]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_lo_2 = {fillBySeg_hi_lo_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_lo_hi_lo_2 = {{3{maskForGroupWire[37]}}, {3{maskForGroupWire[36]}}};
  wire [5:0]       fillBySeg_hi_lo_lo_hi_hi_2 = {{3{maskForGroupWire[39]}}, {3{maskForGroupWire[38]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_hi_2 = {fillBySeg_hi_lo_lo_hi_hi_2, fillBySeg_hi_lo_lo_hi_lo_2};
  wire [23:0]      fillBySeg_hi_lo_lo_2 = {fillBySeg_hi_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_hi_lo_lo_2 = {{3{maskForGroupWire[41]}}, {3{maskForGroupWire[40]}}};
  wire [5:0]       fillBySeg_hi_lo_hi_lo_hi_2 = {{3{maskForGroupWire[43]}}, {3{maskForGroupWire[42]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_lo_2 = {fillBySeg_hi_lo_hi_lo_hi_2, fillBySeg_hi_lo_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_hi_hi_lo_2 = {{3{maskForGroupWire[45]}}, {3{maskForGroupWire[44]}}};
  wire [5:0]       fillBySeg_hi_lo_hi_hi_hi_2 = {{3{maskForGroupWire[47]}}, {3{maskForGroupWire[46]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_hi_2 = {fillBySeg_hi_lo_hi_hi_hi_2, fillBySeg_hi_lo_hi_hi_lo_2};
  wire [23:0]      fillBySeg_hi_lo_hi_2 = {fillBySeg_hi_lo_hi_hi_2, fillBySeg_hi_lo_hi_lo_2};
  wire [47:0]      fillBySeg_hi_lo_2 = {fillBySeg_hi_lo_hi_2, fillBySeg_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_lo_lo_lo_2 = {{3{maskForGroupWire[49]}}, {3{maskForGroupWire[48]}}};
  wire [5:0]       fillBySeg_hi_hi_lo_lo_hi_2 = {{3{maskForGroupWire[51]}}, {3{maskForGroupWire[50]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_lo_2 = {fillBySeg_hi_hi_lo_lo_hi_2, fillBySeg_hi_hi_lo_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_lo_hi_lo_2 = {{3{maskForGroupWire[53]}}, {3{maskForGroupWire[52]}}};
  wire [5:0]       fillBySeg_hi_hi_lo_hi_hi_2 = {{3{maskForGroupWire[55]}}, {3{maskForGroupWire[54]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_hi_2 = {fillBySeg_hi_hi_lo_hi_hi_2, fillBySeg_hi_hi_lo_hi_lo_2};
  wire [23:0]      fillBySeg_hi_hi_lo_2 = {fillBySeg_hi_hi_lo_hi_2, fillBySeg_hi_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_hi_lo_lo_2 = {{3{maskForGroupWire[57]}}, {3{maskForGroupWire[56]}}};
  wire [5:0]       fillBySeg_hi_hi_hi_lo_hi_2 = {{3{maskForGroupWire[59]}}, {3{maskForGroupWire[58]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_lo_2 = {fillBySeg_hi_hi_hi_lo_hi_2, fillBySeg_hi_hi_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_hi_hi_lo_2 = {{3{maskForGroupWire[61]}}, {3{maskForGroupWire[60]}}};
  wire [5:0]       fillBySeg_hi_hi_hi_hi_hi_2 = {{3{maskForGroupWire[63]}}, {3{maskForGroupWire[62]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_hi_lo_2};
  wire [23:0]      fillBySeg_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_lo_2};
  wire [47:0]      fillBySeg_hi_hi_2 = {fillBySeg_hi_hi_hi_2, fillBySeg_hi_hi_lo_2};
  wire [95:0]      fillBySeg_hi_2 = {fillBySeg_hi_hi_2, fillBySeg_hi_lo_2};
  wire [7:0]       fillBySeg_lo_lo_lo_lo_lo_3 = {{4{maskForGroupWire[1]}}, {4{maskForGroupWire[0]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_lo_hi_3 = {{4{maskForGroupWire[3]}}, {4{maskForGroupWire[2]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_lo_lo_hi_lo_3 = {{4{maskForGroupWire[5]}}, {4{maskForGroupWire[4]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_hi_hi_3 = {{4{maskForGroupWire[7]}}, {4{maskForGroupWire[6]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_hi_3 = {fillBySeg_lo_lo_lo_hi_hi_3, fillBySeg_lo_lo_lo_hi_lo_3};
  wire [31:0]      fillBySeg_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_lo_hi_lo_lo_3 = {{4{maskForGroupWire[9]}}, {4{maskForGroupWire[8]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_lo_hi_3 = {{4{maskForGroupWire[11]}}, {4{maskForGroupWire[10]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_lo_3 = {fillBySeg_lo_lo_hi_lo_hi_3, fillBySeg_lo_lo_hi_lo_lo_3};
  wire [7:0]       fillBySeg_lo_lo_hi_hi_lo_3 = {{4{maskForGroupWire[13]}}, {4{maskForGroupWire[12]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_hi_hi_3 = {{4{maskForGroupWire[15]}}, {4{maskForGroupWire[14]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_hi_3 = {fillBySeg_lo_lo_hi_hi_hi_3, fillBySeg_lo_lo_hi_hi_lo_3};
  wire [31:0]      fillBySeg_lo_lo_hi_3 = {fillBySeg_lo_lo_hi_hi_3, fillBySeg_lo_lo_hi_lo_3};
  wire [63:0]      fillBySeg_lo_lo_3 = {fillBySeg_lo_lo_hi_3, fillBySeg_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_lo_lo_lo_3 = {{4{maskForGroupWire[17]}}, {4{maskForGroupWire[16]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_lo_hi_3 = {{4{maskForGroupWire[19]}}, {4{maskForGroupWire[18]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_lo_3 = {fillBySeg_lo_hi_lo_lo_hi_3, fillBySeg_lo_hi_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_lo_hi_lo_3 = {{4{maskForGroupWire[21]}}, {4{maskForGroupWire[20]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_hi_hi_3 = {{4{maskForGroupWire[23]}}, {4{maskForGroupWire[22]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_hi_3 = {fillBySeg_lo_hi_lo_hi_hi_3, fillBySeg_lo_hi_lo_hi_lo_3};
  wire [31:0]      fillBySeg_lo_hi_lo_3 = {fillBySeg_lo_hi_lo_hi_3, fillBySeg_lo_hi_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_hi_lo_lo_3 = {{4{maskForGroupWire[25]}}, {4{maskForGroupWire[24]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_lo_hi_3 = {{4{maskForGroupWire[27]}}, {4{maskForGroupWire[26]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_lo_3 = {fillBySeg_lo_hi_hi_lo_hi_3, fillBySeg_lo_hi_hi_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_hi_hi_lo_3 = {{4{maskForGroupWire[29]}}, {4{maskForGroupWire[28]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_hi_hi_3 = {{4{maskForGroupWire[31]}}, {4{maskForGroupWire[30]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_hi_3, fillBySeg_lo_hi_hi_hi_lo_3};
  wire [31:0]      fillBySeg_lo_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_3, fillBySeg_lo_hi_hi_lo_3};
  wire [63:0]      fillBySeg_lo_hi_3 = {fillBySeg_lo_hi_hi_3, fillBySeg_lo_hi_lo_3};
  wire [127:0]     fillBySeg_lo_3 = {fillBySeg_lo_hi_3, fillBySeg_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_lo_lo_lo_3 = {{4{maskForGroupWire[33]}}, {4{maskForGroupWire[32]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_lo_hi_3 = {{4{maskForGroupWire[35]}}, {4{maskForGroupWire[34]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_lo_3 = {fillBySeg_hi_lo_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_lo_hi_lo_3 = {{4{maskForGroupWire[37]}}, {4{maskForGroupWire[36]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_hi_hi_3 = {{4{maskForGroupWire[39]}}, {4{maskForGroupWire[38]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_hi_3 = {fillBySeg_hi_lo_lo_hi_hi_3, fillBySeg_hi_lo_lo_hi_lo_3};
  wire [31:0]      fillBySeg_hi_lo_lo_3 = {fillBySeg_hi_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_hi_lo_lo_3 = {{4{maskForGroupWire[41]}}, {4{maskForGroupWire[40]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_lo_hi_3 = {{4{maskForGroupWire[43]}}, {4{maskForGroupWire[42]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_lo_3 = {fillBySeg_hi_lo_hi_lo_hi_3, fillBySeg_hi_lo_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_hi_hi_lo_3 = {{4{maskForGroupWire[45]}}, {4{maskForGroupWire[44]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_hi_hi_3 = {{4{maskForGroupWire[47]}}, {4{maskForGroupWire[46]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_hi_3 = {fillBySeg_hi_lo_hi_hi_hi_3, fillBySeg_hi_lo_hi_hi_lo_3};
  wire [31:0]      fillBySeg_hi_lo_hi_3 = {fillBySeg_hi_lo_hi_hi_3, fillBySeg_hi_lo_hi_lo_3};
  wire [63:0]      fillBySeg_hi_lo_3 = {fillBySeg_hi_lo_hi_3, fillBySeg_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_lo_lo_lo_3 = {{4{maskForGroupWire[49]}}, {4{maskForGroupWire[48]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_lo_hi_3 = {{4{maskForGroupWire[51]}}, {4{maskForGroupWire[50]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_lo_3 = {fillBySeg_hi_hi_lo_lo_hi_3, fillBySeg_hi_hi_lo_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_lo_hi_lo_3 = {{4{maskForGroupWire[53]}}, {4{maskForGroupWire[52]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_hi_hi_3 = {{4{maskForGroupWire[55]}}, {4{maskForGroupWire[54]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_hi_3 = {fillBySeg_hi_hi_lo_hi_hi_3, fillBySeg_hi_hi_lo_hi_lo_3};
  wire [31:0]      fillBySeg_hi_hi_lo_3 = {fillBySeg_hi_hi_lo_hi_3, fillBySeg_hi_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_hi_lo_lo_3 = {{4{maskForGroupWire[57]}}, {4{maskForGroupWire[56]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_lo_hi_3 = {{4{maskForGroupWire[59]}}, {4{maskForGroupWire[58]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_lo_3 = {fillBySeg_hi_hi_hi_lo_hi_3, fillBySeg_hi_hi_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_hi_hi_lo_3 = {{4{maskForGroupWire[61]}}, {4{maskForGroupWire[60]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_hi_hi_3 = {{4{maskForGroupWire[63]}}, {4{maskForGroupWire[62]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_hi_lo_3};
  wire [31:0]      fillBySeg_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_lo_3};
  wire [63:0]      fillBySeg_hi_hi_3 = {fillBySeg_hi_hi_hi_3, fillBySeg_hi_hi_lo_3};
  wire [127:0]     fillBySeg_hi_3 = {fillBySeg_hi_hi_3, fillBySeg_hi_lo_3};
  wire [9:0]       fillBySeg_lo_lo_lo_lo_lo_4 = {{5{maskForGroupWire[1]}}, {5{maskForGroupWire[0]}}};
  wire [9:0]       fillBySeg_lo_lo_lo_lo_hi_4 = {{5{maskForGroupWire[3]}}, {5{maskForGroupWire[2]}}};
  wire [19:0]      fillBySeg_lo_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_lo_lo_hi_lo_4 = {{5{maskForGroupWire[5]}}, {5{maskForGroupWire[4]}}};
  wire [9:0]       fillBySeg_lo_lo_lo_hi_hi_4 = {{5{maskForGroupWire[7]}}, {5{maskForGroupWire[6]}}};
  wire [19:0]      fillBySeg_lo_lo_lo_hi_4 = {fillBySeg_lo_lo_lo_hi_hi_4, fillBySeg_lo_lo_lo_hi_lo_4};
  wire [39:0]      fillBySeg_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_lo_hi_lo_lo_4 = {{5{maskForGroupWire[9]}}, {5{maskForGroupWire[8]}}};
  wire [9:0]       fillBySeg_lo_lo_hi_lo_hi_4 = {{5{maskForGroupWire[11]}}, {5{maskForGroupWire[10]}}};
  wire [19:0]      fillBySeg_lo_lo_hi_lo_4 = {fillBySeg_lo_lo_hi_lo_hi_4, fillBySeg_lo_lo_hi_lo_lo_4};
  wire [9:0]       fillBySeg_lo_lo_hi_hi_lo_4 = {{5{maskForGroupWire[13]}}, {5{maskForGroupWire[12]}}};
  wire [9:0]       fillBySeg_lo_lo_hi_hi_hi_4 = {{5{maskForGroupWire[15]}}, {5{maskForGroupWire[14]}}};
  wire [19:0]      fillBySeg_lo_lo_hi_hi_4 = {fillBySeg_lo_lo_hi_hi_hi_4, fillBySeg_lo_lo_hi_hi_lo_4};
  wire [39:0]      fillBySeg_lo_lo_hi_4 = {fillBySeg_lo_lo_hi_hi_4, fillBySeg_lo_lo_hi_lo_4};
  wire [79:0]      fillBySeg_lo_lo_4 = {fillBySeg_lo_lo_hi_4, fillBySeg_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_lo_lo_lo_4 = {{5{maskForGroupWire[17]}}, {5{maskForGroupWire[16]}}};
  wire [9:0]       fillBySeg_lo_hi_lo_lo_hi_4 = {{5{maskForGroupWire[19]}}, {5{maskForGroupWire[18]}}};
  wire [19:0]      fillBySeg_lo_hi_lo_lo_4 = {fillBySeg_lo_hi_lo_lo_hi_4, fillBySeg_lo_hi_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_lo_hi_lo_4 = {{5{maskForGroupWire[21]}}, {5{maskForGroupWire[20]}}};
  wire [9:0]       fillBySeg_lo_hi_lo_hi_hi_4 = {{5{maskForGroupWire[23]}}, {5{maskForGroupWire[22]}}};
  wire [19:0]      fillBySeg_lo_hi_lo_hi_4 = {fillBySeg_lo_hi_lo_hi_hi_4, fillBySeg_lo_hi_lo_hi_lo_4};
  wire [39:0]      fillBySeg_lo_hi_lo_4 = {fillBySeg_lo_hi_lo_hi_4, fillBySeg_lo_hi_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_hi_lo_lo_4 = {{5{maskForGroupWire[25]}}, {5{maskForGroupWire[24]}}};
  wire [9:0]       fillBySeg_lo_hi_hi_lo_hi_4 = {{5{maskForGroupWire[27]}}, {5{maskForGroupWire[26]}}};
  wire [19:0]      fillBySeg_lo_hi_hi_lo_4 = {fillBySeg_lo_hi_hi_lo_hi_4, fillBySeg_lo_hi_hi_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_hi_hi_lo_4 = {{5{maskForGroupWire[29]}}, {5{maskForGroupWire[28]}}};
  wire [9:0]       fillBySeg_lo_hi_hi_hi_hi_4 = {{5{maskForGroupWire[31]}}, {5{maskForGroupWire[30]}}};
  wire [19:0]      fillBySeg_lo_hi_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_hi_4, fillBySeg_lo_hi_hi_hi_lo_4};
  wire [39:0]      fillBySeg_lo_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_4, fillBySeg_lo_hi_hi_lo_4};
  wire [79:0]      fillBySeg_lo_hi_4 = {fillBySeg_lo_hi_hi_4, fillBySeg_lo_hi_lo_4};
  wire [159:0]     fillBySeg_lo_4 = {fillBySeg_lo_hi_4, fillBySeg_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_lo_lo_lo_4 = {{5{maskForGroupWire[33]}}, {5{maskForGroupWire[32]}}};
  wire [9:0]       fillBySeg_hi_lo_lo_lo_hi_4 = {{5{maskForGroupWire[35]}}, {5{maskForGroupWire[34]}}};
  wire [19:0]      fillBySeg_hi_lo_lo_lo_4 = {fillBySeg_hi_lo_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_lo_hi_lo_4 = {{5{maskForGroupWire[37]}}, {5{maskForGroupWire[36]}}};
  wire [9:0]       fillBySeg_hi_lo_lo_hi_hi_4 = {{5{maskForGroupWire[39]}}, {5{maskForGroupWire[38]}}};
  wire [19:0]      fillBySeg_hi_lo_lo_hi_4 = {fillBySeg_hi_lo_lo_hi_hi_4, fillBySeg_hi_lo_lo_hi_lo_4};
  wire [39:0]      fillBySeg_hi_lo_lo_4 = {fillBySeg_hi_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_hi_lo_lo_4 = {{5{maskForGroupWire[41]}}, {5{maskForGroupWire[40]}}};
  wire [9:0]       fillBySeg_hi_lo_hi_lo_hi_4 = {{5{maskForGroupWire[43]}}, {5{maskForGroupWire[42]}}};
  wire [19:0]      fillBySeg_hi_lo_hi_lo_4 = {fillBySeg_hi_lo_hi_lo_hi_4, fillBySeg_hi_lo_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_hi_hi_lo_4 = {{5{maskForGroupWire[45]}}, {5{maskForGroupWire[44]}}};
  wire [9:0]       fillBySeg_hi_lo_hi_hi_hi_4 = {{5{maskForGroupWire[47]}}, {5{maskForGroupWire[46]}}};
  wire [19:0]      fillBySeg_hi_lo_hi_hi_4 = {fillBySeg_hi_lo_hi_hi_hi_4, fillBySeg_hi_lo_hi_hi_lo_4};
  wire [39:0]      fillBySeg_hi_lo_hi_4 = {fillBySeg_hi_lo_hi_hi_4, fillBySeg_hi_lo_hi_lo_4};
  wire [79:0]      fillBySeg_hi_lo_4 = {fillBySeg_hi_lo_hi_4, fillBySeg_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_lo_lo_lo_4 = {{5{maskForGroupWire[49]}}, {5{maskForGroupWire[48]}}};
  wire [9:0]       fillBySeg_hi_hi_lo_lo_hi_4 = {{5{maskForGroupWire[51]}}, {5{maskForGroupWire[50]}}};
  wire [19:0]      fillBySeg_hi_hi_lo_lo_4 = {fillBySeg_hi_hi_lo_lo_hi_4, fillBySeg_hi_hi_lo_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_lo_hi_lo_4 = {{5{maskForGroupWire[53]}}, {5{maskForGroupWire[52]}}};
  wire [9:0]       fillBySeg_hi_hi_lo_hi_hi_4 = {{5{maskForGroupWire[55]}}, {5{maskForGroupWire[54]}}};
  wire [19:0]      fillBySeg_hi_hi_lo_hi_4 = {fillBySeg_hi_hi_lo_hi_hi_4, fillBySeg_hi_hi_lo_hi_lo_4};
  wire [39:0]      fillBySeg_hi_hi_lo_4 = {fillBySeg_hi_hi_lo_hi_4, fillBySeg_hi_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_hi_lo_lo_4 = {{5{maskForGroupWire[57]}}, {5{maskForGroupWire[56]}}};
  wire [9:0]       fillBySeg_hi_hi_hi_lo_hi_4 = {{5{maskForGroupWire[59]}}, {5{maskForGroupWire[58]}}};
  wire [19:0]      fillBySeg_hi_hi_hi_lo_4 = {fillBySeg_hi_hi_hi_lo_hi_4, fillBySeg_hi_hi_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_hi_hi_lo_4 = {{5{maskForGroupWire[61]}}, {5{maskForGroupWire[60]}}};
  wire [9:0]       fillBySeg_hi_hi_hi_hi_hi_4 = {{5{maskForGroupWire[63]}}, {5{maskForGroupWire[62]}}};
  wire [19:0]      fillBySeg_hi_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_hi_lo_4};
  wire [39:0]      fillBySeg_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_lo_4};
  wire [79:0]      fillBySeg_hi_hi_4 = {fillBySeg_hi_hi_hi_4, fillBySeg_hi_hi_lo_4};
  wire [159:0]     fillBySeg_hi_4 = {fillBySeg_hi_hi_4, fillBySeg_hi_lo_4};
  wire [11:0]      fillBySeg_lo_lo_lo_lo_lo_5 = {{6{maskForGroupWire[1]}}, {6{maskForGroupWire[0]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_lo_hi_5 = {{6{maskForGroupWire[3]}}, {6{maskForGroupWire[2]}}};
  wire [23:0]      fillBySeg_lo_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_lo_lo_hi_lo_5 = {{6{maskForGroupWire[5]}}, {6{maskForGroupWire[4]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_hi_hi_5 = {{6{maskForGroupWire[7]}}, {6{maskForGroupWire[6]}}};
  wire [23:0]      fillBySeg_lo_lo_lo_hi_5 = {fillBySeg_lo_lo_lo_hi_hi_5, fillBySeg_lo_lo_lo_hi_lo_5};
  wire [47:0]      fillBySeg_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_lo_hi_lo_lo_5 = {{6{maskForGroupWire[9]}}, {6{maskForGroupWire[8]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_lo_hi_5 = {{6{maskForGroupWire[11]}}, {6{maskForGroupWire[10]}}};
  wire [23:0]      fillBySeg_lo_lo_hi_lo_5 = {fillBySeg_lo_lo_hi_lo_hi_5, fillBySeg_lo_lo_hi_lo_lo_5};
  wire [11:0]      fillBySeg_lo_lo_hi_hi_lo_5 = {{6{maskForGroupWire[13]}}, {6{maskForGroupWire[12]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_hi_hi_5 = {{6{maskForGroupWire[15]}}, {6{maskForGroupWire[14]}}};
  wire [23:0]      fillBySeg_lo_lo_hi_hi_5 = {fillBySeg_lo_lo_hi_hi_hi_5, fillBySeg_lo_lo_hi_hi_lo_5};
  wire [47:0]      fillBySeg_lo_lo_hi_5 = {fillBySeg_lo_lo_hi_hi_5, fillBySeg_lo_lo_hi_lo_5};
  wire [95:0]      fillBySeg_lo_lo_5 = {fillBySeg_lo_lo_hi_5, fillBySeg_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_lo_lo_lo_5 = {{6{maskForGroupWire[17]}}, {6{maskForGroupWire[16]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_lo_hi_5 = {{6{maskForGroupWire[19]}}, {6{maskForGroupWire[18]}}};
  wire [23:0]      fillBySeg_lo_hi_lo_lo_5 = {fillBySeg_lo_hi_lo_lo_hi_5, fillBySeg_lo_hi_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_lo_hi_lo_5 = {{6{maskForGroupWire[21]}}, {6{maskForGroupWire[20]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_hi_hi_5 = {{6{maskForGroupWire[23]}}, {6{maskForGroupWire[22]}}};
  wire [23:0]      fillBySeg_lo_hi_lo_hi_5 = {fillBySeg_lo_hi_lo_hi_hi_5, fillBySeg_lo_hi_lo_hi_lo_5};
  wire [47:0]      fillBySeg_lo_hi_lo_5 = {fillBySeg_lo_hi_lo_hi_5, fillBySeg_lo_hi_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_hi_lo_lo_5 = {{6{maskForGroupWire[25]}}, {6{maskForGroupWire[24]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_lo_hi_5 = {{6{maskForGroupWire[27]}}, {6{maskForGroupWire[26]}}};
  wire [23:0]      fillBySeg_lo_hi_hi_lo_5 = {fillBySeg_lo_hi_hi_lo_hi_5, fillBySeg_lo_hi_hi_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_hi_hi_lo_5 = {{6{maskForGroupWire[29]}}, {6{maskForGroupWire[28]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_hi_hi_5 = {{6{maskForGroupWire[31]}}, {6{maskForGroupWire[30]}}};
  wire [23:0]      fillBySeg_lo_hi_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_hi_5, fillBySeg_lo_hi_hi_hi_lo_5};
  wire [47:0]      fillBySeg_lo_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_5, fillBySeg_lo_hi_hi_lo_5};
  wire [95:0]      fillBySeg_lo_hi_5 = {fillBySeg_lo_hi_hi_5, fillBySeg_lo_hi_lo_5};
  wire [191:0]     fillBySeg_lo_5 = {fillBySeg_lo_hi_5, fillBySeg_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_lo_lo_lo_5 = {{6{maskForGroupWire[33]}}, {6{maskForGroupWire[32]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_lo_hi_5 = {{6{maskForGroupWire[35]}}, {6{maskForGroupWire[34]}}};
  wire [23:0]      fillBySeg_hi_lo_lo_lo_5 = {fillBySeg_hi_lo_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_lo_hi_lo_5 = {{6{maskForGroupWire[37]}}, {6{maskForGroupWire[36]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_hi_hi_5 = {{6{maskForGroupWire[39]}}, {6{maskForGroupWire[38]}}};
  wire [23:0]      fillBySeg_hi_lo_lo_hi_5 = {fillBySeg_hi_lo_lo_hi_hi_5, fillBySeg_hi_lo_lo_hi_lo_5};
  wire [47:0]      fillBySeg_hi_lo_lo_5 = {fillBySeg_hi_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_hi_lo_lo_5 = {{6{maskForGroupWire[41]}}, {6{maskForGroupWire[40]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_lo_hi_5 = {{6{maskForGroupWire[43]}}, {6{maskForGroupWire[42]}}};
  wire [23:0]      fillBySeg_hi_lo_hi_lo_5 = {fillBySeg_hi_lo_hi_lo_hi_5, fillBySeg_hi_lo_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_hi_hi_lo_5 = {{6{maskForGroupWire[45]}}, {6{maskForGroupWire[44]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_hi_hi_5 = {{6{maskForGroupWire[47]}}, {6{maskForGroupWire[46]}}};
  wire [23:0]      fillBySeg_hi_lo_hi_hi_5 = {fillBySeg_hi_lo_hi_hi_hi_5, fillBySeg_hi_lo_hi_hi_lo_5};
  wire [47:0]      fillBySeg_hi_lo_hi_5 = {fillBySeg_hi_lo_hi_hi_5, fillBySeg_hi_lo_hi_lo_5};
  wire [95:0]      fillBySeg_hi_lo_5 = {fillBySeg_hi_lo_hi_5, fillBySeg_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_lo_lo_lo_5 = {{6{maskForGroupWire[49]}}, {6{maskForGroupWire[48]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_lo_hi_5 = {{6{maskForGroupWire[51]}}, {6{maskForGroupWire[50]}}};
  wire [23:0]      fillBySeg_hi_hi_lo_lo_5 = {fillBySeg_hi_hi_lo_lo_hi_5, fillBySeg_hi_hi_lo_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_lo_hi_lo_5 = {{6{maskForGroupWire[53]}}, {6{maskForGroupWire[52]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_hi_hi_5 = {{6{maskForGroupWire[55]}}, {6{maskForGroupWire[54]}}};
  wire [23:0]      fillBySeg_hi_hi_lo_hi_5 = {fillBySeg_hi_hi_lo_hi_hi_5, fillBySeg_hi_hi_lo_hi_lo_5};
  wire [47:0]      fillBySeg_hi_hi_lo_5 = {fillBySeg_hi_hi_lo_hi_5, fillBySeg_hi_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_hi_lo_lo_5 = {{6{maskForGroupWire[57]}}, {6{maskForGroupWire[56]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_lo_hi_5 = {{6{maskForGroupWire[59]}}, {6{maskForGroupWire[58]}}};
  wire [23:0]      fillBySeg_hi_hi_hi_lo_5 = {fillBySeg_hi_hi_hi_lo_hi_5, fillBySeg_hi_hi_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_hi_hi_lo_5 = {{6{maskForGroupWire[61]}}, {6{maskForGroupWire[60]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_hi_hi_5 = {{6{maskForGroupWire[63]}}, {6{maskForGroupWire[62]}}};
  wire [23:0]      fillBySeg_hi_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_hi_lo_5};
  wire [47:0]      fillBySeg_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_lo_5};
  wire [95:0]      fillBySeg_hi_hi_5 = {fillBySeg_hi_hi_hi_5, fillBySeg_hi_hi_lo_5};
  wire [191:0]     fillBySeg_hi_5 = {fillBySeg_hi_hi_5, fillBySeg_hi_lo_5};
  wire [13:0]      fillBySeg_lo_lo_lo_lo_lo_6 = {{7{maskForGroupWire[1]}}, {7{maskForGroupWire[0]}}};
  wire [13:0]      fillBySeg_lo_lo_lo_lo_hi_6 = {{7{maskForGroupWire[3]}}, {7{maskForGroupWire[2]}}};
  wire [27:0]      fillBySeg_lo_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_lo_lo_hi_lo_6 = {{7{maskForGroupWire[5]}}, {7{maskForGroupWire[4]}}};
  wire [13:0]      fillBySeg_lo_lo_lo_hi_hi_6 = {{7{maskForGroupWire[7]}}, {7{maskForGroupWire[6]}}};
  wire [27:0]      fillBySeg_lo_lo_lo_hi_6 = {fillBySeg_lo_lo_lo_hi_hi_6, fillBySeg_lo_lo_lo_hi_lo_6};
  wire [55:0]      fillBySeg_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_lo_hi_lo_lo_6 = {{7{maskForGroupWire[9]}}, {7{maskForGroupWire[8]}}};
  wire [13:0]      fillBySeg_lo_lo_hi_lo_hi_6 = {{7{maskForGroupWire[11]}}, {7{maskForGroupWire[10]}}};
  wire [27:0]      fillBySeg_lo_lo_hi_lo_6 = {fillBySeg_lo_lo_hi_lo_hi_6, fillBySeg_lo_lo_hi_lo_lo_6};
  wire [13:0]      fillBySeg_lo_lo_hi_hi_lo_6 = {{7{maskForGroupWire[13]}}, {7{maskForGroupWire[12]}}};
  wire [13:0]      fillBySeg_lo_lo_hi_hi_hi_6 = {{7{maskForGroupWire[15]}}, {7{maskForGroupWire[14]}}};
  wire [27:0]      fillBySeg_lo_lo_hi_hi_6 = {fillBySeg_lo_lo_hi_hi_hi_6, fillBySeg_lo_lo_hi_hi_lo_6};
  wire [55:0]      fillBySeg_lo_lo_hi_6 = {fillBySeg_lo_lo_hi_hi_6, fillBySeg_lo_lo_hi_lo_6};
  wire [111:0]     fillBySeg_lo_lo_6 = {fillBySeg_lo_lo_hi_6, fillBySeg_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_lo_lo_lo_6 = {{7{maskForGroupWire[17]}}, {7{maskForGroupWire[16]}}};
  wire [13:0]      fillBySeg_lo_hi_lo_lo_hi_6 = {{7{maskForGroupWire[19]}}, {7{maskForGroupWire[18]}}};
  wire [27:0]      fillBySeg_lo_hi_lo_lo_6 = {fillBySeg_lo_hi_lo_lo_hi_6, fillBySeg_lo_hi_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_lo_hi_lo_6 = {{7{maskForGroupWire[21]}}, {7{maskForGroupWire[20]}}};
  wire [13:0]      fillBySeg_lo_hi_lo_hi_hi_6 = {{7{maskForGroupWire[23]}}, {7{maskForGroupWire[22]}}};
  wire [27:0]      fillBySeg_lo_hi_lo_hi_6 = {fillBySeg_lo_hi_lo_hi_hi_6, fillBySeg_lo_hi_lo_hi_lo_6};
  wire [55:0]      fillBySeg_lo_hi_lo_6 = {fillBySeg_lo_hi_lo_hi_6, fillBySeg_lo_hi_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_hi_lo_lo_6 = {{7{maskForGroupWire[25]}}, {7{maskForGroupWire[24]}}};
  wire [13:0]      fillBySeg_lo_hi_hi_lo_hi_6 = {{7{maskForGroupWire[27]}}, {7{maskForGroupWire[26]}}};
  wire [27:0]      fillBySeg_lo_hi_hi_lo_6 = {fillBySeg_lo_hi_hi_lo_hi_6, fillBySeg_lo_hi_hi_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_hi_hi_lo_6 = {{7{maskForGroupWire[29]}}, {7{maskForGroupWire[28]}}};
  wire [13:0]      fillBySeg_lo_hi_hi_hi_hi_6 = {{7{maskForGroupWire[31]}}, {7{maskForGroupWire[30]}}};
  wire [27:0]      fillBySeg_lo_hi_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_hi_6, fillBySeg_lo_hi_hi_hi_lo_6};
  wire [55:0]      fillBySeg_lo_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_6, fillBySeg_lo_hi_hi_lo_6};
  wire [111:0]     fillBySeg_lo_hi_6 = {fillBySeg_lo_hi_hi_6, fillBySeg_lo_hi_lo_6};
  wire [223:0]     fillBySeg_lo_6 = {fillBySeg_lo_hi_6, fillBySeg_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_lo_lo_lo_6 = {{7{maskForGroupWire[33]}}, {7{maskForGroupWire[32]}}};
  wire [13:0]      fillBySeg_hi_lo_lo_lo_hi_6 = {{7{maskForGroupWire[35]}}, {7{maskForGroupWire[34]}}};
  wire [27:0]      fillBySeg_hi_lo_lo_lo_6 = {fillBySeg_hi_lo_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_lo_hi_lo_6 = {{7{maskForGroupWire[37]}}, {7{maskForGroupWire[36]}}};
  wire [13:0]      fillBySeg_hi_lo_lo_hi_hi_6 = {{7{maskForGroupWire[39]}}, {7{maskForGroupWire[38]}}};
  wire [27:0]      fillBySeg_hi_lo_lo_hi_6 = {fillBySeg_hi_lo_lo_hi_hi_6, fillBySeg_hi_lo_lo_hi_lo_6};
  wire [55:0]      fillBySeg_hi_lo_lo_6 = {fillBySeg_hi_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_hi_lo_lo_6 = {{7{maskForGroupWire[41]}}, {7{maskForGroupWire[40]}}};
  wire [13:0]      fillBySeg_hi_lo_hi_lo_hi_6 = {{7{maskForGroupWire[43]}}, {7{maskForGroupWire[42]}}};
  wire [27:0]      fillBySeg_hi_lo_hi_lo_6 = {fillBySeg_hi_lo_hi_lo_hi_6, fillBySeg_hi_lo_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_hi_hi_lo_6 = {{7{maskForGroupWire[45]}}, {7{maskForGroupWire[44]}}};
  wire [13:0]      fillBySeg_hi_lo_hi_hi_hi_6 = {{7{maskForGroupWire[47]}}, {7{maskForGroupWire[46]}}};
  wire [27:0]      fillBySeg_hi_lo_hi_hi_6 = {fillBySeg_hi_lo_hi_hi_hi_6, fillBySeg_hi_lo_hi_hi_lo_6};
  wire [55:0]      fillBySeg_hi_lo_hi_6 = {fillBySeg_hi_lo_hi_hi_6, fillBySeg_hi_lo_hi_lo_6};
  wire [111:0]     fillBySeg_hi_lo_6 = {fillBySeg_hi_lo_hi_6, fillBySeg_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_lo_lo_lo_6 = {{7{maskForGroupWire[49]}}, {7{maskForGroupWire[48]}}};
  wire [13:0]      fillBySeg_hi_hi_lo_lo_hi_6 = {{7{maskForGroupWire[51]}}, {7{maskForGroupWire[50]}}};
  wire [27:0]      fillBySeg_hi_hi_lo_lo_6 = {fillBySeg_hi_hi_lo_lo_hi_6, fillBySeg_hi_hi_lo_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_lo_hi_lo_6 = {{7{maskForGroupWire[53]}}, {7{maskForGroupWire[52]}}};
  wire [13:0]      fillBySeg_hi_hi_lo_hi_hi_6 = {{7{maskForGroupWire[55]}}, {7{maskForGroupWire[54]}}};
  wire [27:0]      fillBySeg_hi_hi_lo_hi_6 = {fillBySeg_hi_hi_lo_hi_hi_6, fillBySeg_hi_hi_lo_hi_lo_6};
  wire [55:0]      fillBySeg_hi_hi_lo_6 = {fillBySeg_hi_hi_lo_hi_6, fillBySeg_hi_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_hi_lo_lo_6 = {{7{maskForGroupWire[57]}}, {7{maskForGroupWire[56]}}};
  wire [13:0]      fillBySeg_hi_hi_hi_lo_hi_6 = {{7{maskForGroupWire[59]}}, {7{maskForGroupWire[58]}}};
  wire [27:0]      fillBySeg_hi_hi_hi_lo_6 = {fillBySeg_hi_hi_hi_lo_hi_6, fillBySeg_hi_hi_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_hi_hi_lo_6 = {{7{maskForGroupWire[61]}}, {7{maskForGroupWire[60]}}};
  wire [13:0]      fillBySeg_hi_hi_hi_hi_hi_6 = {{7{maskForGroupWire[63]}}, {7{maskForGroupWire[62]}}};
  wire [27:0]      fillBySeg_hi_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_hi_lo_6};
  wire [55:0]      fillBySeg_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_lo_6};
  wire [111:0]     fillBySeg_hi_hi_6 = {fillBySeg_hi_hi_hi_6, fillBySeg_hi_hi_lo_6};
  wire [223:0]     fillBySeg_hi_6 = {fillBySeg_hi_hi_6, fillBySeg_hi_lo_6};
  wire [15:0]      fillBySeg_lo_lo_lo_lo_lo_7 = {{8{maskForGroupWire[1]}}, {8{maskForGroupWire[0]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_lo_hi_7 = {{8{maskForGroupWire[3]}}, {8{maskForGroupWire[2]}}};
  wire [31:0]      fillBySeg_lo_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_lo_lo_hi_lo_7 = {{8{maskForGroupWire[5]}}, {8{maskForGroupWire[4]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_hi_hi_7 = {{8{maskForGroupWire[7]}}, {8{maskForGroupWire[6]}}};
  wire [31:0]      fillBySeg_lo_lo_lo_hi_7 = {fillBySeg_lo_lo_lo_hi_hi_7, fillBySeg_lo_lo_lo_hi_lo_7};
  wire [63:0]      fillBySeg_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_lo_hi_lo_lo_7 = {{8{maskForGroupWire[9]}}, {8{maskForGroupWire[8]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_lo_hi_7 = {{8{maskForGroupWire[11]}}, {8{maskForGroupWire[10]}}};
  wire [31:0]      fillBySeg_lo_lo_hi_lo_7 = {fillBySeg_lo_lo_hi_lo_hi_7, fillBySeg_lo_lo_hi_lo_lo_7};
  wire [15:0]      fillBySeg_lo_lo_hi_hi_lo_7 = {{8{maskForGroupWire[13]}}, {8{maskForGroupWire[12]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_hi_hi_7 = {{8{maskForGroupWire[15]}}, {8{maskForGroupWire[14]}}};
  wire [31:0]      fillBySeg_lo_lo_hi_hi_7 = {fillBySeg_lo_lo_hi_hi_hi_7, fillBySeg_lo_lo_hi_hi_lo_7};
  wire [63:0]      fillBySeg_lo_lo_hi_7 = {fillBySeg_lo_lo_hi_hi_7, fillBySeg_lo_lo_hi_lo_7};
  wire [127:0]     fillBySeg_lo_lo_7 = {fillBySeg_lo_lo_hi_7, fillBySeg_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_lo_lo_lo_7 = {{8{maskForGroupWire[17]}}, {8{maskForGroupWire[16]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_lo_hi_7 = {{8{maskForGroupWire[19]}}, {8{maskForGroupWire[18]}}};
  wire [31:0]      fillBySeg_lo_hi_lo_lo_7 = {fillBySeg_lo_hi_lo_lo_hi_7, fillBySeg_lo_hi_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_lo_hi_lo_7 = {{8{maskForGroupWire[21]}}, {8{maskForGroupWire[20]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_hi_hi_7 = {{8{maskForGroupWire[23]}}, {8{maskForGroupWire[22]}}};
  wire [31:0]      fillBySeg_lo_hi_lo_hi_7 = {fillBySeg_lo_hi_lo_hi_hi_7, fillBySeg_lo_hi_lo_hi_lo_7};
  wire [63:0]      fillBySeg_lo_hi_lo_7 = {fillBySeg_lo_hi_lo_hi_7, fillBySeg_lo_hi_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_hi_lo_lo_7 = {{8{maskForGroupWire[25]}}, {8{maskForGroupWire[24]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_lo_hi_7 = {{8{maskForGroupWire[27]}}, {8{maskForGroupWire[26]}}};
  wire [31:0]      fillBySeg_lo_hi_hi_lo_7 = {fillBySeg_lo_hi_hi_lo_hi_7, fillBySeg_lo_hi_hi_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_hi_hi_lo_7 = {{8{maskForGroupWire[29]}}, {8{maskForGroupWire[28]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_hi_hi_7 = {{8{maskForGroupWire[31]}}, {8{maskForGroupWire[30]}}};
  wire [31:0]      fillBySeg_lo_hi_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_hi_7, fillBySeg_lo_hi_hi_hi_lo_7};
  wire [63:0]      fillBySeg_lo_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_7, fillBySeg_lo_hi_hi_lo_7};
  wire [127:0]     fillBySeg_lo_hi_7 = {fillBySeg_lo_hi_hi_7, fillBySeg_lo_hi_lo_7};
  wire [255:0]     fillBySeg_lo_7 = {fillBySeg_lo_hi_7, fillBySeg_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_lo_lo_lo_7 = {{8{maskForGroupWire[33]}}, {8{maskForGroupWire[32]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_lo_hi_7 = {{8{maskForGroupWire[35]}}, {8{maskForGroupWire[34]}}};
  wire [31:0]      fillBySeg_hi_lo_lo_lo_7 = {fillBySeg_hi_lo_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_lo_hi_lo_7 = {{8{maskForGroupWire[37]}}, {8{maskForGroupWire[36]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_hi_hi_7 = {{8{maskForGroupWire[39]}}, {8{maskForGroupWire[38]}}};
  wire [31:0]      fillBySeg_hi_lo_lo_hi_7 = {fillBySeg_hi_lo_lo_hi_hi_7, fillBySeg_hi_lo_lo_hi_lo_7};
  wire [63:0]      fillBySeg_hi_lo_lo_7 = {fillBySeg_hi_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_hi_lo_lo_7 = {{8{maskForGroupWire[41]}}, {8{maskForGroupWire[40]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_lo_hi_7 = {{8{maskForGroupWire[43]}}, {8{maskForGroupWire[42]}}};
  wire [31:0]      fillBySeg_hi_lo_hi_lo_7 = {fillBySeg_hi_lo_hi_lo_hi_7, fillBySeg_hi_lo_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_hi_hi_lo_7 = {{8{maskForGroupWire[45]}}, {8{maskForGroupWire[44]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_hi_hi_7 = {{8{maskForGroupWire[47]}}, {8{maskForGroupWire[46]}}};
  wire [31:0]      fillBySeg_hi_lo_hi_hi_7 = {fillBySeg_hi_lo_hi_hi_hi_7, fillBySeg_hi_lo_hi_hi_lo_7};
  wire [63:0]      fillBySeg_hi_lo_hi_7 = {fillBySeg_hi_lo_hi_hi_7, fillBySeg_hi_lo_hi_lo_7};
  wire [127:0]     fillBySeg_hi_lo_7 = {fillBySeg_hi_lo_hi_7, fillBySeg_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_lo_lo_lo_7 = {{8{maskForGroupWire[49]}}, {8{maskForGroupWire[48]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_lo_hi_7 = {{8{maskForGroupWire[51]}}, {8{maskForGroupWire[50]}}};
  wire [31:0]      fillBySeg_hi_hi_lo_lo_7 = {fillBySeg_hi_hi_lo_lo_hi_7, fillBySeg_hi_hi_lo_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_lo_hi_lo_7 = {{8{maskForGroupWire[53]}}, {8{maskForGroupWire[52]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_hi_hi_7 = {{8{maskForGroupWire[55]}}, {8{maskForGroupWire[54]}}};
  wire [31:0]      fillBySeg_hi_hi_lo_hi_7 = {fillBySeg_hi_hi_lo_hi_hi_7, fillBySeg_hi_hi_lo_hi_lo_7};
  wire [63:0]      fillBySeg_hi_hi_lo_7 = {fillBySeg_hi_hi_lo_hi_7, fillBySeg_hi_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_hi_lo_lo_7 = {{8{maskForGroupWire[57]}}, {8{maskForGroupWire[56]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_lo_hi_7 = {{8{maskForGroupWire[59]}}, {8{maskForGroupWire[58]}}};
  wire [31:0]      fillBySeg_hi_hi_hi_lo_7 = {fillBySeg_hi_hi_hi_lo_hi_7, fillBySeg_hi_hi_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_hi_hi_lo_7 = {{8{maskForGroupWire[61]}}, {8{maskForGroupWire[60]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_hi_hi_7 = {{8{maskForGroupWire[63]}}, {8{maskForGroupWire[62]}}};
  wire [31:0]      fillBySeg_hi_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_hi_lo_7};
  wire [63:0]      fillBySeg_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_lo_7};
  wire [127:0]     fillBySeg_hi_hi_7 = {fillBySeg_hi_hi_hi_7, fillBySeg_hi_hi_lo_7};
  wire [255:0]     fillBySeg_hi_7 = {fillBySeg_hi_hi_7, fillBySeg_hi_lo_7};
  wire [511:0]     fillBySeg =
    {64'h0,
     {64'h0,
      {64'h0,
       {64'h0,
        {64'h0, {64'h0, {64'h0, _fillBySeg_T[0] ? {fillBySeg_hi, fillBySeg_lo} : 64'h0} | (_fillBySeg_T[1] ? {fillBySeg_hi_1, fillBySeg_lo_1} : 128'h0)} | (_fillBySeg_T[2] ? {fillBySeg_hi_2, fillBySeg_lo_2} : 192'h0)}
          | (_fillBySeg_T[3] ? {fillBySeg_hi_3, fillBySeg_lo_3} : 256'h0)} | (_fillBySeg_T[4] ? {fillBySeg_hi_4, fillBySeg_lo_4} : 320'h0)} | (_fillBySeg_T[5] ? {fillBySeg_hi_5, fillBySeg_lo_5} : 384'h0)}
       | (_fillBySeg_T[6] ? {fillBySeg_hi_6, fillBySeg_lo_6} : 448'h0)} | (_fillBySeg_T[7] ? {fillBySeg_hi_7, fillBySeg_lo_7} : 512'h0);
  wire [7:0]       dataRegroupBySew_0_0 = bufferStageEnqueueData_0[7:0];
  wire [7:0]       dataRegroupBySew_0_1 = bufferStageEnqueueData_0[15:8];
  wire [7:0]       dataRegroupBySew_0_2 = bufferStageEnqueueData_0[23:16];
  wire [7:0]       dataRegroupBySew_0_3 = bufferStageEnqueueData_0[31:24];
  wire [7:0]       dataRegroupBySew_0_4 = bufferStageEnqueueData_0[39:32];
  wire [7:0]       dataRegroupBySew_0_5 = bufferStageEnqueueData_0[47:40];
  wire [7:0]       dataRegroupBySew_0_6 = bufferStageEnqueueData_0[55:48];
  wire [7:0]       dataRegroupBySew_0_7 = bufferStageEnqueueData_0[63:56];
  wire [7:0]       dataRegroupBySew_0_8 = bufferStageEnqueueData_0[71:64];
  wire [7:0]       dataRegroupBySew_0_9 = bufferStageEnqueueData_0[79:72];
  wire [7:0]       dataRegroupBySew_0_10 = bufferStageEnqueueData_0[87:80];
  wire [7:0]       dataRegroupBySew_0_11 = bufferStageEnqueueData_0[95:88];
  wire [7:0]       dataRegroupBySew_0_12 = bufferStageEnqueueData_0[103:96];
  wire [7:0]       dataRegroupBySew_0_13 = bufferStageEnqueueData_0[111:104];
  wire [7:0]       dataRegroupBySew_0_14 = bufferStageEnqueueData_0[119:112];
  wire [7:0]       dataRegroupBySew_0_15 = bufferStageEnqueueData_0[127:120];
  wire [7:0]       dataRegroupBySew_0_16 = bufferStageEnqueueData_0[135:128];
  wire [7:0]       dataRegroupBySew_0_17 = bufferStageEnqueueData_0[143:136];
  wire [7:0]       dataRegroupBySew_0_18 = bufferStageEnqueueData_0[151:144];
  wire [7:0]       dataRegroupBySew_0_19 = bufferStageEnqueueData_0[159:152];
  wire [7:0]       dataRegroupBySew_0_20 = bufferStageEnqueueData_0[167:160];
  wire [7:0]       dataRegroupBySew_0_21 = bufferStageEnqueueData_0[175:168];
  wire [7:0]       dataRegroupBySew_0_22 = bufferStageEnqueueData_0[183:176];
  wire [7:0]       dataRegroupBySew_0_23 = bufferStageEnqueueData_0[191:184];
  wire [7:0]       dataRegroupBySew_0_24 = bufferStageEnqueueData_0[199:192];
  wire [7:0]       dataRegroupBySew_0_25 = bufferStageEnqueueData_0[207:200];
  wire [7:0]       dataRegroupBySew_0_26 = bufferStageEnqueueData_0[215:208];
  wire [7:0]       dataRegroupBySew_0_27 = bufferStageEnqueueData_0[223:216];
  wire [7:0]       dataRegroupBySew_0_28 = bufferStageEnqueueData_0[231:224];
  wire [7:0]       dataRegroupBySew_0_29 = bufferStageEnqueueData_0[239:232];
  wire [7:0]       dataRegroupBySew_0_30 = bufferStageEnqueueData_0[247:240];
  wire [7:0]       dataRegroupBySew_0_31 = bufferStageEnqueueData_0[255:248];
  wire [7:0]       dataRegroupBySew_0_32 = bufferStageEnqueueData_0[263:256];
  wire [7:0]       dataRegroupBySew_0_33 = bufferStageEnqueueData_0[271:264];
  wire [7:0]       dataRegroupBySew_0_34 = bufferStageEnqueueData_0[279:272];
  wire [7:0]       dataRegroupBySew_0_35 = bufferStageEnqueueData_0[287:280];
  wire [7:0]       dataRegroupBySew_0_36 = bufferStageEnqueueData_0[295:288];
  wire [7:0]       dataRegroupBySew_0_37 = bufferStageEnqueueData_0[303:296];
  wire [7:0]       dataRegroupBySew_0_38 = bufferStageEnqueueData_0[311:304];
  wire [7:0]       dataRegroupBySew_0_39 = bufferStageEnqueueData_0[319:312];
  wire [7:0]       dataRegroupBySew_0_40 = bufferStageEnqueueData_0[327:320];
  wire [7:0]       dataRegroupBySew_0_41 = bufferStageEnqueueData_0[335:328];
  wire [7:0]       dataRegroupBySew_0_42 = bufferStageEnqueueData_0[343:336];
  wire [7:0]       dataRegroupBySew_0_43 = bufferStageEnqueueData_0[351:344];
  wire [7:0]       dataRegroupBySew_0_44 = bufferStageEnqueueData_0[359:352];
  wire [7:0]       dataRegroupBySew_0_45 = bufferStageEnqueueData_0[367:360];
  wire [7:0]       dataRegroupBySew_0_46 = bufferStageEnqueueData_0[375:368];
  wire [7:0]       dataRegroupBySew_0_47 = bufferStageEnqueueData_0[383:376];
  wire [7:0]       dataRegroupBySew_0_48 = bufferStageEnqueueData_0[391:384];
  wire [7:0]       dataRegroupBySew_0_49 = bufferStageEnqueueData_0[399:392];
  wire [7:0]       dataRegroupBySew_0_50 = bufferStageEnqueueData_0[407:400];
  wire [7:0]       dataRegroupBySew_0_51 = bufferStageEnqueueData_0[415:408];
  wire [7:0]       dataRegroupBySew_0_52 = bufferStageEnqueueData_0[423:416];
  wire [7:0]       dataRegroupBySew_0_53 = bufferStageEnqueueData_0[431:424];
  wire [7:0]       dataRegroupBySew_0_54 = bufferStageEnqueueData_0[439:432];
  wire [7:0]       dataRegroupBySew_0_55 = bufferStageEnqueueData_0[447:440];
  wire [7:0]       dataRegroupBySew_0_56 = bufferStageEnqueueData_0[455:448];
  wire [7:0]       dataRegroupBySew_0_57 = bufferStageEnqueueData_0[463:456];
  wire [7:0]       dataRegroupBySew_0_58 = bufferStageEnqueueData_0[471:464];
  wire [7:0]       dataRegroupBySew_0_59 = bufferStageEnqueueData_0[479:472];
  wire [7:0]       dataRegroupBySew_0_60 = bufferStageEnqueueData_0[487:480];
  wire [7:0]       dataRegroupBySew_0_61 = bufferStageEnqueueData_0[495:488];
  wire [7:0]       dataRegroupBySew_0_62 = bufferStageEnqueueData_0[503:496];
  wire [7:0]       dataRegroupBySew_0_63 = bufferStageEnqueueData_0[511:504];
  wire [7:0]       dataRegroupBySew_1_0 = bufferStageEnqueueData_1[7:0];
  wire [7:0]       dataRegroupBySew_1_1 = bufferStageEnqueueData_1[15:8];
  wire [7:0]       dataRegroupBySew_1_2 = bufferStageEnqueueData_1[23:16];
  wire [7:0]       dataRegroupBySew_1_3 = bufferStageEnqueueData_1[31:24];
  wire [7:0]       dataRegroupBySew_1_4 = bufferStageEnqueueData_1[39:32];
  wire [7:0]       dataRegroupBySew_1_5 = bufferStageEnqueueData_1[47:40];
  wire [7:0]       dataRegroupBySew_1_6 = bufferStageEnqueueData_1[55:48];
  wire [7:0]       dataRegroupBySew_1_7 = bufferStageEnqueueData_1[63:56];
  wire [7:0]       dataRegroupBySew_1_8 = bufferStageEnqueueData_1[71:64];
  wire [7:0]       dataRegroupBySew_1_9 = bufferStageEnqueueData_1[79:72];
  wire [7:0]       dataRegroupBySew_1_10 = bufferStageEnqueueData_1[87:80];
  wire [7:0]       dataRegroupBySew_1_11 = bufferStageEnqueueData_1[95:88];
  wire [7:0]       dataRegroupBySew_1_12 = bufferStageEnqueueData_1[103:96];
  wire [7:0]       dataRegroupBySew_1_13 = bufferStageEnqueueData_1[111:104];
  wire [7:0]       dataRegroupBySew_1_14 = bufferStageEnqueueData_1[119:112];
  wire [7:0]       dataRegroupBySew_1_15 = bufferStageEnqueueData_1[127:120];
  wire [7:0]       dataRegroupBySew_1_16 = bufferStageEnqueueData_1[135:128];
  wire [7:0]       dataRegroupBySew_1_17 = bufferStageEnqueueData_1[143:136];
  wire [7:0]       dataRegroupBySew_1_18 = bufferStageEnqueueData_1[151:144];
  wire [7:0]       dataRegroupBySew_1_19 = bufferStageEnqueueData_1[159:152];
  wire [7:0]       dataRegroupBySew_1_20 = bufferStageEnqueueData_1[167:160];
  wire [7:0]       dataRegroupBySew_1_21 = bufferStageEnqueueData_1[175:168];
  wire [7:0]       dataRegroupBySew_1_22 = bufferStageEnqueueData_1[183:176];
  wire [7:0]       dataRegroupBySew_1_23 = bufferStageEnqueueData_1[191:184];
  wire [7:0]       dataRegroupBySew_1_24 = bufferStageEnqueueData_1[199:192];
  wire [7:0]       dataRegroupBySew_1_25 = bufferStageEnqueueData_1[207:200];
  wire [7:0]       dataRegroupBySew_1_26 = bufferStageEnqueueData_1[215:208];
  wire [7:0]       dataRegroupBySew_1_27 = bufferStageEnqueueData_1[223:216];
  wire [7:0]       dataRegroupBySew_1_28 = bufferStageEnqueueData_1[231:224];
  wire [7:0]       dataRegroupBySew_1_29 = bufferStageEnqueueData_1[239:232];
  wire [7:0]       dataRegroupBySew_1_30 = bufferStageEnqueueData_1[247:240];
  wire [7:0]       dataRegroupBySew_1_31 = bufferStageEnqueueData_1[255:248];
  wire [7:0]       dataRegroupBySew_1_32 = bufferStageEnqueueData_1[263:256];
  wire [7:0]       dataRegroupBySew_1_33 = bufferStageEnqueueData_1[271:264];
  wire [7:0]       dataRegroupBySew_1_34 = bufferStageEnqueueData_1[279:272];
  wire [7:0]       dataRegroupBySew_1_35 = bufferStageEnqueueData_1[287:280];
  wire [7:0]       dataRegroupBySew_1_36 = bufferStageEnqueueData_1[295:288];
  wire [7:0]       dataRegroupBySew_1_37 = bufferStageEnqueueData_1[303:296];
  wire [7:0]       dataRegroupBySew_1_38 = bufferStageEnqueueData_1[311:304];
  wire [7:0]       dataRegroupBySew_1_39 = bufferStageEnqueueData_1[319:312];
  wire [7:0]       dataRegroupBySew_1_40 = bufferStageEnqueueData_1[327:320];
  wire [7:0]       dataRegroupBySew_1_41 = bufferStageEnqueueData_1[335:328];
  wire [7:0]       dataRegroupBySew_1_42 = bufferStageEnqueueData_1[343:336];
  wire [7:0]       dataRegroupBySew_1_43 = bufferStageEnqueueData_1[351:344];
  wire [7:0]       dataRegroupBySew_1_44 = bufferStageEnqueueData_1[359:352];
  wire [7:0]       dataRegroupBySew_1_45 = bufferStageEnqueueData_1[367:360];
  wire [7:0]       dataRegroupBySew_1_46 = bufferStageEnqueueData_1[375:368];
  wire [7:0]       dataRegroupBySew_1_47 = bufferStageEnqueueData_1[383:376];
  wire [7:0]       dataRegroupBySew_1_48 = bufferStageEnqueueData_1[391:384];
  wire [7:0]       dataRegroupBySew_1_49 = bufferStageEnqueueData_1[399:392];
  wire [7:0]       dataRegroupBySew_1_50 = bufferStageEnqueueData_1[407:400];
  wire [7:0]       dataRegroupBySew_1_51 = bufferStageEnqueueData_1[415:408];
  wire [7:0]       dataRegroupBySew_1_52 = bufferStageEnqueueData_1[423:416];
  wire [7:0]       dataRegroupBySew_1_53 = bufferStageEnqueueData_1[431:424];
  wire [7:0]       dataRegroupBySew_1_54 = bufferStageEnqueueData_1[439:432];
  wire [7:0]       dataRegroupBySew_1_55 = bufferStageEnqueueData_1[447:440];
  wire [7:0]       dataRegroupBySew_1_56 = bufferStageEnqueueData_1[455:448];
  wire [7:0]       dataRegroupBySew_1_57 = bufferStageEnqueueData_1[463:456];
  wire [7:0]       dataRegroupBySew_1_58 = bufferStageEnqueueData_1[471:464];
  wire [7:0]       dataRegroupBySew_1_59 = bufferStageEnqueueData_1[479:472];
  wire [7:0]       dataRegroupBySew_1_60 = bufferStageEnqueueData_1[487:480];
  wire [7:0]       dataRegroupBySew_1_61 = bufferStageEnqueueData_1[495:488];
  wire [7:0]       dataRegroupBySew_1_62 = bufferStageEnqueueData_1[503:496];
  wire [7:0]       dataRegroupBySew_1_63 = bufferStageEnqueueData_1[511:504];
  wire [7:0]       dataRegroupBySew_2_0 = bufferStageEnqueueData_2[7:0];
  wire [7:0]       dataRegroupBySew_2_1 = bufferStageEnqueueData_2[15:8];
  wire [7:0]       dataRegroupBySew_2_2 = bufferStageEnqueueData_2[23:16];
  wire [7:0]       dataRegroupBySew_2_3 = bufferStageEnqueueData_2[31:24];
  wire [7:0]       dataRegroupBySew_2_4 = bufferStageEnqueueData_2[39:32];
  wire [7:0]       dataRegroupBySew_2_5 = bufferStageEnqueueData_2[47:40];
  wire [7:0]       dataRegroupBySew_2_6 = bufferStageEnqueueData_2[55:48];
  wire [7:0]       dataRegroupBySew_2_7 = bufferStageEnqueueData_2[63:56];
  wire [7:0]       dataRegroupBySew_2_8 = bufferStageEnqueueData_2[71:64];
  wire [7:0]       dataRegroupBySew_2_9 = bufferStageEnqueueData_2[79:72];
  wire [7:0]       dataRegroupBySew_2_10 = bufferStageEnqueueData_2[87:80];
  wire [7:0]       dataRegroupBySew_2_11 = bufferStageEnqueueData_2[95:88];
  wire [7:0]       dataRegroupBySew_2_12 = bufferStageEnqueueData_2[103:96];
  wire [7:0]       dataRegroupBySew_2_13 = bufferStageEnqueueData_2[111:104];
  wire [7:0]       dataRegroupBySew_2_14 = bufferStageEnqueueData_2[119:112];
  wire [7:0]       dataRegroupBySew_2_15 = bufferStageEnqueueData_2[127:120];
  wire [7:0]       dataRegroupBySew_2_16 = bufferStageEnqueueData_2[135:128];
  wire [7:0]       dataRegroupBySew_2_17 = bufferStageEnqueueData_2[143:136];
  wire [7:0]       dataRegroupBySew_2_18 = bufferStageEnqueueData_2[151:144];
  wire [7:0]       dataRegroupBySew_2_19 = bufferStageEnqueueData_2[159:152];
  wire [7:0]       dataRegroupBySew_2_20 = bufferStageEnqueueData_2[167:160];
  wire [7:0]       dataRegroupBySew_2_21 = bufferStageEnqueueData_2[175:168];
  wire [7:0]       dataRegroupBySew_2_22 = bufferStageEnqueueData_2[183:176];
  wire [7:0]       dataRegroupBySew_2_23 = bufferStageEnqueueData_2[191:184];
  wire [7:0]       dataRegroupBySew_2_24 = bufferStageEnqueueData_2[199:192];
  wire [7:0]       dataRegroupBySew_2_25 = bufferStageEnqueueData_2[207:200];
  wire [7:0]       dataRegroupBySew_2_26 = bufferStageEnqueueData_2[215:208];
  wire [7:0]       dataRegroupBySew_2_27 = bufferStageEnqueueData_2[223:216];
  wire [7:0]       dataRegroupBySew_2_28 = bufferStageEnqueueData_2[231:224];
  wire [7:0]       dataRegroupBySew_2_29 = bufferStageEnqueueData_2[239:232];
  wire [7:0]       dataRegroupBySew_2_30 = bufferStageEnqueueData_2[247:240];
  wire [7:0]       dataRegroupBySew_2_31 = bufferStageEnqueueData_2[255:248];
  wire [7:0]       dataRegroupBySew_2_32 = bufferStageEnqueueData_2[263:256];
  wire [7:0]       dataRegroupBySew_2_33 = bufferStageEnqueueData_2[271:264];
  wire [7:0]       dataRegroupBySew_2_34 = bufferStageEnqueueData_2[279:272];
  wire [7:0]       dataRegroupBySew_2_35 = bufferStageEnqueueData_2[287:280];
  wire [7:0]       dataRegroupBySew_2_36 = bufferStageEnqueueData_2[295:288];
  wire [7:0]       dataRegroupBySew_2_37 = bufferStageEnqueueData_2[303:296];
  wire [7:0]       dataRegroupBySew_2_38 = bufferStageEnqueueData_2[311:304];
  wire [7:0]       dataRegroupBySew_2_39 = bufferStageEnqueueData_2[319:312];
  wire [7:0]       dataRegroupBySew_2_40 = bufferStageEnqueueData_2[327:320];
  wire [7:0]       dataRegroupBySew_2_41 = bufferStageEnqueueData_2[335:328];
  wire [7:0]       dataRegroupBySew_2_42 = bufferStageEnqueueData_2[343:336];
  wire [7:0]       dataRegroupBySew_2_43 = bufferStageEnqueueData_2[351:344];
  wire [7:0]       dataRegroupBySew_2_44 = bufferStageEnqueueData_2[359:352];
  wire [7:0]       dataRegroupBySew_2_45 = bufferStageEnqueueData_2[367:360];
  wire [7:0]       dataRegroupBySew_2_46 = bufferStageEnqueueData_2[375:368];
  wire [7:0]       dataRegroupBySew_2_47 = bufferStageEnqueueData_2[383:376];
  wire [7:0]       dataRegroupBySew_2_48 = bufferStageEnqueueData_2[391:384];
  wire [7:0]       dataRegroupBySew_2_49 = bufferStageEnqueueData_2[399:392];
  wire [7:0]       dataRegroupBySew_2_50 = bufferStageEnqueueData_2[407:400];
  wire [7:0]       dataRegroupBySew_2_51 = bufferStageEnqueueData_2[415:408];
  wire [7:0]       dataRegroupBySew_2_52 = bufferStageEnqueueData_2[423:416];
  wire [7:0]       dataRegroupBySew_2_53 = bufferStageEnqueueData_2[431:424];
  wire [7:0]       dataRegroupBySew_2_54 = bufferStageEnqueueData_2[439:432];
  wire [7:0]       dataRegroupBySew_2_55 = bufferStageEnqueueData_2[447:440];
  wire [7:0]       dataRegroupBySew_2_56 = bufferStageEnqueueData_2[455:448];
  wire [7:0]       dataRegroupBySew_2_57 = bufferStageEnqueueData_2[463:456];
  wire [7:0]       dataRegroupBySew_2_58 = bufferStageEnqueueData_2[471:464];
  wire [7:0]       dataRegroupBySew_2_59 = bufferStageEnqueueData_2[479:472];
  wire [7:0]       dataRegroupBySew_2_60 = bufferStageEnqueueData_2[487:480];
  wire [7:0]       dataRegroupBySew_2_61 = bufferStageEnqueueData_2[495:488];
  wire [7:0]       dataRegroupBySew_2_62 = bufferStageEnqueueData_2[503:496];
  wire [7:0]       dataRegroupBySew_2_63 = bufferStageEnqueueData_2[511:504];
  wire [7:0]       dataRegroupBySew_3_0 = bufferStageEnqueueData_3[7:0];
  wire [7:0]       dataRegroupBySew_3_1 = bufferStageEnqueueData_3[15:8];
  wire [7:0]       dataRegroupBySew_3_2 = bufferStageEnqueueData_3[23:16];
  wire [7:0]       dataRegroupBySew_3_3 = bufferStageEnqueueData_3[31:24];
  wire [7:0]       dataRegroupBySew_3_4 = bufferStageEnqueueData_3[39:32];
  wire [7:0]       dataRegroupBySew_3_5 = bufferStageEnqueueData_3[47:40];
  wire [7:0]       dataRegroupBySew_3_6 = bufferStageEnqueueData_3[55:48];
  wire [7:0]       dataRegroupBySew_3_7 = bufferStageEnqueueData_3[63:56];
  wire [7:0]       dataRegroupBySew_3_8 = bufferStageEnqueueData_3[71:64];
  wire [7:0]       dataRegroupBySew_3_9 = bufferStageEnqueueData_3[79:72];
  wire [7:0]       dataRegroupBySew_3_10 = bufferStageEnqueueData_3[87:80];
  wire [7:0]       dataRegroupBySew_3_11 = bufferStageEnqueueData_3[95:88];
  wire [7:0]       dataRegroupBySew_3_12 = bufferStageEnqueueData_3[103:96];
  wire [7:0]       dataRegroupBySew_3_13 = bufferStageEnqueueData_3[111:104];
  wire [7:0]       dataRegroupBySew_3_14 = bufferStageEnqueueData_3[119:112];
  wire [7:0]       dataRegroupBySew_3_15 = bufferStageEnqueueData_3[127:120];
  wire [7:0]       dataRegroupBySew_3_16 = bufferStageEnqueueData_3[135:128];
  wire [7:0]       dataRegroupBySew_3_17 = bufferStageEnqueueData_3[143:136];
  wire [7:0]       dataRegroupBySew_3_18 = bufferStageEnqueueData_3[151:144];
  wire [7:0]       dataRegroupBySew_3_19 = bufferStageEnqueueData_3[159:152];
  wire [7:0]       dataRegroupBySew_3_20 = bufferStageEnqueueData_3[167:160];
  wire [7:0]       dataRegroupBySew_3_21 = bufferStageEnqueueData_3[175:168];
  wire [7:0]       dataRegroupBySew_3_22 = bufferStageEnqueueData_3[183:176];
  wire [7:0]       dataRegroupBySew_3_23 = bufferStageEnqueueData_3[191:184];
  wire [7:0]       dataRegroupBySew_3_24 = bufferStageEnqueueData_3[199:192];
  wire [7:0]       dataRegroupBySew_3_25 = bufferStageEnqueueData_3[207:200];
  wire [7:0]       dataRegroupBySew_3_26 = bufferStageEnqueueData_3[215:208];
  wire [7:0]       dataRegroupBySew_3_27 = bufferStageEnqueueData_3[223:216];
  wire [7:0]       dataRegroupBySew_3_28 = bufferStageEnqueueData_3[231:224];
  wire [7:0]       dataRegroupBySew_3_29 = bufferStageEnqueueData_3[239:232];
  wire [7:0]       dataRegroupBySew_3_30 = bufferStageEnqueueData_3[247:240];
  wire [7:0]       dataRegroupBySew_3_31 = bufferStageEnqueueData_3[255:248];
  wire [7:0]       dataRegroupBySew_3_32 = bufferStageEnqueueData_3[263:256];
  wire [7:0]       dataRegroupBySew_3_33 = bufferStageEnqueueData_3[271:264];
  wire [7:0]       dataRegroupBySew_3_34 = bufferStageEnqueueData_3[279:272];
  wire [7:0]       dataRegroupBySew_3_35 = bufferStageEnqueueData_3[287:280];
  wire [7:0]       dataRegroupBySew_3_36 = bufferStageEnqueueData_3[295:288];
  wire [7:0]       dataRegroupBySew_3_37 = bufferStageEnqueueData_3[303:296];
  wire [7:0]       dataRegroupBySew_3_38 = bufferStageEnqueueData_3[311:304];
  wire [7:0]       dataRegroupBySew_3_39 = bufferStageEnqueueData_3[319:312];
  wire [7:0]       dataRegroupBySew_3_40 = bufferStageEnqueueData_3[327:320];
  wire [7:0]       dataRegroupBySew_3_41 = bufferStageEnqueueData_3[335:328];
  wire [7:0]       dataRegroupBySew_3_42 = bufferStageEnqueueData_3[343:336];
  wire [7:0]       dataRegroupBySew_3_43 = bufferStageEnqueueData_3[351:344];
  wire [7:0]       dataRegroupBySew_3_44 = bufferStageEnqueueData_3[359:352];
  wire [7:0]       dataRegroupBySew_3_45 = bufferStageEnqueueData_3[367:360];
  wire [7:0]       dataRegroupBySew_3_46 = bufferStageEnqueueData_3[375:368];
  wire [7:0]       dataRegroupBySew_3_47 = bufferStageEnqueueData_3[383:376];
  wire [7:0]       dataRegroupBySew_3_48 = bufferStageEnqueueData_3[391:384];
  wire [7:0]       dataRegroupBySew_3_49 = bufferStageEnqueueData_3[399:392];
  wire [7:0]       dataRegroupBySew_3_50 = bufferStageEnqueueData_3[407:400];
  wire [7:0]       dataRegroupBySew_3_51 = bufferStageEnqueueData_3[415:408];
  wire [7:0]       dataRegroupBySew_3_52 = bufferStageEnqueueData_3[423:416];
  wire [7:0]       dataRegroupBySew_3_53 = bufferStageEnqueueData_3[431:424];
  wire [7:0]       dataRegroupBySew_3_54 = bufferStageEnqueueData_3[439:432];
  wire [7:0]       dataRegroupBySew_3_55 = bufferStageEnqueueData_3[447:440];
  wire [7:0]       dataRegroupBySew_3_56 = bufferStageEnqueueData_3[455:448];
  wire [7:0]       dataRegroupBySew_3_57 = bufferStageEnqueueData_3[463:456];
  wire [7:0]       dataRegroupBySew_3_58 = bufferStageEnqueueData_3[471:464];
  wire [7:0]       dataRegroupBySew_3_59 = bufferStageEnqueueData_3[479:472];
  wire [7:0]       dataRegroupBySew_3_60 = bufferStageEnqueueData_3[487:480];
  wire [7:0]       dataRegroupBySew_3_61 = bufferStageEnqueueData_3[495:488];
  wire [7:0]       dataRegroupBySew_3_62 = bufferStageEnqueueData_3[503:496];
  wire [7:0]       dataRegroupBySew_3_63 = bufferStageEnqueueData_3[511:504];
  wire [7:0]       dataRegroupBySew_4_0 = bufferStageEnqueueData_4[7:0];
  wire [7:0]       dataRegroupBySew_4_1 = bufferStageEnqueueData_4[15:8];
  wire [7:0]       dataRegroupBySew_4_2 = bufferStageEnqueueData_4[23:16];
  wire [7:0]       dataRegroupBySew_4_3 = bufferStageEnqueueData_4[31:24];
  wire [7:0]       dataRegroupBySew_4_4 = bufferStageEnqueueData_4[39:32];
  wire [7:0]       dataRegroupBySew_4_5 = bufferStageEnqueueData_4[47:40];
  wire [7:0]       dataRegroupBySew_4_6 = bufferStageEnqueueData_4[55:48];
  wire [7:0]       dataRegroupBySew_4_7 = bufferStageEnqueueData_4[63:56];
  wire [7:0]       dataRegroupBySew_4_8 = bufferStageEnqueueData_4[71:64];
  wire [7:0]       dataRegroupBySew_4_9 = bufferStageEnqueueData_4[79:72];
  wire [7:0]       dataRegroupBySew_4_10 = bufferStageEnqueueData_4[87:80];
  wire [7:0]       dataRegroupBySew_4_11 = bufferStageEnqueueData_4[95:88];
  wire [7:0]       dataRegroupBySew_4_12 = bufferStageEnqueueData_4[103:96];
  wire [7:0]       dataRegroupBySew_4_13 = bufferStageEnqueueData_4[111:104];
  wire [7:0]       dataRegroupBySew_4_14 = bufferStageEnqueueData_4[119:112];
  wire [7:0]       dataRegroupBySew_4_15 = bufferStageEnqueueData_4[127:120];
  wire [7:0]       dataRegroupBySew_4_16 = bufferStageEnqueueData_4[135:128];
  wire [7:0]       dataRegroupBySew_4_17 = bufferStageEnqueueData_4[143:136];
  wire [7:0]       dataRegroupBySew_4_18 = bufferStageEnqueueData_4[151:144];
  wire [7:0]       dataRegroupBySew_4_19 = bufferStageEnqueueData_4[159:152];
  wire [7:0]       dataRegroupBySew_4_20 = bufferStageEnqueueData_4[167:160];
  wire [7:0]       dataRegroupBySew_4_21 = bufferStageEnqueueData_4[175:168];
  wire [7:0]       dataRegroupBySew_4_22 = bufferStageEnqueueData_4[183:176];
  wire [7:0]       dataRegroupBySew_4_23 = bufferStageEnqueueData_4[191:184];
  wire [7:0]       dataRegroupBySew_4_24 = bufferStageEnqueueData_4[199:192];
  wire [7:0]       dataRegroupBySew_4_25 = bufferStageEnqueueData_4[207:200];
  wire [7:0]       dataRegroupBySew_4_26 = bufferStageEnqueueData_4[215:208];
  wire [7:0]       dataRegroupBySew_4_27 = bufferStageEnqueueData_4[223:216];
  wire [7:0]       dataRegroupBySew_4_28 = bufferStageEnqueueData_4[231:224];
  wire [7:0]       dataRegroupBySew_4_29 = bufferStageEnqueueData_4[239:232];
  wire [7:0]       dataRegroupBySew_4_30 = bufferStageEnqueueData_4[247:240];
  wire [7:0]       dataRegroupBySew_4_31 = bufferStageEnqueueData_4[255:248];
  wire [7:0]       dataRegroupBySew_4_32 = bufferStageEnqueueData_4[263:256];
  wire [7:0]       dataRegroupBySew_4_33 = bufferStageEnqueueData_4[271:264];
  wire [7:0]       dataRegroupBySew_4_34 = bufferStageEnqueueData_4[279:272];
  wire [7:0]       dataRegroupBySew_4_35 = bufferStageEnqueueData_4[287:280];
  wire [7:0]       dataRegroupBySew_4_36 = bufferStageEnqueueData_4[295:288];
  wire [7:0]       dataRegroupBySew_4_37 = bufferStageEnqueueData_4[303:296];
  wire [7:0]       dataRegroupBySew_4_38 = bufferStageEnqueueData_4[311:304];
  wire [7:0]       dataRegroupBySew_4_39 = bufferStageEnqueueData_4[319:312];
  wire [7:0]       dataRegroupBySew_4_40 = bufferStageEnqueueData_4[327:320];
  wire [7:0]       dataRegroupBySew_4_41 = bufferStageEnqueueData_4[335:328];
  wire [7:0]       dataRegroupBySew_4_42 = bufferStageEnqueueData_4[343:336];
  wire [7:0]       dataRegroupBySew_4_43 = bufferStageEnqueueData_4[351:344];
  wire [7:0]       dataRegroupBySew_4_44 = bufferStageEnqueueData_4[359:352];
  wire [7:0]       dataRegroupBySew_4_45 = bufferStageEnqueueData_4[367:360];
  wire [7:0]       dataRegroupBySew_4_46 = bufferStageEnqueueData_4[375:368];
  wire [7:0]       dataRegroupBySew_4_47 = bufferStageEnqueueData_4[383:376];
  wire [7:0]       dataRegroupBySew_4_48 = bufferStageEnqueueData_4[391:384];
  wire [7:0]       dataRegroupBySew_4_49 = bufferStageEnqueueData_4[399:392];
  wire [7:0]       dataRegroupBySew_4_50 = bufferStageEnqueueData_4[407:400];
  wire [7:0]       dataRegroupBySew_4_51 = bufferStageEnqueueData_4[415:408];
  wire [7:0]       dataRegroupBySew_4_52 = bufferStageEnqueueData_4[423:416];
  wire [7:0]       dataRegroupBySew_4_53 = bufferStageEnqueueData_4[431:424];
  wire [7:0]       dataRegroupBySew_4_54 = bufferStageEnqueueData_4[439:432];
  wire [7:0]       dataRegroupBySew_4_55 = bufferStageEnqueueData_4[447:440];
  wire [7:0]       dataRegroupBySew_4_56 = bufferStageEnqueueData_4[455:448];
  wire [7:0]       dataRegroupBySew_4_57 = bufferStageEnqueueData_4[463:456];
  wire [7:0]       dataRegroupBySew_4_58 = bufferStageEnqueueData_4[471:464];
  wire [7:0]       dataRegroupBySew_4_59 = bufferStageEnqueueData_4[479:472];
  wire [7:0]       dataRegroupBySew_4_60 = bufferStageEnqueueData_4[487:480];
  wire [7:0]       dataRegroupBySew_4_61 = bufferStageEnqueueData_4[495:488];
  wire [7:0]       dataRegroupBySew_4_62 = bufferStageEnqueueData_4[503:496];
  wire [7:0]       dataRegroupBySew_4_63 = bufferStageEnqueueData_4[511:504];
  wire [7:0]       dataRegroupBySew_5_0 = bufferStageEnqueueData_5[7:0];
  wire [7:0]       dataRegroupBySew_5_1 = bufferStageEnqueueData_5[15:8];
  wire [7:0]       dataRegroupBySew_5_2 = bufferStageEnqueueData_5[23:16];
  wire [7:0]       dataRegroupBySew_5_3 = bufferStageEnqueueData_5[31:24];
  wire [7:0]       dataRegroupBySew_5_4 = bufferStageEnqueueData_5[39:32];
  wire [7:0]       dataRegroupBySew_5_5 = bufferStageEnqueueData_5[47:40];
  wire [7:0]       dataRegroupBySew_5_6 = bufferStageEnqueueData_5[55:48];
  wire [7:0]       dataRegroupBySew_5_7 = bufferStageEnqueueData_5[63:56];
  wire [7:0]       dataRegroupBySew_5_8 = bufferStageEnqueueData_5[71:64];
  wire [7:0]       dataRegroupBySew_5_9 = bufferStageEnqueueData_5[79:72];
  wire [7:0]       dataRegroupBySew_5_10 = bufferStageEnqueueData_5[87:80];
  wire [7:0]       dataRegroupBySew_5_11 = bufferStageEnqueueData_5[95:88];
  wire [7:0]       dataRegroupBySew_5_12 = bufferStageEnqueueData_5[103:96];
  wire [7:0]       dataRegroupBySew_5_13 = bufferStageEnqueueData_5[111:104];
  wire [7:0]       dataRegroupBySew_5_14 = bufferStageEnqueueData_5[119:112];
  wire [7:0]       dataRegroupBySew_5_15 = bufferStageEnqueueData_5[127:120];
  wire [7:0]       dataRegroupBySew_5_16 = bufferStageEnqueueData_5[135:128];
  wire [7:0]       dataRegroupBySew_5_17 = bufferStageEnqueueData_5[143:136];
  wire [7:0]       dataRegroupBySew_5_18 = bufferStageEnqueueData_5[151:144];
  wire [7:0]       dataRegroupBySew_5_19 = bufferStageEnqueueData_5[159:152];
  wire [7:0]       dataRegroupBySew_5_20 = bufferStageEnqueueData_5[167:160];
  wire [7:0]       dataRegroupBySew_5_21 = bufferStageEnqueueData_5[175:168];
  wire [7:0]       dataRegroupBySew_5_22 = bufferStageEnqueueData_5[183:176];
  wire [7:0]       dataRegroupBySew_5_23 = bufferStageEnqueueData_5[191:184];
  wire [7:0]       dataRegroupBySew_5_24 = bufferStageEnqueueData_5[199:192];
  wire [7:0]       dataRegroupBySew_5_25 = bufferStageEnqueueData_5[207:200];
  wire [7:0]       dataRegroupBySew_5_26 = bufferStageEnqueueData_5[215:208];
  wire [7:0]       dataRegroupBySew_5_27 = bufferStageEnqueueData_5[223:216];
  wire [7:0]       dataRegroupBySew_5_28 = bufferStageEnqueueData_5[231:224];
  wire [7:0]       dataRegroupBySew_5_29 = bufferStageEnqueueData_5[239:232];
  wire [7:0]       dataRegroupBySew_5_30 = bufferStageEnqueueData_5[247:240];
  wire [7:0]       dataRegroupBySew_5_31 = bufferStageEnqueueData_5[255:248];
  wire [7:0]       dataRegroupBySew_5_32 = bufferStageEnqueueData_5[263:256];
  wire [7:0]       dataRegroupBySew_5_33 = bufferStageEnqueueData_5[271:264];
  wire [7:0]       dataRegroupBySew_5_34 = bufferStageEnqueueData_5[279:272];
  wire [7:0]       dataRegroupBySew_5_35 = bufferStageEnqueueData_5[287:280];
  wire [7:0]       dataRegroupBySew_5_36 = bufferStageEnqueueData_5[295:288];
  wire [7:0]       dataRegroupBySew_5_37 = bufferStageEnqueueData_5[303:296];
  wire [7:0]       dataRegroupBySew_5_38 = bufferStageEnqueueData_5[311:304];
  wire [7:0]       dataRegroupBySew_5_39 = bufferStageEnqueueData_5[319:312];
  wire [7:0]       dataRegroupBySew_5_40 = bufferStageEnqueueData_5[327:320];
  wire [7:0]       dataRegroupBySew_5_41 = bufferStageEnqueueData_5[335:328];
  wire [7:0]       dataRegroupBySew_5_42 = bufferStageEnqueueData_5[343:336];
  wire [7:0]       dataRegroupBySew_5_43 = bufferStageEnqueueData_5[351:344];
  wire [7:0]       dataRegroupBySew_5_44 = bufferStageEnqueueData_5[359:352];
  wire [7:0]       dataRegroupBySew_5_45 = bufferStageEnqueueData_5[367:360];
  wire [7:0]       dataRegroupBySew_5_46 = bufferStageEnqueueData_5[375:368];
  wire [7:0]       dataRegroupBySew_5_47 = bufferStageEnqueueData_5[383:376];
  wire [7:0]       dataRegroupBySew_5_48 = bufferStageEnqueueData_5[391:384];
  wire [7:0]       dataRegroupBySew_5_49 = bufferStageEnqueueData_5[399:392];
  wire [7:0]       dataRegroupBySew_5_50 = bufferStageEnqueueData_5[407:400];
  wire [7:0]       dataRegroupBySew_5_51 = bufferStageEnqueueData_5[415:408];
  wire [7:0]       dataRegroupBySew_5_52 = bufferStageEnqueueData_5[423:416];
  wire [7:0]       dataRegroupBySew_5_53 = bufferStageEnqueueData_5[431:424];
  wire [7:0]       dataRegroupBySew_5_54 = bufferStageEnqueueData_5[439:432];
  wire [7:0]       dataRegroupBySew_5_55 = bufferStageEnqueueData_5[447:440];
  wire [7:0]       dataRegroupBySew_5_56 = bufferStageEnqueueData_5[455:448];
  wire [7:0]       dataRegroupBySew_5_57 = bufferStageEnqueueData_5[463:456];
  wire [7:0]       dataRegroupBySew_5_58 = bufferStageEnqueueData_5[471:464];
  wire [7:0]       dataRegroupBySew_5_59 = bufferStageEnqueueData_5[479:472];
  wire [7:0]       dataRegroupBySew_5_60 = bufferStageEnqueueData_5[487:480];
  wire [7:0]       dataRegroupBySew_5_61 = bufferStageEnqueueData_5[495:488];
  wire [7:0]       dataRegroupBySew_5_62 = bufferStageEnqueueData_5[503:496];
  wire [7:0]       dataRegroupBySew_5_63 = bufferStageEnqueueData_5[511:504];
  wire [7:0]       dataRegroupBySew_6_0 = bufferStageEnqueueData_6[7:0];
  wire [7:0]       dataRegroupBySew_6_1 = bufferStageEnqueueData_6[15:8];
  wire [7:0]       dataRegroupBySew_6_2 = bufferStageEnqueueData_6[23:16];
  wire [7:0]       dataRegroupBySew_6_3 = bufferStageEnqueueData_6[31:24];
  wire [7:0]       dataRegroupBySew_6_4 = bufferStageEnqueueData_6[39:32];
  wire [7:0]       dataRegroupBySew_6_5 = bufferStageEnqueueData_6[47:40];
  wire [7:0]       dataRegroupBySew_6_6 = bufferStageEnqueueData_6[55:48];
  wire [7:0]       dataRegroupBySew_6_7 = bufferStageEnqueueData_6[63:56];
  wire [7:0]       dataRegroupBySew_6_8 = bufferStageEnqueueData_6[71:64];
  wire [7:0]       dataRegroupBySew_6_9 = bufferStageEnqueueData_6[79:72];
  wire [7:0]       dataRegroupBySew_6_10 = bufferStageEnqueueData_6[87:80];
  wire [7:0]       dataRegroupBySew_6_11 = bufferStageEnqueueData_6[95:88];
  wire [7:0]       dataRegroupBySew_6_12 = bufferStageEnqueueData_6[103:96];
  wire [7:0]       dataRegroupBySew_6_13 = bufferStageEnqueueData_6[111:104];
  wire [7:0]       dataRegroupBySew_6_14 = bufferStageEnqueueData_6[119:112];
  wire [7:0]       dataRegroupBySew_6_15 = bufferStageEnqueueData_6[127:120];
  wire [7:0]       dataRegroupBySew_6_16 = bufferStageEnqueueData_6[135:128];
  wire [7:0]       dataRegroupBySew_6_17 = bufferStageEnqueueData_6[143:136];
  wire [7:0]       dataRegroupBySew_6_18 = bufferStageEnqueueData_6[151:144];
  wire [7:0]       dataRegroupBySew_6_19 = bufferStageEnqueueData_6[159:152];
  wire [7:0]       dataRegroupBySew_6_20 = bufferStageEnqueueData_6[167:160];
  wire [7:0]       dataRegroupBySew_6_21 = bufferStageEnqueueData_6[175:168];
  wire [7:0]       dataRegroupBySew_6_22 = bufferStageEnqueueData_6[183:176];
  wire [7:0]       dataRegroupBySew_6_23 = bufferStageEnqueueData_6[191:184];
  wire [7:0]       dataRegroupBySew_6_24 = bufferStageEnqueueData_6[199:192];
  wire [7:0]       dataRegroupBySew_6_25 = bufferStageEnqueueData_6[207:200];
  wire [7:0]       dataRegroupBySew_6_26 = bufferStageEnqueueData_6[215:208];
  wire [7:0]       dataRegroupBySew_6_27 = bufferStageEnqueueData_6[223:216];
  wire [7:0]       dataRegroupBySew_6_28 = bufferStageEnqueueData_6[231:224];
  wire [7:0]       dataRegroupBySew_6_29 = bufferStageEnqueueData_6[239:232];
  wire [7:0]       dataRegroupBySew_6_30 = bufferStageEnqueueData_6[247:240];
  wire [7:0]       dataRegroupBySew_6_31 = bufferStageEnqueueData_6[255:248];
  wire [7:0]       dataRegroupBySew_6_32 = bufferStageEnqueueData_6[263:256];
  wire [7:0]       dataRegroupBySew_6_33 = bufferStageEnqueueData_6[271:264];
  wire [7:0]       dataRegroupBySew_6_34 = bufferStageEnqueueData_6[279:272];
  wire [7:0]       dataRegroupBySew_6_35 = bufferStageEnqueueData_6[287:280];
  wire [7:0]       dataRegroupBySew_6_36 = bufferStageEnqueueData_6[295:288];
  wire [7:0]       dataRegroupBySew_6_37 = bufferStageEnqueueData_6[303:296];
  wire [7:0]       dataRegroupBySew_6_38 = bufferStageEnqueueData_6[311:304];
  wire [7:0]       dataRegroupBySew_6_39 = bufferStageEnqueueData_6[319:312];
  wire [7:0]       dataRegroupBySew_6_40 = bufferStageEnqueueData_6[327:320];
  wire [7:0]       dataRegroupBySew_6_41 = bufferStageEnqueueData_6[335:328];
  wire [7:0]       dataRegroupBySew_6_42 = bufferStageEnqueueData_6[343:336];
  wire [7:0]       dataRegroupBySew_6_43 = bufferStageEnqueueData_6[351:344];
  wire [7:0]       dataRegroupBySew_6_44 = bufferStageEnqueueData_6[359:352];
  wire [7:0]       dataRegroupBySew_6_45 = bufferStageEnqueueData_6[367:360];
  wire [7:0]       dataRegroupBySew_6_46 = bufferStageEnqueueData_6[375:368];
  wire [7:0]       dataRegroupBySew_6_47 = bufferStageEnqueueData_6[383:376];
  wire [7:0]       dataRegroupBySew_6_48 = bufferStageEnqueueData_6[391:384];
  wire [7:0]       dataRegroupBySew_6_49 = bufferStageEnqueueData_6[399:392];
  wire [7:0]       dataRegroupBySew_6_50 = bufferStageEnqueueData_6[407:400];
  wire [7:0]       dataRegroupBySew_6_51 = bufferStageEnqueueData_6[415:408];
  wire [7:0]       dataRegroupBySew_6_52 = bufferStageEnqueueData_6[423:416];
  wire [7:0]       dataRegroupBySew_6_53 = bufferStageEnqueueData_6[431:424];
  wire [7:0]       dataRegroupBySew_6_54 = bufferStageEnqueueData_6[439:432];
  wire [7:0]       dataRegroupBySew_6_55 = bufferStageEnqueueData_6[447:440];
  wire [7:0]       dataRegroupBySew_6_56 = bufferStageEnqueueData_6[455:448];
  wire [7:0]       dataRegroupBySew_6_57 = bufferStageEnqueueData_6[463:456];
  wire [7:0]       dataRegroupBySew_6_58 = bufferStageEnqueueData_6[471:464];
  wire [7:0]       dataRegroupBySew_6_59 = bufferStageEnqueueData_6[479:472];
  wire [7:0]       dataRegroupBySew_6_60 = bufferStageEnqueueData_6[487:480];
  wire [7:0]       dataRegroupBySew_6_61 = bufferStageEnqueueData_6[495:488];
  wire [7:0]       dataRegroupBySew_6_62 = bufferStageEnqueueData_6[503:496];
  wire [7:0]       dataRegroupBySew_6_63 = bufferStageEnqueueData_6[511:504];
  wire [7:0]       dataRegroupBySew_7_0 = bufferStageEnqueueData_7[7:0];
  wire [7:0]       dataRegroupBySew_7_1 = bufferStageEnqueueData_7[15:8];
  wire [7:0]       dataRegroupBySew_7_2 = bufferStageEnqueueData_7[23:16];
  wire [7:0]       dataRegroupBySew_7_3 = bufferStageEnqueueData_7[31:24];
  wire [7:0]       dataRegroupBySew_7_4 = bufferStageEnqueueData_7[39:32];
  wire [7:0]       dataRegroupBySew_7_5 = bufferStageEnqueueData_7[47:40];
  wire [7:0]       dataRegroupBySew_7_6 = bufferStageEnqueueData_7[55:48];
  wire [7:0]       dataRegroupBySew_7_7 = bufferStageEnqueueData_7[63:56];
  wire [7:0]       dataRegroupBySew_7_8 = bufferStageEnqueueData_7[71:64];
  wire [7:0]       dataRegroupBySew_7_9 = bufferStageEnqueueData_7[79:72];
  wire [7:0]       dataRegroupBySew_7_10 = bufferStageEnqueueData_7[87:80];
  wire [7:0]       dataRegroupBySew_7_11 = bufferStageEnqueueData_7[95:88];
  wire [7:0]       dataRegroupBySew_7_12 = bufferStageEnqueueData_7[103:96];
  wire [7:0]       dataRegroupBySew_7_13 = bufferStageEnqueueData_7[111:104];
  wire [7:0]       dataRegroupBySew_7_14 = bufferStageEnqueueData_7[119:112];
  wire [7:0]       dataRegroupBySew_7_15 = bufferStageEnqueueData_7[127:120];
  wire [7:0]       dataRegroupBySew_7_16 = bufferStageEnqueueData_7[135:128];
  wire [7:0]       dataRegroupBySew_7_17 = bufferStageEnqueueData_7[143:136];
  wire [7:0]       dataRegroupBySew_7_18 = bufferStageEnqueueData_7[151:144];
  wire [7:0]       dataRegroupBySew_7_19 = bufferStageEnqueueData_7[159:152];
  wire [7:0]       dataRegroupBySew_7_20 = bufferStageEnqueueData_7[167:160];
  wire [7:0]       dataRegroupBySew_7_21 = bufferStageEnqueueData_7[175:168];
  wire [7:0]       dataRegroupBySew_7_22 = bufferStageEnqueueData_7[183:176];
  wire [7:0]       dataRegroupBySew_7_23 = bufferStageEnqueueData_7[191:184];
  wire [7:0]       dataRegroupBySew_7_24 = bufferStageEnqueueData_7[199:192];
  wire [7:0]       dataRegroupBySew_7_25 = bufferStageEnqueueData_7[207:200];
  wire [7:0]       dataRegroupBySew_7_26 = bufferStageEnqueueData_7[215:208];
  wire [7:0]       dataRegroupBySew_7_27 = bufferStageEnqueueData_7[223:216];
  wire [7:0]       dataRegroupBySew_7_28 = bufferStageEnqueueData_7[231:224];
  wire [7:0]       dataRegroupBySew_7_29 = bufferStageEnqueueData_7[239:232];
  wire [7:0]       dataRegroupBySew_7_30 = bufferStageEnqueueData_7[247:240];
  wire [7:0]       dataRegroupBySew_7_31 = bufferStageEnqueueData_7[255:248];
  wire [7:0]       dataRegroupBySew_7_32 = bufferStageEnqueueData_7[263:256];
  wire [7:0]       dataRegroupBySew_7_33 = bufferStageEnqueueData_7[271:264];
  wire [7:0]       dataRegroupBySew_7_34 = bufferStageEnqueueData_7[279:272];
  wire [7:0]       dataRegroupBySew_7_35 = bufferStageEnqueueData_7[287:280];
  wire [7:0]       dataRegroupBySew_7_36 = bufferStageEnqueueData_7[295:288];
  wire [7:0]       dataRegroupBySew_7_37 = bufferStageEnqueueData_7[303:296];
  wire [7:0]       dataRegroupBySew_7_38 = bufferStageEnqueueData_7[311:304];
  wire [7:0]       dataRegroupBySew_7_39 = bufferStageEnqueueData_7[319:312];
  wire [7:0]       dataRegroupBySew_7_40 = bufferStageEnqueueData_7[327:320];
  wire [7:0]       dataRegroupBySew_7_41 = bufferStageEnqueueData_7[335:328];
  wire [7:0]       dataRegroupBySew_7_42 = bufferStageEnqueueData_7[343:336];
  wire [7:0]       dataRegroupBySew_7_43 = bufferStageEnqueueData_7[351:344];
  wire [7:0]       dataRegroupBySew_7_44 = bufferStageEnqueueData_7[359:352];
  wire [7:0]       dataRegroupBySew_7_45 = bufferStageEnqueueData_7[367:360];
  wire [7:0]       dataRegroupBySew_7_46 = bufferStageEnqueueData_7[375:368];
  wire [7:0]       dataRegroupBySew_7_47 = bufferStageEnqueueData_7[383:376];
  wire [7:0]       dataRegroupBySew_7_48 = bufferStageEnqueueData_7[391:384];
  wire [7:0]       dataRegroupBySew_7_49 = bufferStageEnqueueData_7[399:392];
  wire [7:0]       dataRegroupBySew_7_50 = bufferStageEnqueueData_7[407:400];
  wire [7:0]       dataRegroupBySew_7_51 = bufferStageEnqueueData_7[415:408];
  wire [7:0]       dataRegroupBySew_7_52 = bufferStageEnqueueData_7[423:416];
  wire [7:0]       dataRegroupBySew_7_53 = bufferStageEnqueueData_7[431:424];
  wire [7:0]       dataRegroupBySew_7_54 = bufferStageEnqueueData_7[439:432];
  wire [7:0]       dataRegroupBySew_7_55 = bufferStageEnqueueData_7[447:440];
  wire [7:0]       dataRegroupBySew_7_56 = bufferStageEnqueueData_7[455:448];
  wire [7:0]       dataRegroupBySew_7_57 = bufferStageEnqueueData_7[463:456];
  wire [7:0]       dataRegroupBySew_7_58 = bufferStageEnqueueData_7[471:464];
  wire [7:0]       dataRegroupBySew_7_59 = bufferStageEnqueueData_7[479:472];
  wire [7:0]       dataRegroupBySew_7_60 = bufferStageEnqueueData_7[487:480];
  wire [7:0]       dataRegroupBySew_7_61 = bufferStageEnqueueData_7[495:488];
  wire [7:0]       dataRegroupBySew_7_62 = bufferStageEnqueueData_7[503:496];
  wire [7:0]       dataRegroupBySew_7_63 = bufferStageEnqueueData_7[511:504];
  wire [15:0]      dataInMem_lo_lo_lo_lo_lo = {dataRegroupBySew_0_1, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_lo_lo_lo_hi = {dataRegroupBySew_0_3, dataRegroupBySew_0_2};
  wire [31:0]      dataInMem_lo_lo_lo_lo = {dataInMem_lo_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo_lo};
  wire [15:0]      dataInMem_lo_lo_lo_hi_lo = {dataRegroupBySew_0_5, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_lo_lo_hi_hi = {dataRegroupBySew_0_7, dataRegroupBySew_0_6};
  wire [31:0]      dataInMem_lo_lo_lo_hi = {dataInMem_lo_lo_lo_hi_hi, dataInMem_lo_lo_lo_hi_lo};
  wire [63:0]      dataInMem_lo_lo_lo = {dataInMem_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo};
  wire [15:0]      dataInMem_lo_lo_hi_lo_lo = {dataRegroupBySew_0_9, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_lo_lo_hi_lo_hi = {dataRegroupBySew_0_11, dataRegroupBySew_0_10};
  wire [31:0]      dataInMem_lo_lo_hi_lo = {dataInMem_lo_lo_hi_lo_hi, dataInMem_lo_lo_hi_lo_lo};
  wire [15:0]      dataInMem_lo_lo_hi_hi_lo = {dataRegroupBySew_0_13, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_lo_lo_hi_hi_hi = {dataRegroupBySew_0_15, dataRegroupBySew_0_14};
  wire [31:0]      dataInMem_lo_lo_hi_hi = {dataInMem_lo_lo_hi_hi_hi, dataInMem_lo_lo_hi_hi_lo};
  wire [63:0]      dataInMem_lo_lo_hi = {dataInMem_lo_lo_hi_hi, dataInMem_lo_lo_hi_lo};
  wire [127:0]     dataInMem_lo_lo = {dataInMem_lo_lo_hi, dataInMem_lo_lo_lo};
  wire [15:0]      dataInMem_lo_hi_lo_lo_lo = {dataRegroupBySew_0_17, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_lo_hi_lo_lo_hi = {dataRegroupBySew_0_19, dataRegroupBySew_0_18};
  wire [31:0]      dataInMem_lo_hi_lo_lo = {dataInMem_lo_hi_lo_lo_hi, dataInMem_lo_hi_lo_lo_lo};
  wire [15:0]      dataInMem_lo_hi_lo_hi_lo = {dataRegroupBySew_0_21, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_lo_hi_lo_hi_hi = {dataRegroupBySew_0_23, dataRegroupBySew_0_22};
  wire [31:0]      dataInMem_lo_hi_lo_hi = {dataInMem_lo_hi_lo_hi_hi, dataInMem_lo_hi_lo_hi_lo};
  wire [63:0]      dataInMem_lo_hi_lo = {dataInMem_lo_hi_lo_hi, dataInMem_lo_hi_lo_lo};
  wire [15:0]      dataInMem_lo_hi_hi_lo_lo = {dataRegroupBySew_0_25, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_lo_hi_hi_lo_hi = {dataRegroupBySew_0_27, dataRegroupBySew_0_26};
  wire [31:0]      dataInMem_lo_hi_hi_lo = {dataInMem_lo_hi_hi_lo_hi, dataInMem_lo_hi_hi_lo_lo};
  wire [15:0]      dataInMem_lo_hi_hi_hi_lo = {dataRegroupBySew_0_29, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_lo_hi_hi_hi_hi = {dataRegroupBySew_0_31, dataRegroupBySew_0_30};
  wire [31:0]      dataInMem_lo_hi_hi_hi = {dataInMem_lo_hi_hi_hi_hi, dataInMem_lo_hi_hi_hi_lo};
  wire [63:0]      dataInMem_lo_hi_hi = {dataInMem_lo_hi_hi_hi, dataInMem_lo_hi_hi_lo};
  wire [127:0]     dataInMem_lo_hi = {dataInMem_lo_hi_hi, dataInMem_lo_hi_lo};
  wire [255:0]     dataInMem_lo = {dataInMem_lo_hi, dataInMem_lo_lo};
  wire [15:0]      dataInMem_hi_lo_lo_lo_lo = {dataRegroupBySew_0_33, dataRegroupBySew_0_32};
  wire [15:0]      dataInMem_hi_lo_lo_lo_hi = {dataRegroupBySew_0_35, dataRegroupBySew_0_34};
  wire [31:0]      dataInMem_hi_lo_lo_lo = {dataInMem_hi_lo_lo_lo_hi, dataInMem_hi_lo_lo_lo_lo};
  wire [15:0]      dataInMem_hi_lo_lo_hi_lo = {dataRegroupBySew_0_37, dataRegroupBySew_0_36};
  wire [15:0]      dataInMem_hi_lo_lo_hi_hi = {dataRegroupBySew_0_39, dataRegroupBySew_0_38};
  wire [31:0]      dataInMem_hi_lo_lo_hi = {dataInMem_hi_lo_lo_hi_hi, dataInMem_hi_lo_lo_hi_lo};
  wire [63:0]      dataInMem_hi_lo_lo = {dataInMem_hi_lo_lo_hi, dataInMem_hi_lo_lo_lo};
  wire [15:0]      dataInMem_hi_lo_hi_lo_lo = {dataRegroupBySew_0_41, dataRegroupBySew_0_40};
  wire [15:0]      dataInMem_hi_lo_hi_lo_hi = {dataRegroupBySew_0_43, dataRegroupBySew_0_42};
  wire [31:0]      dataInMem_hi_lo_hi_lo = {dataInMem_hi_lo_hi_lo_hi, dataInMem_hi_lo_hi_lo_lo};
  wire [15:0]      dataInMem_hi_lo_hi_hi_lo = {dataRegroupBySew_0_45, dataRegroupBySew_0_44};
  wire [15:0]      dataInMem_hi_lo_hi_hi_hi = {dataRegroupBySew_0_47, dataRegroupBySew_0_46};
  wire [31:0]      dataInMem_hi_lo_hi_hi = {dataInMem_hi_lo_hi_hi_hi, dataInMem_hi_lo_hi_hi_lo};
  wire [63:0]      dataInMem_hi_lo_hi = {dataInMem_hi_lo_hi_hi, dataInMem_hi_lo_hi_lo};
  wire [127:0]     dataInMem_hi_lo = {dataInMem_hi_lo_hi, dataInMem_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_lo_lo_lo = {dataRegroupBySew_0_49, dataRegroupBySew_0_48};
  wire [15:0]      dataInMem_hi_hi_lo_lo_hi = {dataRegroupBySew_0_51, dataRegroupBySew_0_50};
  wire [31:0]      dataInMem_hi_hi_lo_lo = {dataInMem_hi_hi_lo_lo_hi, dataInMem_hi_hi_lo_lo_lo};
  wire [15:0]      dataInMem_hi_hi_lo_hi_lo = {dataRegroupBySew_0_53, dataRegroupBySew_0_52};
  wire [15:0]      dataInMem_hi_hi_lo_hi_hi = {dataRegroupBySew_0_55, dataRegroupBySew_0_54};
  wire [31:0]      dataInMem_hi_hi_lo_hi = {dataInMem_hi_hi_lo_hi_hi, dataInMem_hi_hi_lo_hi_lo};
  wire [63:0]      dataInMem_hi_hi_lo = {dataInMem_hi_hi_lo_hi, dataInMem_hi_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_hi_lo_lo = {dataRegroupBySew_0_57, dataRegroupBySew_0_56};
  wire [15:0]      dataInMem_hi_hi_hi_lo_hi = {dataRegroupBySew_0_59, dataRegroupBySew_0_58};
  wire [31:0]      dataInMem_hi_hi_hi_lo = {dataInMem_hi_hi_hi_lo_hi, dataInMem_hi_hi_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_hi_hi_lo = {dataRegroupBySew_0_61, dataRegroupBySew_0_60};
  wire [15:0]      dataInMem_hi_hi_hi_hi_hi = {dataRegroupBySew_0_63, dataRegroupBySew_0_62};
  wire [31:0]      dataInMem_hi_hi_hi_hi = {dataInMem_hi_hi_hi_hi_hi, dataInMem_hi_hi_hi_hi_lo};
  wire [63:0]      dataInMem_hi_hi_hi = {dataInMem_hi_hi_hi_hi, dataInMem_hi_hi_hi_lo};
  wire [127:0]     dataInMem_hi_hi = {dataInMem_hi_hi_hi, dataInMem_hi_hi_lo};
  wire [255:0]     dataInMem_hi = {dataInMem_hi_hi, dataInMem_hi_lo};
  wire [511:0]     dataInMem = {dataInMem_hi, dataInMem_lo};
  wire [511:0]     regroupCacheLine_0 = dataInMem;
  wire [511:0]     res = regroupCacheLine_0;
  wire [1023:0]    lo_lo = {512'h0, res};
  wire [2047:0]    lo = {1024'h0, lo_lo};
  wire [4095:0]    regroupLoadData_0_0 = {2048'h0, lo};
  wire [31:0]      dataInMem_lo_lo_lo_lo_lo_1 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1, dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [31:0]      dataInMem_lo_lo_lo_lo_hi_1 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3, dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [63:0]      dataInMem_lo_lo_lo_lo_1 = {dataInMem_lo_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_lo_lo_hi_lo_1 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5, dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [31:0]      dataInMem_lo_lo_lo_hi_hi_1 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7, dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [63:0]      dataInMem_lo_lo_lo_hi_1 = {dataInMem_lo_lo_lo_hi_hi_1, dataInMem_lo_lo_lo_hi_lo_1};
  wire [127:0]     dataInMem_lo_lo_lo_1 = {dataInMem_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_lo_hi_lo_lo_1 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9, dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [31:0]      dataInMem_lo_lo_hi_lo_hi_1 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11, dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [63:0]      dataInMem_lo_lo_hi_lo_1 = {dataInMem_lo_lo_hi_lo_hi_1, dataInMem_lo_lo_hi_lo_lo_1};
  wire [31:0]      dataInMem_lo_lo_hi_hi_lo_1 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13, dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [31:0]      dataInMem_lo_lo_hi_hi_hi_1 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15, dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [63:0]      dataInMem_lo_lo_hi_hi_1 = {dataInMem_lo_lo_hi_hi_hi_1, dataInMem_lo_lo_hi_hi_lo_1};
  wire [127:0]     dataInMem_lo_lo_hi_1 = {dataInMem_lo_lo_hi_hi_1, dataInMem_lo_lo_hi_lo_1};
  wire [255:0]     dataInMem_lo_lo_1 = {dataInMem_lo_lo_hi_1, dataInMem_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_lo_lo_lo_1 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17, dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [31:0]      dataInMem_lo_hi_lo_lo_hi_1 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19, dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [63:0]      dataInMem_lo_hi_lo_lo_1 = {dataInMem_lo_hi_lo_lo_hi_1, dataInMem_lo_hi_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_lo_hi_lo_1 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21, dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [31:0]      dataInMem_lo_hi_lo_hi_hi_1 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23, dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [63:0]      dataInMem_lo_hi_lo_hi_1 = {dataInMem_lo_hi_lo_hi_hi_1, dataInMem_lo_hi_lo_hi_lo_1};
  wire [127:0]     dataInMem_lo_hi_lo_1 = {dataInMem_lo_hi_lo_hi_1, dataInMem_lo_hi_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_hi_lo_lo_1 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25, dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [31:0]      dataInMem_lo_hi_hi_lo_hi_1 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27, dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [63:0]      dataInMem_lo_hi_hi_lo_1 = {dataInMem_lo_hi_hi_lo_hi_1, dataInMem_lo_hi_hi_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_hi_hi_lo_1 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29, dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [31:0]      dataInMem_lo_hi_hi_hi_hi_1 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31, dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [63:0]      dataInMem_lo_hi_hi_hi_1 = {dataInMem_lo_hi_hi_hi_hi_1, dataInMem_lo_hi_hi_hi_lo_1};
  wire [127:0]     dataInMem_lo_hi_hi_1 = {dataInMem_lo_hi_hi_hi_1, dataInMem_lo_hi_hi_lo_1};
  wire [255:0]     dataInMem_lo_hi_1 = {dataInMem_lo_hi_hi_1, dataInMem_lo_hi_lo_1};
  wire [511:0]     dataInMem_lo_1 = {dataInMem_lo_hi_1, dataInMem_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_lo_lo_lo_1 = {dataRegroupBySew_1_33, dataRegroupBySew_0_33, dataRegroupBySew_1_32, dataRegroupBySew_0_32};
  wire [31:0]      dataInMem_hi_lo_lo_lo_hi_1 = {dataRegroupBySew_1_35, dataRegroupBySew_0_35, dataRegroupBySew_1_34, dataRegroupBySew_0_34};
  wire [63:0]      dataInMem_hi_lo_lo_lo_1 = {dataInMem_hi_lo_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_lo_hi_lo_1 = {dataRegroupBySew_1_37, dataRegroupBySew_0_37, dataRegroupBySew_1_36, dataRegroupBySew_0_36};
  wire [31:0]      dataInMem_hi_lo_lo_hi_hi_1 = {dataRegroupBySew_1_39, dataRegroupBySew_0_39, dataRegroupBySew_1_38, dataRegroupBySew_0_38};
  wire [63:0]      dataInMem_hi_lo_lo_hi_1 = {dataInMem_hi_lo_lo_hi_hi_1, dataInMem_hi_lo_lo_hi_lo_1};
  wire [127:0]     dataInMem_hi_lo_lo_1 = {dataInMem_hi_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_hi_lo_lo_1 = {dataRegroupBySew_1_41, dataRegroupBySew_0_41, dataRegroupBySew_1_40, dataRegroupBySew_0_40};
  wire [31:0]      dataInMem_hi_lo_hi_lo_hi_1 = {dataRegroupBySew_1_43, dataRegroupBySew_0_43, dataRegroupBySew_1_42, dataRegroupBySew_0_42};
  wire [63:0]      dataInMem_hi_lo_hi_lo_1 = {dataInMem_hi_lo_hi_lo_hi_1, dataInMem_hi_lo_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_hi_hi_lo_1 = {dataRegroupBySew_1_45, dataRegroupBySew_0_45, dataRegroupBySew_1_44, dataRegroupBySew_0_44};
  wire [31:0]      dataInMem_hi_lo_hi_hi_hi_1 = {dataRegroupBySew_1_47, dataRegroupBySew_0_47, dataRegroupBySew_1_46, dataRegroupBySew_0_46};
  wire [63:0]      dataInMem_hi_lo_hi_hi_1 = {dataInMem_hi_lo_hi_hi_hi_1, dataInMem_hi_lo_hi_hi_lo_1};
  wire [127:0]     dataInMem_hi_lo_hi_1 = {dataInMem_hi_lo_hi_hi_1, dataInMem_hi_lo_hi_lo_1};
  wire [255:0]     dataInMem_hi_lo_1 = {dataInMem_hi_lo_hi_1, dataInMem_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_lo_lo_lo_1 = {dataRegroupBySew_1_49, dataRegroupBySew_0_49, dataRegroupBySew_1_48, dataRegroupBySew_0_48};
  wire [31:0]      dataInMem_hi_hi_lo_lo_hi_1 = {dataRegroupBySew_1_51, dataRegroupBySew_0_51, dataRegroupBySew_1_50, dataRegroupBySew_0_50};
  wire [63:0]      dataInMem_hi_hi_lo_lo_1 = {dataInMem_hi_hi_lo_lo_hi_1, dataInMem_hi_hi_lo_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_lo_hi_lo_1 = {dataRegroupBySew_1_53, dataRegroupBySew_0_53, dataRegroupBySew_1_52, dataRegroupBySew_0_52};
  wire [31:0]      dataInMem_hi_hi_lo_hi_hi_1 = {dataRegroupBySew_1_55, dataRegroupBySew_0_55, dataRegroupBySew_1_54, dataRegroupBySew_0_54};
  wire [63:0]      dataInMem_hi_hi_lo_hi_1 = {dataInMem_hi_hi_lo_hi_hi_1, dataInMem_hi_hi_lo_hi_lo_1};
  wire [127:0]     dataInMem_hi_hi_lo_1 = {dataInMem_hi_hi_lo_hi_1, dataInMem_hi_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_hi_lo_lo_1 = {dataRegroupBySew_1_57, dataRegroupBySew_0_57, dataRegroupBySew_1_56, dataRegroupBySew_0_56};
  wire [31:0]      dataInMem_hi_hi_hi_lo_hi_1 = {dataRegroupBySew_1_59, dataRegroupBySew_0_59, dataRegroupBySew_1_58, dataRegroupBySew_0_58};
  wire [63:0]      dataInMem_hi_hi_hi_lo_1 = {dataInMem_hi_hi_hi_lo_hi_1, dataInMem_hi_hi_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_hi_hi_lo_1 = {dataRegroupBySew_1_61, dataRegroupBySew_0_61, dataRegroupBySew_1_60, dataRegroupBySew_0_60};
  wire [31:0]      dataInMem_hi_hi_hi_hi_hi_1 = {dataRegroupBySew_1_63, dataRegroupBySew_0_63, dataRegroupBySew_1_62, dataRegroupBySew_0_62};
  wire [63:0]      dataInMem_hi_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_hi_lo_1};
  wire [127:0]     dataInMem_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_lo_1};
  wire [255:0]     dataInMem_hi_hi_1 = {dataInMem_hi_hi_hi_1, dataInMem_hi_hi_lo_1};
  wire [511:0]     dataInMem_hi_1 = {dataInMem_hi_hi_1, dataInMem_hi_lo_1};
  wire [1023:0]    dataInMem_1 = {dataInMem_hi_1, dataInMem_lo_1};
  wire [511:0]     regroupCacheLine_1_0 = dataInMem_1[511:0];
  wire [511:0]     regroupCacheLine_1_1 = dataInMem_1[1023:512];
  wire [511:0]     res_8 = regroupCacheLine_1_0;
  wire [511:0]     res_9 = regroupCacheLine_1_1;
  wire [1023:0]    lo_lo_1 = {res_9, res_8};
  wire [2047:0]    lo_1 = {1024'h0, lo_lo_1};
  wire [4095:0]    regroupLoadData_0_1 = {2048'h0, lo_1};
  wire [15:0]      _GEN_5 = {dataRegroupBySew_2_0, dataRegroupBySew_1_0};
  wire [15:0]      dataInMem_hi_2;
  assign dataInMem_hi_2 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_5;
  assign dataInMem_lo_hi_5 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_70;
  assign dataInMem_lo_hi_70 = _GEN_5;
  wire [15:0]      _GEN_6 = {dataRegroupBySew_2_1, dataRegroupBySew_1_1};
  wire [15:0]      dataInMem_hi_3;
  assign dataInMem_hi_3 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_6;
  assign dataInMem_lo_hi_6 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_71;
  assign dataInMem_lo_hi_71 = _GEN_6;
  wire [15:0]      _GEN_7 = {dataRegroupBySew_2_2, dataRegroupBySew_1_2};
  wire [15:0]      dataInMem_hi_4;
  assign dataInMem_hi_4 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_7;
  assign dataInMem_lo_hi_7 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_72;
  assign dataInMem_lo_hi_72 = _GEN_7;
  wire [15:0]      _GEN_8 = {dataRegroupBySew_2_3, dataRegroupBySew_1_3};
  wire [15:0]      dataInMem_hi_5;
  assign dataInMem_hi_5 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_8;
  assign dataInMem_lo_hi_8 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_73;
  assign dataInMem_lo_hi_73 = _GEN_8;
  wire [15:0]      _GEN_9 = {dataRegroupBySew_2_4, dataRegroupBySew_1_4};
  wire [15:0]      dataInMem_hi_6;
  assign dataInMem_hi_6 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_9;
  assign dataInMem_lo_hi_9 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_74;
  assign dataInMem_lo_hi_74 = _GEN_9;
  wire [15:0]      _GEN_10 = {dataRegroupBySew_2_5, dataRegroupBySew_1_5};
  wire [15:0]      dataInMem_hi_7;
  assign dataInMem_hi_7 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_10;
  assign dataInMem_lo_hi_10 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_75;
  assign dataInMem_lo_hi_75 = _GEN_10;
  wire [15:0]      _GEN_11 = {dataRegroupBySew_2_6, dataRegroupBySew_1_6};
  wire [15:0]      dataInMem_hi_8;
  assign dataInMem_hi_8 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_11;
  assign dataInMem_lo_hi_11 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_76;
  assign dataInMem_lo_hi_76 = _GEN_11;
  wire [15:0]      _GEN_12 = {dataRegroupBySew_2_7, dataRegroupBySew_1_7};
  wire [15:0]      dataInMem_hi_9;
  assign dataInMem_hi_9 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_12;
  assign dataInMem_lo_hi_12 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_77;
  assign dataInMem_lo_hi_77 = _GEN_12;
  wire [15:0]      _GEN_13 = {dataRegroupBySew_2_8, dataRegroupBySew_1_8};
  wire [15:0]      dataInMem_hi_10;
  assign dataInMem_hi_10 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_13;
  assign dataInMem_lo_hi_13 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_78;
  assign dataInMem_lo_hi_78 = _GEN_13;
  wire [15:0]      _GEN_14 = {dataRegroupBySew_2_9, dataRegroupBySew_1_9};
  wire [15:0]      dataInMem_hi_11;
  assign dataInMem_hi_11 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_14;
  assign dataInMem_lo_hi_14 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_79;
  assign dataInMem_lo_hi_79 = _GEN_14;
  wire [15:0]      _GEN_15 = {dataRegroupBySew_2_10, dataRegroupBySew_1_10};
  wire [15:0]      dataInMem_hi_12;
  assign dataInMem_hi_12 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_15;
  assign dataInMem_lo_hi_15 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_80;
  assign dataInMem_lo_hi_80 = _GEN_15;
  wire [15:0]      _GEN_16 = {dataRegroupBySew_2_11, dataRegroupBySew_1_11};
  wire [15:0]      dataInMem_hi_13;
  assign dataInMem_hi_13 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_16;
  assign dataInMem_lo_hi_16 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_81;
  assign dataInMem_lo_hi_81 = _GEN_16;
  wire [15:0]      _GEN_17 = {dataRegroupBySew_2_12, dataRegroupBySew_1_12};
  wire [15:0]      dataInMem_hi_14;
  assign dataInMem_hi_14 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_17;
  assign dataInMem_lo_hi_17 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_82;
  assign dataInMem_lo_hi_82 = _GEN_17;
  wire [15:0]      _GEN_18 = {dataRegroupBySew_2_13, dataRegroupBySew_1_13};
  wire [15:0]      dataInMem_hi_15;
  assign dataInMem_hi_15 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_18;
  assign dataInMem_lo_hi_18 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_83;
  assign dataInMem_lo_hi_83 = _GEN_18;
  wire [15:0]      _GEN_19 = {dataRegroupBySew_2_14, dataRegroupBySew_1_14};
  wire [15:0]      dataInMem_hi_16;
  assign dataInMem_hi_16 = _GEN_19;
  wire [15:0]      dataInMem_lo_hi_19;
  assign dataInMem_lo_hi_19 = _GEN_19;
  wire [15:0]      dataInMem_lo_hi_84;
  assign dataInMem_lo_hi_84 = _GEN_19;
  wire [15:0]      _GEN_20 = {dataRegroupBySew_2_15, dataRegroupBySew_1_15};
  wire [15:0]      dataInMem_hi_17;
  assign dataInMem_hi_17 = _GEN_20;
  wire [15:0]      dataInMem_lo_hi_20;
  assign dataInMem_lo_hi_20 = _GEN_20;
  wire [15:0]      dataInMem_lo_hi_85;
  assign dataInMem_lo_hi_85 = _GEN_20;
  wire [15:0]      _GEN_21 = {dataRegroupBySew_2_16, dataRegroupBySew_1_16};
  wire [15:0]      dataInMem_hi_18;
  assign dataInMem_hi_18 = _GEN_21;
  wire [15:0]      dataInMem_lo_hi_21;
  assign dataInMem_lo_hi_21 = _GEN_21;
  wire [15:0]      dataInMem_lo_hi_86;
  assign dataInMem_lo_hi_86 = _GEN_21;
  wire [15:0]      _GEN_22 = {dataRegroupBySew_2_17, dataRegroupBySew_1_17};
  wire [15:0]      dataInMem_hi_19;
  assign dataInMem_hi_19 = _GEN_22;
  wire [15:0]      dataInMem_lo_hi_22;
  assign dataInMem_lo_hi_22 = _GEN_22;
  wire [15:0]      dataInMem_lo_hi_87;
  assign dataInMem_lo_hi_87 = _GEN_22;
  wire [15:0]      _GEN_23 = {dataRegroupBySew_2_18, dataRegroupBySew_1_18};
  wire [15:0]      dataInMem_hi_20;
  assign dataInMem_hi_20 = _GEN_23;
  wire [15:0]      dataInMem_lo_hi_23;
  assign dataInMem_lo_hi_23 = _GEN_23;
  wire [15:0]      dataInMem_lo_hi_88;
  assign dataInMem_lo_hi_88 = _GEN_23;
  wire [15:0]      _GEN_24 = {dataRegroupBySew_2_19, dataRegroupBySew_1_19};
  wire [15:0]      dataInMem_hi_21;
  assign dataInMem_hi_21 = _GEN_24;
  wire [15:0]      dataInMem_lo_hi_24;
  assign dataInMem_lo_hi_24 = _GEN_24;
  wire [15:0]      dataInMem_lo_hi_89;
  assign dataInMem_lo_hi_89 = _GEN_24;
  wire [15:0]      _GEN_25 = {dataRegroupBySew_2_20, dataRegroupBySew_1_20};
  wire [15:0]      dataInMem_hi_22;
  assign dataInMem_hi_22 = _GEN_25;
  wire [15:0]      dataInMem_lo_hi_25;
  assign dataInMem_lo_hi_25 = _GEN_25;
  wire [15:0]      dataInMem_lo_hi_90;
  assign dataInMem_lo_hi_90 = _GEN_25;
  wire [15:0]      _GEN_26 = {dataRegroupBySew_2_21, dataRegroupBySew_1_21};
  wire [15:0]      dataInMem_hi_23;
  assign dataInMem_hi_23 = _GEN_26;
  wire [15:0]      dataInMem_lo_hi_26;
  assign dataInMem_lo_hi_26 = _GEN_26;
  wire [15:0]      dataInMem_lo_hi_91;
  assign dataInMem_lo_hi_91 = _GEN_26;
  wire [15:0]      _GEN_27 = {dataRegroupBySew_2_22, dataRegroupBySew_1_22};
  wire [15:0]      dataInMem_hi_24;
  assign dataInMem_hi_24 = _GEN_27;
  wire [15:0]      dataInMem_lo_hi_27;
  assign dataInMem_lo_hi_27 = _GEN_27;
  wire [15:0]      dataInMem_lo_hi_92;
  assign dataInMem_lo_hi_92 = _GEN_27;
  wire [15:0]      _GEN_28 = {dataRegroupBySew_2_23, dataRegroupBySew_1_23};
  wire [15:0]      dataInMem_hi_25;
  assign dataInMem_hi_25 = _GEN_28;
  wire [15:0]      dataInMem_lo_hi_28;
  assign dataInMem_lo_hi_28 = _GEN_28;
  wire [15:0]      dataInMem_lo_hi_93;
  assign dataInMem_lo_hi_93 = _GEN_28;
  wire [15:0]      _GEN_29 = {dataRegroupBySew_2_24, dataRegroupBySew_1_24};
  wire [15:0]      dataInMem_hi_26;
  assign dataInMem_hi_26 = _GEN_29;
  wire [15:0]      dataInMem_lo_hi_29;
  assign dataInMem_lo_hi_29 = _GEN_29;
  wire [15:0]      dataInMem_lo_hi_94;
  assign dataInMem_lo_hi_94 = _GEN_29;
  wire [15:0]      _GEN_30 = {dataRegroupBySew_2_25, dataRegroupBySew_1_25};
  wire [15:0]      dataInMem_hi_27;
  assign dataInMem_hi_27 = _GEN_30;
  wire [15:0]      dataInMem_lo_hi_30;
  assign dataInMem_lo_hi_30 = _GEN_30;
  wire [15:0]      dataInMem_lo_hi_95;
  assign dataInMem_lo_hi_95 = _GEN_30;
  wire [15:0]      _GEN_31 = {dataRegroupBySew_2_26, dataRegroupBySew_1_26};
  wire [15:0]      dataInMem_hi_28;
  assign dataInMem_hi_28 = _GEN_31;
  wire [15:0]      dataInMem_lo_hi_31;
  assign dataInMem_lo_hi_31 = _GEN_31;
  wire [15:0]      dataInMem_lo_hi_96;
  assign dataInMem_lo_hi_96 = _GEN_31;
  wire [15:0]      _GEN_32 = {dataRegroupBySew_2_27, dataRegroupBySew_1_27};
  wire [15:0]      dataInMem_hi_29;
  assign dataInMem_hi_29 = _GEN_32;
  wire [15:0]      dataInMem_lo_hi_32;
  assign dataInMem_lo_hi_32 = _GEN_32;
  wire [15:0]      dataInMem_lo_hi_97;
  assign dataInMem_lo_hi_97 = _GEN_32;
  wire [15:0]      _GEN_33 = {dataRegroupBySew_2_28, dataRegroupBySew_1_28};
  wire [15:0]      dataInMem_hi_30;
  assign dataInMem_hi_30 = _GEN_33;
  wire [15:0]      dataInMem_lo_hi_33;
  assign dataInMem_lo_hi_33 = _GEN_33;
  wire [15:0]      dataInMem_lo_hi_98;
  assign dataInMem_lo_hi_98 = _GEN_33;
  wire [15:0]      _GEN_34 = {dataRegroupBySew_2_29, dataRegroupBySew_1_29};
  wire [15:0]      dataInMem_hi_31;
  assign dataInMem_hi_31 = _GEN_34;
  wire [15:0]      dataInMem_lo_hi_34;
  assign dataInMem_lo_hi_34 = _GEN_34;
  wire [15:0]      dataInMem_lo_hi_99;
  assign dataInMem_lo_hi_99 = _GEN_34;
  wire [15:0]      _GEN_35 = {dataRegroupBySew_2_30, dataRegroupBySew_1_30};
  wire [15:0]      dataInMem_hi_32;
  assign dataInMem_hi_32 = _GEN_35;
  wire [15:0]      dataInMem_lo_hi_35;
  assign dataInMem_lo_hi_35 = _GEN_35;
  wire [15:0]      dataInMem_lo_hi_100;
  assign dataInMem_lo_hi_100 = _GEN_35;
  wire [15:0]      _GEN_36 = {dataRegroupBySew_2_31, dataRegroupBySew_1_31};
  wire [15:0]      dataInMem_hi_33;
  assign dataInMem_hi_33 = _GEN_36;
  wire [15:0]      dataInMem_lo_hi_36;
  assign dataInMem_lo_hi_36 = _GEN_36;
  wire [15:0]      dataInMem_lo_hi_101;
  assign dataInMem_lo_hi_101 = _GEN_36;
  wire [15:0]      _GEN_37 = {dataRegroupBySew_2_32, dataRegroupBySew_1_32};
  wire [15:0]      dataInMem_hi_34;
  assign dataInMem_hi_34 = _GEN_37;
  wire [15:0]      dataInMem_lo_hi_37;
  assign dataInMem_lo_hi_37 = _GEN_37;
  wire [15:0]      dataInMem_lo_hi_102;
  assign dataInMem_lo_hi_102 = _GEN_37;
  wire [15:0]      _GEN_38 = {dataRegroupBySew_2_33, dataRegroupBySew_1_33};
  wire [15:0]      dataInMem_hi_35;
  assign dataInMem_hi_35 = _GEN_38;
  wire [15:0]      dataInMem_lo_hi_38;
  assign dataInMem_lo_hi_38 = _GEN_38;
  wire [15:0]      dataInMem_lo_hi_103;
  assign dataInMem_lo_hi_103 = _GEN_38;
  wire [15:0]      _GEN_39 = {dataRegroupBySew_2_34, dataRegroupBySew_1_34};
  wire [15:0]      dataInMem_hi_36;
  assign dataInMem_hi_36 = _GEN_39;
  wire [15:0]      dataInMem_lo_hi_39;
  assign dataInMem_lo_hi_39 = _GEN_39;
  wire [15:0]      dataInMem_lo_hi_104;
  assign dataInMem_lo_hi_104 = _GEN_39;
  wire [15:0]      _GEN_40 = {dataRegroupBySew_2_35, dataRegroupBySew_1_35};
  wire [15:0]      dataInMem_hi_37;
  assign dataInMem_hi_37 = _GEN_40;
  wire [15:0]      dataInMem_lo_hi_40;
  assign dataInMem_lo_hi_40 = _GEN_40;
  wire [15:0]      dataInMem_lo_hi_105;
  assign dataInMem_lo_hi_105 = _GEN_40;
  wire [15:0]      _GEN_41 = {dataRegroupBySew_2_36, dataRegroupBySew_1_36};
  wire [15:0]      dataInMem_hi_38;
  assign dataInMem_hi_38 = _GEN_41;
  wire [15:0]      dataInMem_lo_hi_41;
  assign dataInMem_lo_hi_41 = _GEN_41;
  wire [15:0]      dataInMem_lo_hi_106;
  assign dataInMem_lo_hi_106 = _GEN_41;
  wire [15:0]      _GEN_42 = {dataRegroupBySew_2_37, dataRegroupBySew_1_37};
  wire [15:0]      dataInMem_hi_39;
  assign dataInMem_hi_39 = _GEN_42;
  wire [15:0]      dataInMem_lo_hi_42;
  assign dataInMem_lo_hi_42 = _GEN_42;
  wire [15:0]      dataInMem_lo_hi_107;
  assign dataInMem_lo_hi_107 = _GEN_42;
  wire [15:0]      _GEN_43 = {dataRegroupBySew_2_38, dataRegroupBySew_1_38};
  wire [15:0]      dataInMem_hi_40;
  assign dataInMem_hi_40 = _GEN_43;
  wire [15:0]      dataInMem_lo_hi_43;
  assign dataInMem_lo_hi_43 = _GEN_43;
  wire [15:0]      dataInMem_lo_hi_108;
  assign dataInMem_lo_hi_108 = _GEN_43;
  wire [15:0]      _GEN_44 = {dataRegroupBySew_2_39, dataRegroupBySew_1_39};
  wire [15:0]      dataInMem_hi_41;
  assign dataInMem_hi_41 = _GEN_44;
  wire [15:0]      dataInMem_lo_hi_44;
  assign dataInMem_lo_hi_44 = _GEN_44;
  wire [15:0]      dataInMem_lo_hi_109;
  assign dataInMem_lo_hi_109 = _GEN_44;
  wire [15:0]      _GEN_45 = {dataRegroupBySew_2_40, dataRegroupBySew_1_40};
  wire [15:0]      dataInMem_hi_42;
  assign dataInMem_hi_42 = _GEN_45;
  wire [15:0]      dataInMem_lo_hi_45;
  assign dataInMem_lo_hi_45 = _GEN_45;
  wire [15:0]      dataInMem_lo_hi_110;
  assign dataInMem_lo_hi_110 = _GEN_45;
  wire [15:0]      _GEN_46 = {dataRegroupBySew_2_41, dataRegroupBySew_1_41};
  wire [15:0]      dataInMem_hi_43;
  assign dataInMem_hi_43 = _GEN_46;
  wire [15:0]      dataInMem_lo_hi_46;
  assign dataInMem_lo_hi_46 = _GEN_46;
  wire [15:0]      dataInMem_lo_hi_111;
  assign dataInMem_lo_hi_111 = _GEN_46;
  wire [15:0]      _GEN_47 = {dataRegroupBySew_2_42, dataRegroupBySew_1_42};
  wire [15:0]      dataInMem_hi_44;
  assign dataInMem_hi_44 = _GEN_47;
  wire [15:0]      dataInMem_lo_hi_47;
  assign dataInMem_lo_hi_47 = _GEN_47;
  wire [15:0]      dataInMem_lo_hi_112;
  assign dataInMem_lo_hi_112 = _GEN_47;
  wire [15:0]      _GEN_48 = {dataRegroupBySew_2_43, dataRegroupBySew_1_43};
  wire [15:0]      dataInMem_hi_45;
  assign dataInMem_hi_45 = _GEN_48;
  wire [15:0]      dataInMem_lo_hi_48;
  assign dataInMem_lo_hi_48 = _GEN_48;
  wire [15:0]      dataInMem_lo_hi_113;
  assign dataInMem_lo_hi_113 = _GEN_48;
  wire [15:0]      _GEN_49 = {dataRegroupBySew_2_44, dataRegroupBySew_1_44};
  wire [15:0]      dataInMem_hi_46;
  assign dataInMem_hi_46 = _GEN_49;
  wire [15:0]      dataInMem_lo_hi_49;
  assign dataInMem_lo_hi_49 = _GEN_49;
  wire [15:0]      dataInMem_lo_hi_114;
  assign dataInMem_lo_hi_114 = _GEN_49;
  wire [15:0]      _GEN_50 = {dataRegroupBySew_2_45, dataRegroupBySew_1_45};
  wire [15:0]      dataInMem_hi_47;
  assign dataInMem_hi_47 = _GEN_50;
  wire [15:0]      dataInMem_lo_hi_50;
  assign dataInMem_lo_hi_50 = _GEN_50;
  wire [15:0]      dataInMem_lo_hi_115;
  assign dataInMem_lo_hi_115 = _GEN_50;
  wire [15:0]      _GEN_51 = {dataRegroupBySew_2_46, dataRegroupBySew_1_46};
  wire [15:0]      dataInMem_hi_48;
  assign dataInMem_hi_48 = _GEN_51;
  wire [15:0]      dataInMem_lo_hi_51;
  assign dataInMem_lo_hi_51 = _GEN_51;
  wire [15:0]      dataInMem_lo_hi_116;
  assign dataInMem_lo_hi_116 = _GEN_51;
  wire [15:0]      _GEN_52 = {dataRegroupBySew_2_47, dataRegroupBySew_1_47};
  wire [15:0]      dataInMem_hi_49;
  assign dataInMem_hi_49 = _GEN_52;
  wire [15:0]      dataInMem_lo_hi_52;
  assign dataInMem_lo_hi_52 = _GEN_52;
  wire [15:0]      dataInMem_lo_hi_117;
  assign dataInMem_lo_hi_117 = _GEN_52;
  wire [15:0]      _GEN_53 = {dataRegroupBySew_2_48, dataRegroupBySew_1_48};
  wire [15:0]      dataInMem_hi_50;
  assign dataInMem_hi_50 = _GEN_53;
  wire [15:0]      dataInMem_lo_hi_53;
  assign dataInMem_lo_hi_53 = _GEN_53;
  wire [15:0]      dataInMem_lo_hi_118;
  assign dataInMem_lo_hi_118 = _GEN_53;
  wire [15:0]      _GEN_54 = {dataRegroupBySew_2_49, dataRegroupBySew_1_49};
  wire [15:0]      dataInMem_hi_51;
  assign dataInMem_hi_51 = _GEN_54;
  wire [15:0]      dataInMem_lo_hi_54;
  assign dataInMem_lo_hi_54 = _GEN_54;
  wire [15:0]      dataInMem_lo_hi_119;
  assign dataInMem_lo_hi_119 = _GEN_54;
  wire [15:0]      _GEN_55 = {dataRegroupBySew_2_50, dataRegroupBySew_1_50};
  wire [15:0]      dataInMem_hi_52;
  assign dataInMem_hi_52 = _GEN_55;
  wire [15:0]      dataInMem_lo_hi_55;
  assign dataInMem_lo_hi_55 = _GEN_55;
  wire [15:0]      dataInMem_lo_hi_120;
  assign dataInMem_lo_hi_120 = _GEN_55;
  wire [15:0]      _GEN_56 = {dataRegroupBySew_2_51, dataRegroupBySew_1_51};
  wire [15:0]      dataInMem_hi_53;
  assign dataInMem_hi_53 = _GEN_56;
  wire [15:0]      dataInMem_lo_hi_56;
  assign dataInMem_lo_hi_56 = _GEN_56;
  wire [15:0]      dataInMem_lo_hi_121;
  assign dataInMem_lo_hi_121 = _GEN_56;
  wire [15:0]      _GEN_57 = {dataRegroupBySew_2_52, dataRegroupBySew_1_52};
  wire [15:0]      dataInMem_hi_54;
  assign dataInMem_hi_54 = _GEN_57;
  wire [15:0]      dataInMem_lo_hi_57;
  assign dataInMem_lo_hi_57 = _GEN_57;
  wire [15:0]      dataInMem_lo_hi_122;
  assign dataInMem_lo_hi_122 = _GEN_57;
  wire [15:0]      _GEN_58 = {dataRegroupBySew_2_53, dataRegroupBySew_1_53};
  wire [15:0]      dataInMem_hi_55;
  assign dataInMem_hi_55 = _GEN_58;
  wire [15:0]      dataInMem_lo_hi_58;
  assign dataInMem_lo_hi_58 = _GEN_58;
  wire [15:0]      dataInMem_lo_hi_123;
  assign dataInMem_lo_hi_123 = _GEN_58;
  wire [15:0]      _GEN_59 = {dataRegroupBySew_2_54, dataRegroupBySew_1_54};
  wire [15:0]      dataInMem_hi_56;
  assign dataInMem_hi_56 = _GEN_59;
  wire [15:0]      dataInMem_lo_hi_59;
  assign dataInMem_lo_hi_59 = _GEN_59;
  wire [15:0]      dataInMem_lo_hi_124;
  assign dataInMem_lo_hi_124 = _GEN_59;
  wire [15:0]      _GEN_60 = {dataRegroupBySew_2_55, dataRegroupBySew_1_55};
  wire [15:0]      dataInMem_hi_57;
  assign dataInMem_hi_57 = _GEN_60;
  wire [15:0]      dataInMem_lo_hi_60;
  assign dataInMem_lo_hi_60 = _GEN_60;
  wire [15:0]      dataInMem_lo_hi_125;
  assign dataInMem_lo_hi_125 = _GEN_60;
  wire [15:0]      _GEN_61 = {dataRegroupBySew_2_56, dataRegroupBySew_1_56};
  wire [15:0]      dataInMem_hi_58;
  assign dataInMem_hi_58 = _GEN_61;
  wire [15:0]      dataInMem_lo_hi_61;
  assign dataInMem_lo_hi_61 = _GEN_61;
  wire [15:0]      dataInMem_lo_hi_126;
  assign dataInMem_lo_hi_126 = _GEN_61;
  wire [15:0]      _GEN_62 = {dataRegroupBySew_2_57, dataRegroupBySew_1_57};
  wire [15:0]      dataInMem_hi_59;
  assign dataInMem_hi_59 = _GEN_62;
  wire [15:0]      dataInMem_lo_hi_62;
  assign dataInMem_lo_hi_62 = _GEN_62;
  wire [15:0]      dataInMem_lo_hi_127;
  assign dataInMem_lo_hi_127 = _GEN_62;
  wire [15:0]      _GEN_63 = {dataRegroupBySew_2_58, dataRegroupBySew_1_58};
  wire [15:0]      dataInMem_hi_60;
  assign dataInMem_hi_60 = _GEN_63;
  wire [15:0]      dataInMem_lo_hi_63;
  assign dataInMem_lo_hi_63 = _GEN_63;
  wire [15:0]      dataInMem_lo_hi_128;
  assign dataInMem_lo_hi_128 = _GEN_63;
  wire [15:0]      _GEN_64 = {dataRegroupBySew_2_59, dataRegroupBySew_1_59};
  wire [15:0]      dataInMem_hi_61;
  assign dataInMem_hi_61 = _GEN_64;
  wire [15:0]      dataInMem_lo_hi_64;
  assign dataInMem_lo_hi_64 = _GEN_64;
  wire [15:0]      dataInMem_lo_hi_129;
  assign dataInMem_lo_hi_129 = _GEN_64;
  wire [15:0]      _GEN_65 = {dataRegroupBySew_2_60, dataRegroupBySew_1_60};
  wire [15:0]      dataInMem_hi_62;
  assign dataInMem_hi_62 = _GEN_65;
  wire [15:0]      dataInMem_lo_hi_65;
  assign dataInMem_lo_hi_65 = _GEN_65;
  wire [15:0]      dataInMem_lo_hi_130;
  assign dataInMem_lo_hi_130 = _GEN_65;
  wire [15:0]      _GEN_66 = {dataRegroupBySew_2_61, dataRegroupBySew_1_61};
  wire [15:0]      dataInMem_hi_63;
  assign dataInMem_hi_63 = _GEN_66;
  wire [15:0]      dataInMem_lo_hi_66;
  assign dataInMem_lo_hi_66 = _GEN_66;
  wire [15:0]      dataInMem_lo_hi_131;
  assign dataInMem_lo_hi_131 = _GEN_66;
  wire [15:0]      _GEN_67 = {dataRegroupBySew_2_62, dataRegroupBySew_1_62};
  wire [15:0]      dataInMem_hi_64;
  assign dataInMem_hi_64 = _GEN_67;
  wire [15:0]      dataInMem_lo_hi_67;
  assign dataInMem_lo_hi_67 = _GEN_67;
  wire [15:0]      dataInMem_lo_hi_132;
  assign dataInMem_lo_hi_132 = _GEN_67;
  wire [15:0]      _GEN_68 = {dataRegroupBySew_2_63, dataRegroupBySew_1_63};
  wire [15:0]      dataInMem_hi_65;
  assign dataInMem_hi_65 = _GEN_68;
  wire [15:0]      dataInMem_lo_hi_68;
  assign dataInMem_lo_hi_68 = _GEN_68;
  wire [15:0]      dataInMem_lo_hi_133;
  assign dataInMem_lo_hi_133 = _GEN_68;
  wire [47:0]      dataInMem_lo_lo_lo_lo_lo_2 = {dataInMem_hi_3, dataRegroupBySew_0_1, dataInMem_hi_2, dataRegroupBySew_0_0};
  wire [47:0]      dataInMem_lo_lo_lo_lo_hi_2 = {dataInMem_hi_5, dataRegroupBySew_0_3, dataInMem_hi_4, dataRegroupBySew_0_2};
  wire [95:0]      dataInMem_lo_lo_lo_lo_2 = {dataInMem_lo_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_lo_lo_hi_lo_2 = {dataInMem_hi_7, dataRegroupBySew_0_5, dataInMem_hi_6, dataRegroupBySew_0_4};
  wire [47:0]      dataInMem_lo_lo_lo_hi_hi_2 = {dataInMem_hi_9, dataRegroupBySew_0_7, dataInMem_hi_8, dataRegroupBySew_0_6};
  wire [95:0]      dataInMem_lo_lo_lo_hi_2 = {dataInMem_lo_lo_lo_hi_hi_2, dataInMem_lo_lo_lo_hi_lo_2};
  wire [191:0]     dataInMem_lo_lo_lo_2 = {dataInMem_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_lo_hi_lo_lo_2 = {dataInMem_hi_11, dataRegroupBySew_0_9, dataInMem_hi_10, dataRegroupBySew_0_8};
  wire [47:0]      dataInMem_lo_lo_hi_lo_hi_2 = {dataInMem_hi_13, dataRegroupBySew_0_11, dataInMem_hi_12, dataRegroupBySew_0_10};
  wire [95:0]      dataInMem_lo_lo_hi_lo_2 = {dataInMem_lo_lo_hi_lo_hi_2, dataInMem_lo_lo_hi_lo_lo_2};
  wire [47:0]      dataInMem_lo_lo_hi_hi_lo_2 = {dataInMem_hi_15, dataRegroupBySew_0_13, dataInMem_hi_14, dataRegroupBySew_0_12};
  wire [47:0]      dataInMem_lo_lo_hi_hi_hi_2 = {dataInMem_hi_17, dataRegroupBySew_0_15, dataInMem_hi_16, dataRegroupBySew_0_14};
  wire [95:0]      dataInMem_lo_lo_hi_hi_2 = {dataInMem_lo_lo_hi_hi_hi_2, dataInMem_lo_lo_hi_hi_lo_2};
  wire [191:0]     dataInMem_lo_lo_hi_2 = {dataInMem_lo_lo_hi_hi_2, dataInMem_lo_lo_hi_lo_2};
  wire [383:0]     dataInMem_lo_lo_2 = {dataInMem_lo_lo_hi_2, dataInMem_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_lo_lo_lo_2 = {dataInMem_hi_19, dataRegroupBySew_0_17, dataInMem_hi_18, dataRegroupBySew_0_16};
  wire [47:0]      dataInMem_lo_hi_lo_lo_hi_2 = {dataInMem_hi_21, dataRegroupBySew_0_19, dataInMem_hi_20, dataRegroupBySew_0_18};
  wire [95:0]      dataInMem_lo_hi_lo_lo_2 = {dataInMem_lo_hi_lo_lo_hi_2, dataInMem_lo_hi_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_lo_hi_lo_2 = {dataInMem_hi_23, dataRegroupBySew_0_21, dataInMem_hi_22, dataRegroupBySew_0_20};
  wire [47:0]      dataInMem_lo_hi_lo_hi_hi_2 = {dataInMem_hi_25, dataRegroupBySew_0_23, dataInMem_hi_24, dataRegroupBySew_0_22};
  wire [95:0]      dataInMem_lo_hi_lo_hi_2 = {dataInMem_lo_hi_lo_hi_hi_2, dataInMem_lo_hi_lo_hi_lo_2};
  wire [191:0]     dataInMem_lo_hi_lo_2 = {dataInMem_lo_hi_lo_hi_2, dataInMem_lo_hi_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_hi_lo_lo_2 = {dataInMem_hi_27, dataRegroupBySew_0_25, dataInMem_hi_26, dataRegroupBySew_0_24};
  wire [47:0]      dataInMem_lo_hi_hi_lo_hi_2 = {dataInMem_hi_29, dataRegroupBySew_0_27, dataInMem_hi_28, dataRegroupBySew_0_26};
  wire [95:0]      dataInMem_lo_hi_hi_lo_2 = {dataInMem_lo_hi_hi_lo_hi_2, dataInMem_lo_hi_hi_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_hi_hi_lo_2 = {dataInMem_hi_31, dataRegroupBySew_0_29, dataInMem_hi_30, dataRegroupBySew_0_28};
  wire [47:0]      dataInMem_lo_hi_hi_hi_hi_2 = {dataInMem_hi_33, dataRegroupBySew_0_31, dataInMem_hi_32, dataRegroupBySew_0_30};
  wire [95:0]      dataInMem_lo_hi_hi_hi_2 = {dataInMem_lo_hi_hi_hi_hi_2, dataInMem_lo_hi_hi_hi_lo_2};
  wire [191:0]     dataInMem_lo_hi_hi_2 = {dataInMem_lo_hi_hi_hi_2, dataInMem_lo_hi_hi_lo_2};
  wire [383:0]     dataInMem_lo_hi_2 = {dataInMem_lo_hi_hi_2, dataInMem_lo_hi_lo_2};
  wire [767:0]     dataInMem_lo_2 = {dataInMem_lo_hi_2, dataInMem_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_lo_lo_lo_2 = {dataInMem_hi_35, dataRegroupBySew_0_33, dataInMem_hi_34, dataRegroupBySew_0_32};
  wire [47:0]      dataInMem_hi_lo_lo_lo_hi_2 = {dataInMem_hi_37, dataRegroupBySew_0_35, dataInMem_hi_36, dataRegroupBySew_0_34};
  wire [95:0]      dataInMem_hi_lo_lo_lo_2 = {dataInMem_hi_lo_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_lo_hi_lo_2 = {dataInMem_hi_39, dataRegroupBySew_0_37, dataInMem_hi_38, dataRegroupBySew_0_36};
  wire [47:0]      dataInMem_hi_lo_lo_hi_hi_2 = {dataInMem_hi_41, dataRegroupBySew_0_39, dataInMem_hi_40, dataRegroupBySew_0_38};
  wire [95:0]      dataInMem_hi_lo_lo_hi_2 = {dataInMem_hi_lo_lo_hi_hi_2, dataInMem_hi_lo_lo_hi_lo_2};
  wire [191:0]     dataInMem_hi_lo_lo_2 = {dataInMem_hi_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_hi_lo_lo_2 = {dataInMem_hi_43, dataRegroupBySew_0_41, dataInMem_hi_42, dataRegroupBySew_0_40};
  wire [47:0]      dataInMem_hi_lo_hi_lo_hi_2 = {dataInMem_hi_45, dataRegroupBySew_0_43, dataInMem_hi_44, dataRegroupBySew_0_42};
  wire [95:0]      dataInMem_hi_lo_hi_lo_2 = {dataInMem_hi_lo_hi_lo_hi_2, dataInMem_hi_lo_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_hi_hi_lo_2 = {dataInMem_hi_47, dataRegroupBySew_0_45, dataInMem_hi_46, dataRegroupBySew_0_44};
  wire [47:0]      dataInMem_hi_lo_hi_hi_hi_2 = {dataInMem_hi_49, dataRegroupBySew_0_47, dataInMem_hi_48, dataRegroupBySew_0_46};
  wire [95:0]      dataInMem_hi_lo_hi_hi_2 = {dataInMem_hi_lo_hi_hi_hi_2, dataInMem_hi_lo_hi_hi_lo_2};
  wire [191:0]     dataInMem_hi_lo_hi_2 = {dataInMem_hi_lo_hi_hi_2, dataInMem_hi_lo_hi_lo_2};
  wire [383:0]     dataInMem_hi_lo_2 = {dataInMem_hi_lo_hi_2, dataInMem_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_lo_lo_lo_2 = {dataInMem_hi_51, dataRegroupBySew_0_49, dataInMem_hi_50, dataRegroupBySew_0_48};
  wire [47:0]      dataInMem_hi_hi_lo_lo_hi_2 = {dataInMem_hi_53, dataRegroupBySew_0_51, dataInMem_hi_52, dataRegroupBySew_0_50};
  wire [95:0]      dataInMem_hi_hi_lo_lo_2 = {dataInMem_hi_hi_lo_lo_hi_2, dataInMem_hi_hi_lo_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_lo_hi_lo_2 = {dataInMem_hi_55, dataRegroupBySew_0_53, dataInMem_hi_54, dataRegroupBySew_0_52};
  wire [47:0]      dataInMem_hi_hi_lo_hi_hi_2 = {dataInMem_hi_57, dataRegroupBySew_0_55, dataInMem_hi_56, dataRegroupBySew_0_54};
  wire [95:0]      dataInMem_hi_hi_lo_hi_2 = {dataInMem_hi_hi_lo_hi_hi_2, dataInMem_hi_hi_lo_hi_lo_2};
  wire [191:0]     dataInMem_hi_hi_lo_2 = {dataInMem_hi_hi_lo_hi_2, dataInMem_hi_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_hi_lo_lo_2 = {dataInMem_hi_59, dataRegroupBySew_0_57, dataInMem_hi_58, dataRegroupBySew_0_56};
  wire [47:0]      dataInMem_hi_hi_hi_lo_hi_2 = {dataInMem_hi_61, dataRegroupBySew_0_59, dataInMem_hi_60, dataRegroupBySew_0_58};
  wire [95:0]      dataInMem_hi_hi_hi_lo_2 = {dataInMem_hi_hi_hi_lo_hi_2, dataInMem_hi_hi_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_hi_hi_lo_2 = {dataInMem_hi_63, dataRegroupBySew_0_61, dataInMem_hi_62, dataRegroupBySew_0_60};
  wire [47:0]      dataInMem_hi_hi_hi_hi_hi_2 = {dataInMem_hi_65, dataRegroupBySew_0_63, dataInMem_hi_64, dataRegroupBySew_0_62};
  wire [95:0]      dataInMem_hi_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_hi_lo_2};
  wire [191:0]     dataInMem_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_lo_2};
  wire [383:0]     dataInMem_hi_hi_2 = {dataInMem_hi_hi_hi_2, dataInMem_hi_hi_lo_2};
  wire [767:0]     dataInMem_hi_66 = {dataInMem_hi_hi_2, dataInMem_hi_lo_2};
  wire [1535:0]    dataInMem_2 = {dataInMem_hi_66, dataInMem_lo_2};
  wire [511:0]     regroupCacheLine_2_0 = dataInMem_2[511:0];
  wire [511:0]     regroupCacheLine_2_1 = dataInMem_2[1023:512];
  wire [511:0]     regroupCacheLine_2_2 = dataInMem_2[1535:1024];
  wire [511:0]     res_16 = regroupCacheLine_2_0;
  wire [511:0]     res_17 = regroupCacheLine_2_1;
  wire [511:0]     res_18 = regroupCacheLine_2_2;
  wire [1023:0]    lo_lo_2 = {res_17, res_16};
  wire [1023:0]    lo_hi_2 = {512'h0, res_18};
  wire [2047:0]    lo_2 = {lo_hi_2, lo_lo_2};
  wire [4095:0]    regroupLoadData_0_2 = {2048'h0, lo_2};
  wire [15:0]      _GEN_69 = {dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_3;
  assign dataInMem_lo_3 = _GEN_69;
  wire [15:0]      dataInMem_lo_68;
  assign dataInMem_lo_68 = _GEN_69;
  wire [15:0]      dataInMem_lo_lo_7;
  assign dataInMem_lo_lo_7 = _GEN_69;
  wire [15:0]      _GEN_70 = {dataRegroupBySew_3_0, dataRegroupBySew_2_0};
  wire [15:0]      dataInMem_hi_67;
  assign dataInMem_hi_67 = _GEN_70;
  wire [15:0]      dataInMem_lo_hi_135;
  assign dataInMem_lo_hi_135 = _GEN_70;
  wire [15:0]      _GEN_71 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_lo_4;
  assign dataInMem_lo_4 = _GEN_71;
  wire [15:0]      dataInMem_lo_69;
  assign dataInMem_lo_69 = _GEN_71;
  wire [15:0]      dataInMem_lo_lo_8;
  assign dataInMem_lo_lo_8 = _GEN_71;
  wire [15:0]      _GEN_72 = {dataRegroupBySew_3_1, dataRegroupBySew_2_1};
  wire [15:0]      dataInMem_hi_68;
  assign dataInMem_hi_68 = _GEN_72;
  wire [15:0]      dataInMem_lo_hi_136;
  assign dataInMem_lo_hi_136 = _GEN_72;
  wire [15:0]      _GEN_73 = {dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_lo_5;
  assign dataInMem_lo_5 = _GEN_73;
  wire [15:0]      dataInMem_lo_70;
  assign dataInMem_lo_70 = _GEN_73;
  wire [15:0]      dataInMem_lo_lo_9;
  assign dataInMem_lo_lo_9 = _GEN_73;
  wire [15:0]      _GEN_74 = {dataRegroupBySew_3_2, dataRegroupBySew_2_2};
  wire [15:0]      dataInMem_hi_69;
  assign dataInMem_hi_69 = _GEN_74;
  wire [15:0]      dataInMem_lo_hi_137;
  assign dataInMem_lo_hi_137 = _GEN_74;
  wire [15:0]      _GEN_75 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_lo_6;
  assign dataInMem_lo_6 = _GEN_75;
  wire [15:0]      dataInMem_lo_71;
  assign dataInMem_lo_71 = _GEN_75;
  wire [15:0]      dataInMem_lo_lo_10;
  assign dataInMem_lo_lo_10 = _GEN_75;
  wire [15:0]      _GEN_76 = {dataRegroupBySew_3_3, dataRegroupBySew_2_3};
  wire [15:0]      dataInMem_hi_70;
  assign dataInMem_hi_70 = _GEN_76;
  wire [15:0]      dataInMem_lo_hi_138;
  assign dataInMem_lo_hi_138 = _GEN_76;
  wire [15:0]      _GEN_77 = {dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_7;
  assign dataInMem_lo_7 = _GEN_77;
  wire [15:0]      dataInMem_lo_72;
  assign dataInMem_lo_72 = _GEN_77;
  wire [15:0]      dataInMem_lo_lo_11;
  assign dataInMem_lo_lo_11 = _GEN_77;
  wire [15:0]      _GEN_78 = {dataRegroupBySew_3_4, dataRegroupBySew_2_4};
  wire [15:0]      dataInMem_hi_71;
  assign dataInMem_hi_71 = _GEN_78;
  wire [15:0]      dataInMem_lo_hi_139;
  assign dataInMem_lo_hi_139 = _GEN_78;
  wire [15:0]      _GEN_79 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_lo_8;
  assign dataInMem_lo_8 = _GEN_79;
  wire [15:0]      dataInMem_lo_73;
  assign dataInMem_lo_73 = _GEN_79;
  wire [15:0]      dataInMem_lo_lo_12;
  assign dataInMem_lo_lo_12 = _GEN_79;
  wire [15:0]      _GEN_80 = {dataRegroupBySew_3_5, dataRegroupBySew_2_5};
  wire [15:0]      dataInMem_hi_72;
  assign dataInMem_hi_72 = _GEN_80;
  wire [15:0]      dataInMem_lo_hi_140;
  assign dataInMem_lo_hi_140 = _GEN_80;
  wire [15:0]      _GEN_81 = {dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_lo_9;
  assign dataInMem_lo_9 = _GEN_81;
  wire [15:0]      dataInMem_lo_74;
  assign dataInMem_lo_74 = _GEN_81;
  wire [15:0]      dataInMem_lo_lo_13;
  assign dataInMem_lo_lo_13 = _GEN_81;
  wire [15:0]      _GEN_82 = {dataRegroupBySew_3_6, dataRegroupBySew_2_6};
  wire [15:0]      dataInMem_hi_73;
  assign dataInMem_hi_73 = _GEN_82;
  wire [15:0]      dataInMem_lo_hi_141;
  assign dataInMem_lo_hi_141 = _GEN_82;
  wire [15:0]      _GEN_83 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_lo_10;
  assign dataInMem_lo_10 = _GEN_83;
  wire [15:0]      dataInMem_lo_75;
  assign dataInMem_lo_75 = _GEN_83;
  wire [15:0]      dataInMem_lo_lo_14;
  assign dataInMem_lo_lo_14 = _GEN_83;
  wire [15:0]      _GEN_84 = {dataRegroupBySew_3_7, dataRegroupBySew_2_7};
  wire [15:0]      dataInMem_hi_74;
  assign dataInMem_hi_74 = _GEN_84;
  wire [15:0]      dataInMem_lo_hi_142;
  assign dataInMem_lo_hi_142 = _GEN_84;
  wire [15:0]      _GEN_85 = {dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_lo_11;
  assign dataInMem_lo_11 = _GEN_85;
  wire [15:0]      dataInMem_lo_76;
  assign dataInMem_lo_76 = _GEN_85;
  wire [15:0]      dataInMem_lo_lo_15;
  assign dataInMem_lo_lo_15 = _GEN_85;
  wire [15:0]      _GEN_86 = {dataRegroupBySew_3_8, dataRegroupBySew_2_8};
  wire [15:0]      dataInMem_hi_75;
  assign dataInMem_hi_75 = _GEN_86;
  wire [15:0]      dataInMem_lo_hi_143;
  assign dataInMem_lo_hi_143 = _GEN_86;
  wire [15:0]      _GEN_87 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_lo_12;
  assign dataInMem_lo_12 = _GEN_87;
  wire [15:0]      dataInMem_lo_77;
  assign dataInMem_lo_77 = _GEN_87;
  wire [15:0]      dataInMem_lo_lo_16;
  assign dataInMem_lo_lo_16 = _GEN_87;
  wire [15:0]      _GEN_88 = {dataRegroupBySew_3_9, dataRegroupBySew_2_9};
  wire [15:0]      dataInMem_hi_76;
  assign dataInMem_hi_76 = _GEN_88;
  wire [15:0]      dataInMem_lo_hi_144;
  assign dataInMem_lo_hi_144 = _GEN_88;
  wire [15:0]      _GEN_89 = {dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_lo_13;
  assign dataInMem_lo_13 = _GEN_89;
  wire [15:0]      dataInMem_lo_78;
  assign dataInMem_lo_78 = _GEN_89;
  wire [15:0]      dataInMem_lo_lo_17;
  assign dataInMem_lo_lo_17 = _GEN_89;
  wire [15:0]      _GEN_90 = {dataRegroupBySew_3_10, dataRegroupBySew_2_10};
  wire [15:0]      dataInMem_hi_77;
  assign dataInMem_hi_77 = _GEN_90;
  wire [15:0]      dataInMem_lo_hi_145;
  assign dataInMem_lo_hi_145 = _GEN_90;
  wire [15:0]      _GEN_91 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_lo_14;
  assign dataInMem_lo_14 = _GEN_91;
  wire [15:0]      dataInMem_lo_79;
  assign dataInMem_lo_79 = _GEN_91;
  wire [15:0]      dataInMem_lo_lo_18;
  assign dataInMem_lo_lo_18 = _GEN_91;
  wire [15:0]      _GEN_92 = {dataRegroupBySew_3_11, dataRegroupBySew_2_11};
  wire [15:0]      dataInMem_hi_78;
  assign dataInMem_hi_78 = _GEN_92;
  wire [15:0]      dataInMem_lo_hi_146;
  assign dataInMem_lo_hi_146 = _GEN_92;
  wire [15:0]      _GEN_93 = {dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_lo_15;
  assign dataInMem_lo_15 = _GEN_93;
  wire [15:0]      dataInMem_lo_80;
  assign dataInMem_lo_80 = _GEN_93;
  wire [15:0]      dataInMem_lo_lo_19;
  assign dataInMem_lo_lo_19 = _GEN_93;
  wire [15:0]      _GEN_94 = {dataRegroupBySew_3_12, dataRegroupBySew_2_12};
  wire [15:0]      dataInMem_hi_79;
  assign dataInMem_hi_79 = _GEN_94;
  wire [15:0]      dataInMem_lo_hi_147;
  assign dataInMem_lo_hi_147 = _GEN_94;
  wire [15:0]      _GEN_95 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_lo_16;
  assign dataInMem_lo_16 = _GEN_95;
  wire [15:0]      dataInMem_lo_81;
  assign dataInMem_lo_81 = _GEN_95;
  wire [15:0]      dataInMem_lo_lo_20;
  assign dataInMem_lo_lo_20 = _GEN_95;
  wire [15:0]      _GEN_96 = {dataRegroupBySew_3_13, dataRegroupBySew_2_13};
  wire [15:0]      dataInMem_hi_80;
  assign dataInMem_hi_80 = _GEN_96;
  wire [15:0]      dataInMem_lo_hi_148;
  assign dataInMem_lo_hi_148 = _GEN_96;
  wire [15:0]      _GEN_97 = {dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_lo_17;
  assign dataInMem_lo_17 = _GEN_97;
  wire [15:0]      dataInMem_lo_82;
  assign dataInMem_lo_82 = _GEN_97;
  wire [15:0]      dataInMem_lo_lo_21;
  assign dataInMem_lo_lo_21 = _GEN_97;
  wire [15:0]      _GEN_98 = {dataRegroupBySew_3_14, dataRegroupBySew_2_14};
  wire [15:0]      dataInMem_hi_81;
  assign dataInMem_hi_81 = _GEN_98;
  wire [15:0]      dataInMem_lo_hi_149;
  assign dataInMem_lo_hi_149 = _GEN_98;
  wire [15:0]      _GEN_99 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_lo_18;
  assign dataInMem_lo_18 = _GEN_99;
  wire [15:0]      dataInMem_lo_83;
  assign dataInMem_lo_83 = _GEN_99;
  wire [15:0]      dataInMem_lo_lo_22;
  assign dataInMem_lo_lo_22 = _GEN_99;
  wire [15:0]      _GEN_100 = {dataRegroupBySew_3_15, dataRegroupBySew_2_15};
  wire [15:0]      dataInMem_hi_82;
  assign dataInMem_hi_82 = _GEN_100;
  wire [15:0]      dataInMem_lo_hi_150;
  assign dataInMem_lo_hi_150 = _GEN_100;
  wire [15:0]      _GEN_101 = {dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_lo_19;
  assign dataInMem_lo_19 = _GEN_101;
  wire [15:0]      dataInMem_lo_84;
  assign dataInMem_lo_84 = _GEN_101;
  wire [15:0]      dataInMem_lo_lo_23;
  assign dataInMem_lo_lo_23 = _GEN_101;
  wire [15:0]      _GEN_102 = {dataRegroupBySew_3_16, dataRegroupBySew_2_16};
  wire [15:0]      dataInMem_hi_83;
  assign dataInMem_hi_83 = _GEN_102;
  wire [15:0]      dataInMem_lo_hi_151;
  assign dataInMem_lo_hi_151 = _GEN_102;
  wire [15:0]      _GEN_103 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17};
  wire [15:0]      dataInMem_lo_20;
  assign dataInMem_lo_20 = _GEN_103;
  wire [15:0]      dataInMem_lo_85;
  assign dataInMem_lo_85 = _GEN_103;
  wire [15:0]      dataInMem_lo_lo_24;
  assign dataInMem_lo_lo_24 = _GEN_103;
  wire [15:0]      _GEN_104 = {dataRegroupBySew_3_17, dataRegroupBySew_2_17};
  wire [15:0]      dataInMem_hi_84;
  assign dataInMem_hi_84 = _GEN_104;
  wire [15:0]      dataInMem_lo_hi_152;
  assign dataInMem_lo_hi_152 = _GEN_104;
  wire [15:0]      _GEN_105 = {dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [15:0]      dataInMem_lo_21;
  assign dataInMem_lo_21 = _GEN_105;
  wire [15:0]      dataInMem_lo_86;
  assign dataInMem_lo_86 = _GEN_105;
  wire [15:0]      dataInMem_lo_lo_25;
  assign dataInMem_lo_lo_25 = _GEN_105;
  wire [15:0]      _GEN_106 = {dataRegroupBySew_3_18, dataRegroupBySew_2_18};
  wire [15:0]      dataInMem_hi_85;
  assign dataInMem_hi_85 = _GEN_106;
  wire [15:0]      dataInMem_lo_hi_153;
  assign dataInMem_lo_hi_153 = _GEN_106;
  wire [15:0]      _GEN_107 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19};
  wire [15:0]      dataInMem_lo_22;
  assign dataInMem_lo_22 = _GEN_107;
  wire [15:0]      dataInMem_lo_87;
  assign dataInMem_lo_87 = _GEN_107;
  wire [15:0]      dataInMem_lo_lo_26;
  assign dataInMem_lo_lo_26 = _GEN_107;
  wire [15:0]      _GEN_108 = {dataRegroupBySew_3_19, dataRegroupBySew_2_19};
  wire [15:0]      dataInMem_hi_86;
  assign dataInMem_hi_86 = _GEN_108;
  wire [15:0]      dataInMem_lo_hi_154;
  assign dataInMem_lo_hi_154 = _GEN_108;
  wire [15:0]      _GEN_109 = {dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_lo_23;
  assign dataInMem_lo_23 = _GEN_109;
  wire [15:0]      dataInMem_lo_88;
  assign dataInMem_lo_88 = _GEN_109;
  wire [15:0]      dataInMem_lo_lo_27;
  assign dataInMem_lo_lo_27 = _GEN_109;
  wire [15:0]      _GEN_110 = {dataRegroupBySew_3_20, dataRegroupBySew_2_20};
  wire [15:0]      dataInMem_hi_87;
  assign dataInMem_hi_87 = _GEN_110;
  wire [15:0]      dataInMem_lo_hi_155;
  assign dataInMem_lo_hi_155 = _GEN_110;
  wire [15:0]      _GEN_111 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21};
  wire [15:0]      dataInMem_lo_24;
  assign dataInMem_lo_24 = _GEN_111;
  wire [15:0]      dataInMem_lo_89;
  assign dataInMem_lo_89 = _GEN_111;
  wire [15:0]      dataInMem_lo_lo_28;
  assign dataInMem_lo_lo_28 = _GEN_111;
  wire [15:0]      _GEN_112 = {dataRegroupBySew_3_21, dataRegroupBySew_2_21};
  wire [15:0]      dataInMem_hi_88;
  assign dataInMem_hi_88 = _GEN_112;
  wire [15:0]      dataInMem_lo_hi_156;
  assign dataInMem_lo_hi_156 = _GEN_112;
  wire [15:0]      _GEN_113 = {dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [15:0]      dataInMem_lo_25;
  assign dataInMem_lo_25 = _GEN_113;
  wire [15:0]      dataInMem_lo_90;
  assign dataInMem_lo_90 = _GEN_113;
  wire [15:0]      dataInMem_lo_lo_29;
  assign dataInMem_lo_lo_29 = _GEN_113;
  wire [15:0]      _GEN_114 = {dataRegroupBySew_3_22, dataRegroupBySew_2_22};
  wire [15:0]      dataInMem_hi_89;
  assign dataInMem_hi_89 = _GEN_114;
  wire [15:0]      dataInMem_lo_hi_157;
  assign dataInMem_lo_hi_157 = _GEN_114;
  wire [15:0]      _GEN_115 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23};
  wire [15:0]      dataInMem_lo_26;
  assign dataInMem_lo_26 = _GEN_115;
  wire [15:0]      dataInMem_lo_91;
  assign dataInMem_lo_91 = _GEN_115;
  wire [15:0]      dataInMem_lo_lo_30;
  assign dataInMem_lo_lo_30 = _GEN_115;
  wire [15:0]      _GEN_116 = {dataRegroupBySew_3_23, dataRegroupBySew_2_23};
  wire [15:0]      dataInMem_hi_90;
  assign dataInMem_hi_90 = _GEN_116;
  wire [15:0]      dataInMem_lo_hi_158;
  assign dataInMem_lo_hi_158 = _GEN_116;
  wire [15:0]      _GEN_117 = {dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_lo_27;
  assign dataInMem_lo_27 = _GEN_117;
  wire [15:0]      dataInMem_lo_92;
  assign dataInMem_lo_92 = _GEN_117;
  wire [15:0]      dataInMem_lo_lo_31;
  assign dataInMem_lo_lo_31 = _GEN_117;
  wire [15:0]      _GEN_118 = {dataRegroupBySew_3_24, dataRegroupBySew_2_24};
  wire [15:0]      dataInMem_hi_91;
  assign dataInMem_hi_91 = _GEN_118;
  wire [15:0]      dataInMem_lo_hi_159;
  assign dataInMem_lo_hi_159 = _GEN_118;
  wire [15:0]      _GEN_119 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25};
  wire [15:0]      dataInMem_lo_28;
  assign dataInMem_lo_28 = _GEN_119;
  wire [15:0]      dataInMem_lo_93;
  assign dataInMem_lo_93 = _GEN_119;
  wire [15:0]      dataInMem_lo_lo_32;
  assign dataInMem_lo_lo_32 = _GEN_119;
  wire [15:0]      _GEN_120 = {dataRegroupBySew_3_25, dataRegroupBySew_2_25};
  wire [15:0]      dataInMem_hi_92;
  assign dataInMem_hi_92 = _GEN_120;
  wire [15:0]      dataInMem_lo_hi_160;
  assign dataInMem_lo_hi_160 = _GEN_120;
  wire [15:0]      _GEN_121 = {dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [15:0]      dataInMem_lo_29;
  assign dataInMem_lo_29 = _GEN_121;
  wire [15:0]      dataInMem_lo_94;
  assign dataInMem_lo_94 = _GEN_121;
  wire [15:0]      dataInMem_lo_lo_33;
  assign dataInMem_lo_lo_33 = _GEN_121;
  wire [15:0]      _GEN_122 = {dataRegroupBySew_3_26, dataRegroupBySew_2_26};
  wire [15:0]      dataInMem_hi_93;
  assign dataInMem_hi_93 = _GEN_122;
  wire [15:0]      dataInMem_lo_hi_161;
  assign dataInMem_lo_hi_161 = _GEN_122;
  wire [15:0]      _GEN_123 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27};
  wire [15:0]      dataInMem_lo_30;
  assign dataInMem_lo_30 = _GEN_123;
  wire [15:0]      dataInMem_lo_95;
  assign dataInMem_lo_95 = _GEN_123;
  wire [15:0]      dataInMem_lo_lo_34;
  assign dataInMem_lo_lo_34 = _GEN_123;
  wire [15:0]      _GEN_124 = {dataRegroupBySew_3_27, dataRegroupBySew_2_27};
  wire [15:0]      dataInMem_hi_94;
  assign dataInMem_hi_94 = _GEN_124;
  wire [15:0]      dataInMem_lo_hi_162;
  assign dataInMem_lo_hi_162 = _GEN_124;
  wire [15:0]      _GEN_125 = {dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_lo_31;
  assign dataInMem_lo_31 = _GEN_125;
  wire [15:0]      dataInMem_lo_96;
  assign dataInMem_lo_96 = _GEN_125;
  wire [15:0]      dataInMem_lo_lo_35;
  assign dataInMem_lo_lo_35 = _GEN_125;
  wire [15:0]      _GEN_126 = {dataRegroupBySew_3_28, dataRegroupBySew_2_28};
  wire [15:0]      dataInMem_hi_95;
  assign dataInMem_hi_95 = _GEN_126;
  wire [15:0]      dataInMem_lo_hi_163;
  assign dataInMem_lo_hi_163 = _GEN_126;
  wire [15:0]      _GEN_127 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29};
  wire [15:0]      dataInMem_lo_32;
  assign dataInMem_lo_32 = _GEN_127;
  wire [15:0]      dataInMem_lo_97;
  assign dataInMem_lo_97 = _GEN_127;
  wire [15:0]      dataInMem_lo_lo_36;
  assign dataInMem_lo_lo_36 = _GEN_127;
  wire [15:0]      _GEN_128 = {dataRegroupBySew_3_29, dataRegroupBySew_2_29};
  wire [15:0]      dataInMem_hi_96;
  assign dataInMem_hi_96 = _GEN_128;
  wire [15:0]      dataInMem_lo_hi_164;
  assign dataInMem_lo_hi_164 = _GEN_128;
  wire [15:0]      _GEN_129 = {dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [15:0]      dataInMem_lo_33;
  assign dataInMem_lo_33 = _GEN_129;
  wire [15:0]      dataInMem_lo_98;
  assign dataInMem_lo_98 = _GEN_129;
  wire [15:0]      dataInMem_lo_lo_37;
  assign dataInMem_lo_lo_37 = _GEN_129;
  wire [15:0]      _GEN_130 = {dataRegroupBySew_3_30, dataRegroupBySew_2_30};
  wire [15:0]      dataInMem_hi_97;
  assign dataInMem_hi_97 = _GEN_130;
  wire [15:0]      dataInMem_lo_hi_165;
  assign dataInMem_lo_hi_165 = _GEN_130;
  wire [15:0]      _GEN_131 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31};
  wire [15:0]      dataInMem_lo_34;
  assign dataInMem_lo_34 = _GEN_131;
  wire [15:0]      dataInMem_lo_99;
  assign dataInMem_lo_99 = _GEN_131;
  wire [15:0]      dataInMem_lo_lo_38;
  assign dataInMem_lo_lo_38 = _GEN_131;
  wire [15:0]      _GEN_132 = {dataRegroupBySew_3_31, dataRegroupBySew_2_31};
  wire [15:0]      dataInMem_hi_98;
  assign dataInMem_hi_98 = _GEN_132;
  wire [15:0]      dataInMem_lo_hi_166;
  assign dataInMem_lo_hi_166 = _GEN_132;
  wire [15:0]      _GEN_133 = {dataRegroupBySew_1_32, dataRegroupBySew_0_32};
  wire [15:0]      dataInMem_lo_35;
  assign dataInMem_lo_35 = _GEN_133;
  wire [15:0]      dataInMem_lo_100;
  assign dataInMem_lo_100 = _GEN_133;
  wire [15:0]      dataInMem_lo_lo_39;
  assign dataInMem_lo_lo_39 = _GEN_133;
  wire [15:0]      _GEN_134 = {dataRegroupBySew_3_32, dataRegroupBySew_2_32};
  wire [15:0]      dataInMem_hi_99;
  assign dataInMem_hi_99 = _GEN_134;
  wire [15:0]      dataInMem_lo_hi_167;
  assign dataInMem_lo_hi_167 = _GEN_134;
  wire [15:0]      _GEN_135 = {dataRegroupBySew_1_33, dataRegroupBySew_0_33};
  wire [15:0]      dataInMem_lo_36;
  assign dataInMem_lo_36 = _GEN_135;
  wire [15:0]      dataInMem_lo_101;
  assign dataInMem_lo_101 = _GEN_135;
  wire [15:0]      dataInMem_lo_lo_40;
  assign dataInMem_lo_lo_40 = _GEN_135;
  wire [15:0]      _GEN_136 = {dataRegroupBySew_3_33, dataRegroupBySew_2_33};
  wire [15:0]      dataInMem_hi_100;
  assign dataInMem_hi_100 = _GEN_136;
  wire [15:0]      dataInMem_lo_hi_168;
  assign dataInMem_lo_hi_168 = _GEN_136;
  wire [15:0]      _GEN_137 = {dataRegroupBySew_1_34, dataRegroupBySew_0_34};
  wire [15:0]      dataInMem_lo_37;
  assign dataInMem_lo_37 = _GEN_137;
  wire [15:0]      dataInMem_lo_102;
  assign dataInMem_lo_102 = _GEN_137;
  wire [15:0]      dataInMem_lo_lo_41;
  assign dataInMem_lo_lo_41 = _GEN_137;
  wire [15:0]      _GEN_138 = {dataRegroupBySew_3_34, dataRegroupBySew_2_34};
  wire [15:0]      dataInMem_hi_101;
  assign dataInMem_hi_101 = _GEN_138;
  wire [15:0]      dataInMem_lo_hi_169;
  assign dataInMem_lo_hi_169 = _GEN_138;
  wire [15:0]      _GEN_139 = {dataRegroupBySew_1_35, dataRegroupBySew_0_35};
  wire [15:0]      dataInMem_lo_38;
  assign dataInMem_lo_38 = _GEN_139;
  wire [15:0]      dataInMem_lo_103;
  assign dataInMem_lo_103 = _GEN_139;
  wire [15:0]      dataInMem_lo_lo_42;
  assign dataInMem_lo_lo_42 = _GEN_139;
  wire [15:0]      _GEN_140 = {dataRegroupBySew_3_35, dataRegroupBySew_2_35};
  wire [15:0]      dataInMem_hi_102;
  assign dataInMem_hi_102 = _GEN_140;
  wire [15:0]      dataInMem_lo_hi_170;
  assign dataInMem_lo_hi_170 = _GEN_140;
  wire [15:0]      _GEN_141 = {dataRegroupBySew_1_36, dataRegroupBySew_0_36};
  wire [15:0]      dataInMem_lo_39;
  assign dataInMem_lo_39 = _GEN_141;
  wire [15:0]      dataInMem_lo_104;
  assign dataInMem_lo_104 = _GEN_141;
  wire [15:0]      dataInMem_lo_lo_43;
  assign dataInMem_lo_lo_43 = _GEN_141;
  wire [15:0]      _GEN_142 = {dataRegroupBySew_3_36, dataRegroupBySew_2_36};
  wire [15:0]      dataInMem_hi_103;
  assign dataInMem_hi_103 = _GEN_142;
  wire [15:0]      dataInMem_lo_hi_171;
  assign dataInMem_lo_hi_171 = _GEN_142;
  wire [15:0]      _GEN_143 = {dataRegroupBySew_1_37, dataRegroupBySew_0_37};
  wire [15:0]      dataInMem_lo_40;
  assign dataInMem_lo_40 = _GEN_143;
  wire [15:0]      dataInMem_lo_105;
  assign dataInMem_lo_105 = _GEN_143;
  wire [15:0]      dataInMem_lo_lo_44;
  assign dataInMem_lo_lo_44 = _GEN_143;
  wire [15:0]      _GEN_144 = {dataRegroupBySew_3_37, dataRegroupBySew_2_37};
  wire [15:0]      dataInMem_hi_104;
  assign dataInMem_hi_104 = _GEN_144;
  wire [15:0]      dataInMem_lo_hi_172;
  assign dataInMem_lo_hi_172 = _GEN_144;
  wire [15:0]      _GEN_145 = {dataRegroupBySew_1_38, dataRegroupBySew_0_38};
  wire [15:0]      dataInMem_lo_41;
  assign dataInMem_lo_41 = _GEN_145;
  wire [15:0]      dataInMem_lo_106;
  assign dataInMem_lo_106 = _GEN_145;
  wire [15:0]      dataInMem_lo_lo_45;
  assign dataInMem_lo_lo_45 = _GEN_145;
  wire [15:0]      _GEN_146 = {dataRegroupBySew_3_38, dataRegroupBySew_2_38};
  wire [15:0]      dataInMem_hi_105;
  assign dataInMem_hi_105 = _GEN_146;
  wire [15:0]      dataInMem_lo_hi_173;
  assign dataInMem_lo_hi_173 = _GEN_146;
  wire [15:0]      _GEN_147 = {dataRegroupBySew_1_39, dataRegroupBySew_0_39};
  wire [15:0]      dataInMem_lo_42;
  assign dataInMem_lo_42 = _GEN_147;
  wire [15:0]      dataInMem_lo_107;
  assign dataInMem_lo_107 = _GEN_147;
  wire [15:0]      dataInMem_lo_lo_46;
  assign dataInMem_lo_lo_46 = _GEN_147;
  wire [15:0]      _GEN_148 = {dataRegroupBySew_3_39, dataRegroupBySew_2_39};
  wire [15:0]      dataInMem_hi_106;
  assign dataInMem_hi_106 = _GEN_148;
  wire [15:0]      dataInMem_lo_hi_174;
  assign dataInMem_lo_hi_174 = _GEN_148;
  wire [15:0]      _GEN_149 = {dataRegroupBySew_1_40, dataRegroupBySew_0_40};
  wire [15:0]      dataInMem_lo_43;
  assign dataInMem_lo_43 = _GEN_149;
  wire [15:0]      dataInMem_lo_108;
  assign dataInMem_lo_108 = _GEN_149;
  wire [15:0]      dataInMem_lo_lo_47;
  assign dataInMem_lo_lo_47 = _GEN_149;
  wire [15:0]      _GEN_150 = {dataRegroupBySew_3_40, dataRegroupBySew_2_40};
  wire [15:0]      dataInMem_hi_107;
  assign dataInMem_hi_107 = _GEN_150;
  wire [15:0]      dataInMem_lo_hi_175;
  assign dataInMem_lo_hi_175 = _GEN_150;
  wire [15:0]      _GEN_151 = {dataRegroupBySew_1_41, dataRegroupBySew_0_41};
  wire [15:0]      dataInMem_lo_44;
  assign dataInMem_lo_44 = _GEN_151;
  wire [15:0]      dataInMem_lo_109;
  assign dataInMem_lo_109 = _GEN_151;
  wire [15:0]      dataInMem_lo_lo_48;
  assign dataInMem_lo_lo_48 = _GEN_151;
  wire [15:0]      _GEN_152 = {dataRegroupBySew_3_41, dataRegroupBySew_2_41};
  wire [15:0]      dataInMem_hi_108;
  assign dataInMem_hi_108 = _GEN_152;
  wire [15:0]      dataInMem_lo_hi_176;
  assign dataInMem_lo_hi_176 = _GEN_152;
  wire [15:0]      _GEN_153 = {dataRegroupBySew_1_42, dataRegroupBySew_0_42};
  wire [15:0]      dataInMem_lo_45;
  assign dataInMem_lo_45 = _GEN_153;
  wire [15:0]      dataInMem_lo_110;
  assign dataInMem_lo_110 = _GEN_153;
  wire [15:0]      dataInMem_lo_lo_49;
  assign dataInMem_lo_lo_49 = _GEN_153;
  wire [15:0]      _GEN_154 = {dataRegroupBySew_3_42, dataRegroupBySew_2_42};
  wire [15:0]      dataInMem_hi_109;
  assign dataInMem_hi_109 = _GEN_154;
  wire [15:0]      dataInMem_lo_hi_177;
  assign dataInMem_lo_hi_177 = _GEN_154;
  wire [15:0]      _GEN_155 = {dataRegroupBySew_1_43, dataRegroupBySew_0_43};
  wire [15:0]      dataInMem_lo_46;
  assign dataInMem_lo_46 = _GEN_155;
  wire [15:0]      dataInMem_lo_111;
  assign dataInMem_lo_111 = _GEN_155;
  wire [15:0]      dataInMem_lo_lo_50;
  assign dataInMem_lo_lo_50 = _GEN_155;
  wire [15:0]      _GEN_156 = {dataRegroupBySew_3_43, dataRegroupBySew_2_43};
  wire [15:0]      dataInMem_hi_110;
  assign dataInMem_hi_110 = _GEN_156;
  wire [15:0]      dataInMem_lo_hi_178;
  assign dataInMem_lo_hi_178 = _GEN_156;
  wire [15:0]      _GEN_157 = {dataRegroupBySew_1_44, dataRegroupBySew_0_44};
  wire [15:0]      dataInMem_lo_47;
  assign dataInMem_lo_47 = _GEN_157;
  wire [15:0]      dataInMem_lo_112;
  assign dataInMem_lo_112 = _GEN_157;
  wire [15:0]      dataInMem_lo_lo_51;
  assign dataInMem_lo_lo_51 = _GEN_157;
  wire [15:0]      _GEN_158 = {dataRegroupBySew_3_44, dataRegroupBySew_2_44};
  wire [15:0]      dataInMem_hi_111;
  assign dataInMem_hi_111 = _GEN_158;
  wire [15:0]      dataInMem_lo_hi_179;
  assign dataInMem_lo_hi_179 = _GEN_158;
  wire [15:0]      _GEN_159 = {dataRegroupBySew_1_45, dataRegroupBySew_0_45};
  wire [15:0]      dataInMem_lo_48;
  assign dataInMem_lo_48 = _GEN_159;
  wire [15:0]      dataInMem_lo_113;
  assign dataInMem_lo_113 = _GEN_159;
  wire [15:0]      dataInMem_lo_lo_52;
  assign dataInMem_lo_lo_52 = _GEN_159;
  wire [15:0]      _GEN_160 = {dataRegroupBySew_3_45, dataRegroupBySew_2_45};
  wire [15:0]      dataInMem_hi_112;
  assign dataInMem_hi_112 = _GEN_160;
  wire [15:0]      dataInMem_lo_hi_180;
  assign dataInMem_lo_hi_180 = _GEN_160;
  wire [15:0]      _GEN_161 = {dataRegroupBySew_1_46, dataRegroupBySew_0_46};
  wire [15:0]      dataInMem_lo_49;
  assign dataInMem_lo_49 = _GEN_161;
  wire [15:0]      dataInMem_lo_114;
  assign dataInMem_lo_114 = _GEN_161;
  wire [15:0]      dataInMem_lo_lo_53;
  assign dataInMem_lo_lo_53 = _GEN_161;
  wire [15:0]      _GEN_162 = {dataRegroupBySew_3_46, dataRegroupBySew_2_46};
  wire [15:0]      dataInMem_hi_113;
  assign dataInMem_hi_113 = _GEN_162;
  wire [15:0]      dataInMem_lo_hi_181;
  assign dataInMem_lo_hi_181 = _GEN_162;
  wire [15:0]      _GEN_163 = {dataRegroupBySew_1_47, dataRegroupBySew_0_47};
  wire [15:0]      dataInMem_lo_50;
  assign dataInMem_lo_50 = _GEN_163;
  wire [15:0]      dataInMem_lo_115;
  assign dataInMem_lo_115 = _GEN_163;
  wire [15:0]      dataInMem_lo_lo_54;
  assign dataInMem_lo_lo_54 = _GEN_163;
  wire [15:0]      _GEN_164 = {dataRegroupBySew_3_47, dataRegroupBySew_2_47};
  wire [15:0]      dataInMem_hi_114;
  assign dataInMem_hi_114 = _GEN_164;
  wire [15:0]      dataInMem_lo_hi_182;
  assign dataInMem_lo_hi_182 = _GEN_164;
  wire [15:0]      _GEN_165 = {dataRegroupBySew_1_48, dataRegroupBySew_0_48};
  wire [15:0]      dataInMem_lo_51;
  assign dataInMem_lo_51 = _GEN_165;
  wire [15:0]      dataInMem_lo_116;
  assign dataInMem_lo_116 = _GEN_165;
  wire [15:0]      dataInMem_lo_lo_55;
  assign dataInMem_lo_lo_55 = _GEN_165;
  wire [15:0]      _GEN_166 = {dataRegroupBySew_3_48, dataRegroupBySew_2_48};
  wire [15:0]      dataInMem_hi_115;
  assign dataInMem_hi_115 = _GEN_166;
  wire [15:0]      dataInMem_lo_hi_183;
  assign dataInMem_lo_hi_183 = _GEN_166;
  wire [15:0]      _GEN_167 = {dataRegroupBySew_1_49, dataRegroupBySew_0_49};
  wire [15:0]      dataInMem_lo_52;
  assign dataInMem_lo_52 = _GEN_167;
  wire [15:0]      dataInMem_lo_117;
  assign dataInMem_lo_117 = _GEN_167;
  wire [15:0]      dataInMem_lo_lo_56;
  assign dataInMem_lo_lo_56 = _GEN_167;
  wire [15:0]      _GEN_168 = {dataRegroupBySew_3_49, dataRegroupBySew_2_49};
  wire [15:0]      dataInMem_hi_116;
  assign dataInMem_hi_116 = _GEN_168;
  wire [15:0]      dataInMem_lo_hi_184;
  assign dataInMem_lo_hi_184 = _GEN_168;
  wire [15:0]      _GEN_169 = {dataRegroupBySew_1_50, dataRegroupBySew_0_50};
  wire [15:0]      dataInMem_lo_53;
  assign dataInMem_lo_53 = _GEN_169;
  wire [15:0]      dataInMem_lo_118;
  assign dataInMem_lo_118 = _GEN_169;
  wire [15:0]      dataInMem_lo_lo_57;
  assign dataInMem_lo_lo_57 = _GEN_169;
  wire [15:0]      _GEN_170 = {dataRegroupBySew_3_50, dataRegroupBySew_2_50};
  wire [15:0]      dataInMem_hi_117;
  assign dataInMem_hi_117 = _GEN_170;
  wire [15:0]      dataInMem_lo_hi_185;
  assign dataInMem_lo_hi_185 = _GEN_170;
  wire [15:0]      _GEN_171 = {dataRegroupBySew_1_51, dataRegroupBySew_0_51};
  wire [15:0]      dataInMem_lo_54;
  assign dataInMem_lo_54 = _GEN_171;
  wire [15:0]      dataInMem_lo_119;
  assign dataInMem_lo_119 = _GEN_171;
  wire [15:0]      dataInMem_lo_lo_58;
  assign dataInMem_lo_lo_58 = _GEN_171;
  wire [15:0]      _GEN_172 = {dataRegroupBySew_3_51, dataRegroupBySew_2_51};
  wire [15:0]      dataInMem_hi_118;
  assign dataInMem_hi_118 = _GEN_172;
  wire [15:0]      dataInMem_lo_hi_186;
  assign dataInMem_lo_hi_186 = _GEN_172;
  wire [15:0]      _GEN_173 = {dataRegroupBySew_1_52, dataRegroupBySew_0_52};
  wire [15:0]      dataInMem_lo_55;
  assign dataInMem_lo_55 = _GEN_173;
  wire [15:0]      dataInMem_lo_120;
  assign dataInMem_lo_120 = _GEN_173;
  wire [15:0]      dataInMem_lo_lo_59;
  assign dataInMem_lo_lo_59 = _GEN_173;
  wire [15:0]      _GEN_174 = {dataRegroupBySew_3_52, dataRegroupBySew_2_52};
  wire [15:0]      dataInMem_hi_119;
  assign dataInMem_hi_119 = _GEN_174;
  wire [15:0]      dataInMem_lo_hi_187;
  assign dataInMem_lo_hi_187 = _GEN_174;
  wire [15:0]      _GEN_175 = {dataRegroupBySew_1_53, dataRegroupBySew_0_53};
  wire [15:0]      dataInMem_lo_56;
  assign dataInMem_lo_56 = _GEN_175;
  wire [15:0]      dataInMem_lo_121;
  assign dataInMem_lo_121 = _GEN_175;
  wire [15:0]      dataInMem_lo_lo_60;
  assign dataInMem_lo_lo_60 = _GEN_175;
  wire [15:0]      _GEN_176 = {dataRegroupBySew_3_53, dataRegroupBySew_2_53};
  wire [15:0]      dataInMem_hi_120;
  assign dataInMem_hi_120 = _GEN_176;
  wire [15:0]      dataInMem_lo_hi_188;
  assign dataInMem_lo_hi_188 = _GEN_176;
  wire [15:0]      _GEN_177 = {dataRegroupBySew_1_54, dataRegroupBySew_0_54};
  wire [15:0]      dataInMem_lo_57;
  assign dataInMem_lo_57 = _GEN_177;
  wire [15:0]      dataInMem_lo_122;
  assign dataInMem_lo_122 = _GEN_177;
  wire [15:0]      dataInMem_lo_lo_61;
  assign dataInMem_lo_lo_61 = _GEN_177;
  wire [15:0]      _GEN_178 = {dataRegroupBySew_3_54, dataRegroupBySew_2_54};
  wire [15:0]      dataInMem_hi_121;
  assign dataInMem_hi_121 = _GEN_178;
  wire [15:0]      dataInMem_lo_hi_189;
  assign dataInMem_lo_hi_189 = _GEN_178;
  wire [15:0]      _GEN_179 = {dataRegroupBySew_1_55, dataRegroupBySew_0_55};
  wire [15:0]      dataInMem_lo_58;
  assign dataInMem_lo_58 = _GEN_179;
  wire [15:0]      dataInMem_lo_123;
  assign dataInMem_lo_123 = _GEN_179;
  wire [15:0]      dataInMem_lo_lo_62;
  assign dataInMem_lo_lo_62 = _GEN_179;
  wire [15:0]      _GEN_180 = {dataRegroupBySew_3_55, dataRegroupBySew_2_55};
  wire [15:0]      dataInMem_hi_122;
  assign dataInMem_hi_122 = _GEN_180;
  wire [15:0]      dataInMem_lo_hi_190;
  assign dataInMem_lo_hi_190 = _GEN_180;
  wire [15:0]      _GEN_181 = {dataRegroupBySew_1_56, dataRegroupBySew_0_56};
  wire [15:0]      dataInMem_lo_59;
  assign dataInMem_lo_59 = _GEN_181;
  wire [15:0]      dataInMem_lo_124;
  assign dataInMem_lo_124 = _GEN_181;
  wire [15:0]      dataInMem_lo_lo_63;
  assign dataInMem_lo_lo_63 = _GEN_181;
  wire [15:0]      _GEN_182 = {dataRegroupBySew_3_56, dataRegroupBySew_2_56};
  wire [15:0]      dataInMem_hi_123;
  assign dataInMem_hi_123 = _GEN_182;
  wire [15:0]      dataInMem_lo_hi_191;
  assign dataInMem_lo_hi_191 = _GEN_182;
  wire [15:0]      _GEN_183 = {dataRegroupBySew_1_57, dataRegroupBySew_0_57};
  wire [15:0]      dataInMem_lo_60;
  assign dataInMem_lo_60 = _GEN_183;
  wire [15:0]      dataInMem_lo_125;
  assign dataInMem_lo_125 = _GEN_183;
  wire [15:0]      dataInMem_lo_lo_64;
  assign dataInMem_lo_lo_64 = _GEN_183;
  wire [15:0]      _GEN_184 = {dataRegroupBySew_3_57, dataRegroupBySew_2_57};
  wire [15:0]      dataInMem_hi_124;
  assign dataInMem_hi_124 = _GEN_184;
  wire [15:0]      dataInMem_lo_hi_192;
  assign dataInMem_lo_hi_192 = _GEN_184;
  wire [15:0]      _GEN_185 = {dataRegroupBySew_1_58, dataRegroupBySew_0_58};
  wire [15:0]      dataInMem_lo_61;
  assign dataInMem_lo_61 = _GEN_185;
  wire [15:0]      dataInMem_lo_126;
  assign dataInMem_lo_126 = _GEN_185;
  wire [15:0]      dataInMem_lo_lo_65;
  assign dataInMem_lo_lo_65 = _GEN_185;
  wire [15:0]      _GEN_186 = {dataRegroupBySew_3_58, dataRegroupBySew_2_58};
  wire [15:0]      dataInMem_hi_125;
  assign dataInMem_hi_125 = _GEN_186;
  wire [15:0]      dataInMem_lo_hi_193;
  assign dataInMem_lo_hi_193 = _GEN_186;
  wire [15:0]      _GEN_187 = {dataRegroupBySew_1_59, dataRegroupBySew_0_59};
  wire [15:0]      dataInMem_lo_62;
  assign dataInMem_lo_62 = _GEN_187;
  wire [15:0]      dataInMem_lo_127;
  assign dataInMem_lo_127 = _GEN_187;
  wire [15:0]      dataInMem_lo_lo_66;
  assign dataInMem_lo_lo_66 = _GEN_187;
  wire [15:0]      _GEN_188 = {dataRegroupBySew_3_59, dataRegroupBySew_2_59};
  wire [15:0]      dataInMem_hi_126;
  assign dataInMem_hi_126 = _GEN_188;
  wire [15:0]      dataInMem_lo_hi_194;
  assign dataInMem_lo_hi_194 = _GEN_188;
  wire [15:0]      _GEN_189 = {dataRegroupBySew_1_60, dataRegroupBySew_0_60};
  wire [15:0]      dataInMem_lo_63;
  assign dataInMem_lo_63 = _GEN_189;
  wire [15:0]      dataInMem_lo_128;
  assign dataInMem_lo_128 = _GEN_189;
  wire [15:0]      dataInMem_lo_lo_67;
  assign dataInMem_lo_lo_67 = _GEN_189;
  wire [15:0]      _GEN_190 = {dataRegroupBySew_3_60, dataRegroupBySew_2_60};
  wire [15:0]      dataInMem_hi_127;
  assign dataInMem_hi_127 = _GEN_190;
  wire [15:0]      dataInMem_lo_hi_195;
  assign dataInMem_lo_hi_195 = _GEN_190;
  wire [15:0]      _GEN_191 = {dataRegroupBySew_1_61, dataRegroupBySew_0_61};
  wire [15:0]      dataInMem_lo_64;
  assign dataInMem_lo_64 = _GEN_191;
  wire [15:0]      dataInMem_lo_129;
  assign dataInMem_lo_129 = _GEN_191;
  wire [15:0]      dataInMem_lo_lo_68;
  assign dataInMem_lo_lo_68 = _GEN_191;
  wire [15:0]      _GEN_192 = {dataRegroupBySew_3_61, dataRegroupBySew_2_61};
  wire [15:0]      dataInMem_hi_128;
  assign dataInMem_hi_128 = _GEN_192;
  wire [15:0]      dataInMem_lo_hi_196;
  assign dataInMem_lo_hi_196 = _GEN_192;
  wire [15:0]      _GEN_193 = {dataRegroupBySew_1_62, dataRegroupBySew_0_62};
  wire [15:0]      dataInMem_lo_65;
  assign dataInMem_lo_65 = _GEN_193;
  wire [15:0]      dataInMem_lo_130;
  assign dataInMem_lo_130 = _GEN_193;
  wire [15:0]      dataInMem_lo_lo_69;
  assign dataInMem_lo_lo_69 = _GEN_193;
  wire [15:0]      _GEN_194 = {dataRegroupBySew_3_62, dataRegroupBySew_2_62};
  wire [15:0]      dataInMem_hi_129;
  assign dataInMem_hi_129 = _GEN_194;
  wire [15:0]      dataInMem_lo_hi_197;
  assign dataInMem_lo_hi_197 = _GEN_194;
  wire [15:0]      _GEN_195 = {dataRegroupBySew_1_63, dataRegroupBySew_0_63};
  wire [15:0]      dataInMem_lo_66;
  assign dataInMem_lo_66 = _GEN_195;
  wire [15:0]      dataInMem_lo_131;
  assign dataInMem_lo_131 = _GEN_195;
  wire [15:0]      dataInMem_lo_lo_70;
  assign dataInMem_lo_lo_70 = _GEN_195;
  wire [15:0]      _GEN_196 = {dataRegroupBySew_3_63, dataRegroupBySew_2_63};
  wire [15:0]      dataInMem_hi_130;
  assign dataInMem_hi_130 = _GEN_196;
  wire [15:0]      dataInMem_lo_hi_198;
  assign dataInMem_lo_hi_198 = _GEN_196;
  wire [63:0]      dataInMem_lo_lo_lo_lo_lo_3 = {dataInMem_hi_68, dataInMem_lo_4, dataInMem_hi_67, dataInMem_lo_3};
  wire [63:0]      dataInMem_lo_lo_lo_lo_hi_3 = {dataInMem_hi_70, dataInMem_lo_6, dataInMem_hi_69, dataInMem_lo_5};
  wire [127:0]     dataInMem_lo_lo_lo_lo_3 = {dataInMem_lo_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_lo_lo_hi_lo_3 = {dataInMem_hi_72, dataInMem_lo_8, dataInMem_hi_71, dataInMem_lo_7};
  wire [63:0]      dataInMem_lo_lo_lo_hi_hi_3 = {dataInMem_hi_74, dataInMem_lo_10, dataInMem_hi_73, dataInMem_lo_9};
  wire [127:0]     dataInMem_lo_lo_lo_hi_3 = {dataInMem_lo_lo_lo_hi_hi_3, dataInMem_lo_lo_lo_hi_lo_3};
  wire [255:0]     dataInMem_lo_lo_lo_3 = {dataInMem_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_lo_hi_lo_lo_3 = {dataInMem_hi_76, dataInMem_lo_12, dataInMem_hi_75, dataInMem_lo_11};
  wire [63:0]      dataInMem_lo_lo_hi_lo_hi_3 = {dataInMem_hi_78, dataInMem_lo_14, dataInMem_hi_77, dataInMem_lo_13};
  wire [127:0]     dataInMem_lo_lo_hi_lo_3 = {dataInMem_lo_lo_hi_lo_hi_3, dataInMem_lo_lo_hi_lo_lo_3};
  wire [63:0]      dataInMem_lo_lo_hi_hi_lo_3 = {dataInMem_hi_80, dataInMem_lo_16, dataInMem_hi_79, dataInMem_lo_15};
  wire [63:0]      dataInMem_lo_lo_hi_hi_hi_3 = {dataInMem_hi_82, dataInMem_lo_18, dataInMem_hi_81, dataInMem_lo_17};
  wire [127:0]     dataInMem_lo_lo_hi_hi_3 = {dataInMem_lo_lo_hi_hi_hi_3, dataInMem_lo_lo_hi_hi_lo_3};
  wire [255:0]     dataInMem_lo_lo_hi_3 = {dataInMem_lo_lo_hi_hi_3, dataInMem_lo_lo_hi_lo_3};
  wire [511:0]     dataInMem_lo_lo_3 = {dataInMem_lo_lo_hi_3, dataInMem_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_lo_lo_lo_3 = {dataInMem_hi_84, dataInMem_lo_20, dataInMem_hi_83, dataInMem_lo_19};
  wire [63:0]      dataInMem_lo_hi_lo_lo_hi_3 = {dataInMem_hi_86, dataInMem_lo_22, dataInMem_hi_85, dataInMem_lo_21};
  wire [127:0]     dataInMem_lo_hi_lo_lo_3 = {dataInMem_lo_hi_lo_lo_hi_3, dataInMem_lo_hi_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_lo_hi_lo_3 = {dataInMem_hi_88, dataInMem_lo_24, dataInMem_hi_87, dataInMem_lo_23};
  wire [63:0]      dataInMem_lo_hi_lo_hi_hi_3 = {dataInMem_hi_90, dataInMem_lo_26, dataInMem_hi_89, dataInMem_lo_25};
  wire [127:0]     dataInMem_lo_hi_lo_hi_3 = {dataInMem_lo_hi_lo_hi_hi_3, dataInMem_lo_hi_lo_hi_lo_3};
  wire [255:0]     dataInMem_lo_hi_lo_3 = {dataInMem_lo_hi_lo_hi_3, dataInMem_lo_hi_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_hi_lo_lo_3 = {dataInMem_hi_92, dataInMem_lo_28, dataInMem_hi_91, dataInMem_lo_27};
  wire [63:0]      dataInMem_lo_hi_hi_lo_hi_3 = {dataInMem_hi_94, dataInMem_lo_30, dataInMem_hi_93, dataInMem_lo_29};
  wire [127:0]     dataInMem_lo_hi_hi_lo_3 = {dataInMem_lo_hi_hi_lo_hi_3, dataInMem_lo_hi_hi_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_hi_hi_lo_3 = {dataInMem_hi_96, dataInMem_lo_32, dataInMem_hi_95, dataInMem_lo_31};
  wire [63:0]      dataInMem_lo_hi_hi_hi_hi_3 = {dataInMem_hi_98, dataInMem_lo_34, dataInMem_hi_97, dataInMem_lo_33};
  wire [127:0]     dataInMem_lo_hi_hi_hi_3 = {dataInMem_lo_hi_hi_hi_hi_3, dataInMem_lo_hi_hi_hi_lo_3};
  wire [255:0]     dataInMem_lo_hi_hi_3 = {dataInMem_lo_hi_hi_hi_3, dataInMem_lo_hi_hi_lo_3};
  wire [511:0]     dataInMem_lo_hi_3 = {dataInMem_lo_hi_hi_3, dataInMem_lo_hi_lo_3};
  wire [1023:0]    dataInMem_lo_67 = {dataInMem_lo_hi_3, dataInMem_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_lo_lo_lo_3 = {dataInMem_hi_100, dataInMem_lo_36, dataInMem_hi_99, dataInMem_lo_35};
  wire [63:0]      dataInMem_hi_lo_lo_lo_hi_3 = {dataInMem_hi_102, dataInMem_lo_38, dataInMem_hi_101, dataInMem_lo_37};
  wire [127:0]     dataInMem_hi_lo_lo_lo_3 = {dataInMem_hi_lo_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_lo_hi_lo_3 = {dataInMem_hi_104, dataInMem_lo_40, dataInMem_hi_103, dataInMem_lo_39};
  wire [63:0]      dataInMem_hi_lo_lo_hi_hi_3 = {dataInMem_hi_106, dataInMem_lo_42, dataInMem_hi_105, dataInMem_lo_41};
  wire [127:0]     dataInMem_hi_lo_lo_hi_3 = {dataInMem_hi_lo_lo_hi_hi_3, dataInMem_hi_lo_lo_hi_lo_3};
  wire [255:0]     dataInMem_hi_lo_lo_3 = {dataInMem_hi_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_hi_lo_lo_3 = {dataInMem_hi_108, dataInMem_lo_44, dataInMem_hi_107, dataInMem_lo_43};
  wire [63:0]      dataInMem_hi_lo_hi_lo_hi_3 = {dataInMem_hi_110, dataInMem_lo_46, dataInMem_hi_109, dataInMem_lo_45};
  wire [127:0]     dataInMem_hi_lo_hi_lo_3 = {dataInMem_hi_lo_hi_lo_hi_3, dataInMem_hi_lo_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_hi_hi_lo_3 = {dataInMem_hi_112, dataInMem_lo_48, dataInMem_hi_111, dataInMem_lo_47};
  wire [63:0]      dataInMem_hi_lo_hi_hi_hi_3 = {dataInMem_hi_114, dataInMem_lo_50, dataInMem_hi_113, dataInMem_lo_49};
  wire [127:0]     dataInMem_hi_lo_hi_hi_3 = {dataInMem_hi_lo_hi_hi_hi_3, dataInMem_hi_lo_hi_hi_lo_3};
  wire [255:0]     dataInMem_hi_lo_hi_3 = {dataInMem_hi_lo_hi_hi_3, dataInMem_hi_lo_hi_lo_3};
  wire [511:0]     dataInMem_hi_lo_3 = {dataInMem_hi_lo_hi_3, dataInMem_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_lo_lo_lo_3 = {dataInMem_hi_116, dataInMem_lo_52, dataInMem_hi_115, dataInMem_lo_51};
  wire [63:0]      dataInMem_hi_hi_lo_lo_hi_3 = {dataInMem_hi_118, dataInMem_lo_54, dataInMem_hi_117, dataInMem_lo_53};
  wire [127:0]     dataInMem_hi_hi_lo_lo_3 = {dataInMem_hi_hi_lo_lo_hi_3, dataInMem_hi_hi_lo_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_lo_hi_lo_3 = {dataInMem_hi_120, dataInMem_lo_56, dataInMem_hi_119, dataInMem_lo_55};
  wire [63:0]      dataInMem_hi_hi_lo_hi_hi_3 = {dataInMem_hi_122, dataInMem_lo_58, dataInMem_hi_121, dataInMem_lo_57};
  wire [127:0]     dataInMem_hi_hi_lo_hi_3 = {dataInMem_hi_hi_lo_hi_hi_3, dataInMem_hi_hi_lo_hi_lo_3};
  wire [255:0]     dataInMem_hi_hi_lo_3 = {dataInMem_hi_hi_lo_hi_3, dataInMem_hi_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_hi_lo_lo_3 = {dataInMem_hi_124, dataInMem_lo_60, dataInMem_hi_123, dataInMem_lo_59};
  wire [63:0]      dataInMem_hi_hi_hi_lo_hi_3 = {dataInMem_hi_126, dataInMem_lo_62, dataInMem_hi_125, dataInMem_lo_61};
  wire [127:0]     dataInMem_hi_hi_hi_lo_3 = {dataInMem_hi_hi_hi_lo_hi_3, dataInMem_hi_hi_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_hi_hi_lo_3 = {dataInMem_hi_128, dataInMem_lo_64, dataInMem_hi_127, dataInMem_lo_63};
  wire [63:0]      dataInMem_hi_hi_hi_hi_hi_3 = {dataInMem_hi_130, dataInMem_lo_66, dataInMem_hi_129, dataInMem_lo_65};
  wire [127:0]     dataInMem_hi_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_hi_lo_3};
  wire [255:0]     dataInMem_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_lo_3};
  wire [511:0]     dataInMem_hi_hi_3 = {dataInMem_hi_hi_hi_3, dataInMem_hi_hi_lo_3};
  wire [1023:0]    dataInMem_hi_131 = {dataInMem_hi_hi_3, dataInMem_hi_lo_3};
  wire [2047:0]    dataInMem_3 = {dataInMem_hi_131, dataInMem_lo_67};
  wire [511:0]     regroupCacheLine_3_0 = dataInMem_3[511:0];
  wire [511:0]     regroupCacheLine_3_1 = dataInMem_3[1023:512];
  wire [511:0]     regroupCacheLine_3_2 = dataInMem_3[1535:1024];
  wire [511:0]     regroupCacheLine_3_3 = dataInMem_3[2047:1536];
  wire [511:0]     res_24 = regroupCacheLine_3_0;
  wire [511:0]     res_25 = regroupCacheLine_3_1;
  wire [511:0]     res_26 = regroupCacheLine_3_2;
  wire [511:0]     res_27 = regroupCacheLine_3_3;
  wire [1023:0]    lo_lo_3 = {res_25, res_24};
  wire [1023:0]    lo_hi_3 = {res_27, res_26};
  wire [2047:0]    lo_3 = {lo_hi_3, lo_lo_3};
  wire [4095:0]    regroupLoadData_0_3 = {2048'h0, lo_3};
  wire [15:0]      _GEN_197 = {dataRegroupBySew_4_0, dataRegroupBySew_3_0};
  wire [15:0]      dataInMem_hi_hi_4;
  assign dataInMem_hi_hi_4 = _GEN_197;
  wire [15:0]      dataInMem_hi_lo_6;
  assign dataInMem_hi_lo_6 = _GEN_197;
  wire [23:0]      dataInMem_hi_132 = {dataInMem_hi_hi_4, dataRegroupBySew_2_0};
  wire [15:0]      _GEN_198 = {dataRegroupBySew_4_1, dataRegroupBySew_3_1};
  wire [15:0]      dataInMem_hi_hi_5;
  assign dataInMem_hi_hi_5 = _GEN_198;
  wire [15:0]      dataInMem_hi_lo_7;
  assign dataInMem_hi_lo_7 = _GEN_198;
  wire [23:0]      dataInMem_hi_133 = {dataInMem_hi_hi_5, dataRegroupBySew_2_1};
  wire [15:0]      _GEN_199 = {dataRegroupBySew_4_2, dataRegroupBySew_3_2};
  wire [15:0]      dataInMem_hi_hi_6;
  assign dataInMem_hi_hi_6 = _GEN_199;
  wire [15:0]      dataInMem_hi_lo_8;
  assign dataInMem_hi_lo_8 = _GEN_199;
  wire [23:0]      dataInMem_hi_134 = {dataInMem_hi_hi_6, dataRegroupBySew_2_2};
  wire [15:0]      _GEN_200 = {dataRegroupBySew_4_3, dataRegroupBySew_3_3};
  wire [15:0]      dataInMem_hi_hi_7;
  assign dataInMem_hi_hi_7 = _GEN_200;
  wire [15:0]      dataInMem_hi_lo_9;
  assign dataInMem_hi_lo_9 = _GEN_200;
  wire [23:0]      dataInMem_hi_135 = {dataInMem_hi_hi_7, dataRegroupBySew_2_3};
  wire [15:0]      _GEN_201 = {dataRegroupBySew_4_4, dataRegroupBySew_3_4};
  wire [15:0]      dataInMem_hi_hi_8;
  assign dataInMem_hi_hi_8 = _GEN_201;
  wire [15:0]      dataInMem_hi_lo_10;
  assign dataInMem_hi_lo_10 = _GEN_201;
  wire [23:0]      dataInMem_hi_136 = {dataInMem_hi_hi_8, dataRegroupBySew_2_4};
  wire [15:0]      _GEN_202 = {dataRegroupBySew_4_5, dataRegroupBySew_3_5};
  wire [15:0]      dataInMem_hi_hi_9;
  assign dataInMem_hi_hi_9 = _GEN_202;
  wire [15:0]      dataInMem_hi_lo_11;
  assign dataInMem_hi_lo_11 = _GEN_202;
  wire [23:0]      dataInMem_hi_137 = {dataInMem_hi_hi_9, dataRegroupBySew_2_5};
  wire [15:0]      _GEN_203 = {dataRegroupBySew_4_6, dataRegroupBySew_3_6};
  wire [15:0]      dataInMem_hi_hi_10;
  assign dataInMem_hi_hi_10 = _GEN_203;
  wire [15:0]      dataInMem_hi_lo_12;
  assign dataInMem_hi_lo_12 = _GEN_203;
  wire [23:0]      dataInMem_hi_138 = {dataInMem_hi_hi_10, dataRegroupBySew_2_6};
  wire [15:0]      _GEN_204 = {dataRegroupBySew_4_7, dataRegroupBySew_3_7};
  wire [15:0]      dataInMem_hi_hi_11;
  assign dataInMem_hi_hi_11 = _GEN_204;
  wire [15:0]      dataInMem_hi_lo_13;
  assign dataInMem_hi_lo_13 = _GEN_204;
  wire [23:0]      dataInMem_hi_139 = {dataInMem_hi_hi_11, dataRegroupBySew_2_7};
  wire [15:0]      _GEN_205 = {dataRegroupBySew_4_8, dataRegroupBySew_3_8};
  wire [15:0]      dataInMem_hi_hi_12;
  assign dataInMem_hi_hi_12 = _GEN_205;
  wire [15:0]      dataInMem_hi_lo_14;
  assign dataInMem_hi_lo_14 = _GEN_205;
  wire [23:0]      dataInMem_hi_140 = {dataInMem_hi_hi_12, dataRegroupBySew_2_8};
  wire [15:0]      _GEN_206 = {dataRegroupBySew_4_9, dataRegroupBySew_3_9};
  wire [15:0]      dataInMem_hi_hi_13;
  assign dataInMem_hi_hi_13 = _GEN_206;
  wire [15:0]      dataInMem_hi_lo_15;
  assign dataInMem_hi_lo_15 = _GEN_206;
  wire [23:0]      dataInMem_hi_141 = {dataInMem_hi_hi_13, dataRegroupBySew_2_9};
  wire [15:0]      _GEN_207 = {dataRegroupBySew_4_10, dataRegroupBySew_3_10};
  wire [15:0]      dataInMem_hi_hi_14;
  assign dataInMem_hi_hi_14 = _GEN_207;
  wire [15:0]      dataInMem_hi_lo_16;
  assign dataInMem_hi_lo_16 = _GEN_207;
  wire [23:0]      dataInMem_hi_142 = {dataInMem_hi_hi_14, dataRegroupBySew_2_10};
  wire [15:0]      _GEN_208 = {dataRegroupBySew_4_11, dataRegroupBySew_3_11};
  wire [15:0]      dataInMem_hi_hi_15;
  assign dataInMem_hi_hi_15 = _GEN_208;
  wire [15:0]      dataInMem_hi_lo_17;
  assign dataInMem_hi_lo_17 = _GEN_208;
  wire [23:0]      dataInMem_hi_143 = {dataInMem_hi_hi_15, dataRegroupBySew_2_11};
  wire [15:0]      _GEN_209 = {dataRegroupBySew_4_12, dataRegroupBySew_3_12};
  wire [15:0]      dataInMem_hi_hi_16;
  assign dataInMem_hi_hi_16 = _GEN_209;
  wire [15:0]      dataInMem_hi_lo_18;
  assign dataInMem_hi_lo_18 = _GEN_209;
  wire [23:0]      dataInMem_hi_144 = {dataInMem_hi_hi_16, dataRegroupBySew_2_12};
  wire [15:0]      _GEN_210 = {dataRegroupBySew_4_13, dataRegroupBySew_3_13};
  wire [15:0]      dataInMem_hi_hi_17;
  assign dataInMem_hi_hi_17 = _GEN_210;
  wire [15:0]      dataInMem_hi_lo_19;
  assign dataInMem_hi_lo_19 = _GEN_210;
  wire [23:0]      dataInMem_hi_145 = {dataInMem_hi_hi_17, dataRegroupBySew_2_13};
  wire [15:0]      _GEN_211 = {dataRegroupBySew_4_14, dataRegroupBySew_3_14};
  wire [15:0]      dataInMem_hi_hi_18;
  assign dataInMem_hi_hi_18 = _GEN_211;
  wire [15:0]      dataInMem_hi_lo_20;
  assign dataInMem_hi_lo_20 = _GEN_211;
  wire [23:0]      dataInMem_hi_146 = {dataInMem_hi_hi_18, dataRegroupBySew_2_14};
  wire [15:0]      _GEN_212 = {dataRegroupBySew_4_15, dataRegroupBySew_3_15};
  wire [15:0]      dataInMem_hi_hi_19;
  assign dataInMem_hi_hi_19 = _GEN_212;
  wire [15:0]      dataInMem_hi_lo_21;
  assign dataInMem_hi_lo_21 = _GEN_212;
  wire [23:0]      dataInMem_hi_147 = {dataInMem_hi_hi_19, dataRegroupBySew_2_15};
  wire [15:0]      _GEN_213 = {dataRegroupBySew_4_16, dataRegroupBySew_3_16};
  wire [15:0]      dataInMem_hi_hi_20;
  assign dataInMem_hi_hi_20 = _GEN_213;
  wire [15:0]      dataInMem_hi_lo_22;
  assign dataInMem_hi_lo_22 = _GEN_213;
  wire [23:0]      dataInMem_hi_148 = {dataInMem_hi_hi_20, dataRegroupBySew_2_16};
  wire [15:0]      _GEN_214 = {dataRegroupBySew_4_17, dataRegroupBySew_3_17};
  wire [15:0]      dataInMem_hi_hi_21;
  assign dataInMem_hi_hi_21 = _GEN_214;
  wire [15:0]      dataInMem_hi_lo_23;
  assign dataInMem_hi_lo_23 = _GEN_214;
  wire [23:0]      dataInMem_hi_149 = {dataInMem_hi_hi_21, dataRegroupBySew_2_17};
  wire [15:0]      _GEN_215 = {dataRegroupBySew_4_18, dataRegroupBySew_3_18};
  wire [15:0]      dataInMem_hi_hi_22;
  assign dataInMem_hi_hi_22 = _GEN_215;
  wire [15:0]      dataInMem_hi_lo_24;
  assign dataInMem_hi_lo_24 = _GEN_215;
  wire [23:0]      dataInMem_hi_150 = {dataInMem_hi_hi_22, dataRegroupBySew_2_18};
  wire [15:0]      _GEN_216 = {dataRegroupBySew_4_19, dataRegroupBySew_3_19};
  wire [15:0]      dataInMem_hi_hi_23;
  assign dataInMem_hi_hi_23 = _GEN_216;
  wire [15:0]      dataInMem_hi_lo_25;
  assign dataInMem_hi_lo_25 = _GEN_216;
  wire [23:0]      dataInMem_hi_151 = {dataInMem_hi_hi_23, dataRegroupBySew_2_19};
  wire [15:0]      _GEN_217 = {dataRegroupBySew_4_20, dataRegroupBySew_3_20};
  wire [15:0]      dataInMem_hi_hi_24;
  assign dataInMem_hi_hi_24 = _GEN_217;
  wire [15:0]      dataInMem_hi_lo_26;
  assign dataInMem_hi_lo_26 = _GEN_217;
  wire [23:0]      dataInMem_hi_152 = {dataInMem_hi_hi_24, dataRegroupBySew_2_20};
  wire [15:0]      _GEN_218 = {dataRegroupBySew_4_21, dataRegroupBySew_3_21};
  wire [15:0]      dataInMem_hi_hi_25;
  assign dataInMem_hi_hi_25 = _GEN_218;
  wire [15:0]      dataInMem_hi_lo_27;
  assign dataInMem_hi_lo_27 = _GEN_218;
  wire [23:0]      dataInMem_hi_153 = {dataInMem_hi_hi_25, dataRegroupBySew_2_21};
  wire [15:0]      _GEN_219 = {dataRegroupBySew_4_22, dataRegroupBySew_3_22};
  wire [15:0]      dataInMem_hi_hi_26;
  assign dataInMem_hi_hi_26 = _GEN_219;
  wire [15:0]      dataInMem_hi_lo_28;
  assign dataInMem_hi_lo_28 = _GEN_219;
  wire [23:0]      dataInMem_hi_154 = {dataInMem_hi_hi_26, dataRegroupBySew_2_22};
  wire [15:0]      _GEN_220 = {dataRegroupBySew_4_23, dataRegroupBySew_3_23};
  wire [15:0]      dataInMem_hi_hi_27;
  assign dataInMem_hi_hi_27 = _GEN_220;
  wire [15:0]      dataInMem_hi_lo_29;
  assign dataInMem_hi_lo_29 = _GEN_220;
  wire [23:0]      dataInMem_hi_155 = {dataInMem_hi_hi_27, dataRegroupBySew_2_23};
  wire [15:0]      _GEN_221 = {dataRegroupBySew_4_24, dataRegroupBySew_3_24};
  wire [15:0]      dataInMem_hi_hi_28;
  assign dataInMem_hi_hi_28 = _GEN_221;
  wire [15:0]      dataInMem_hi_lo_30;
  assign dataInMem_hi_lo_30 = _GEN_221;
  wire [23:0]      dataInMem_hi_156 = {dataInMem_hi_hi_28, dataRegroupBySew_2_24};
  wire [15:0]      _GEN_222 = {dataRegroupBySew_4_25, dataRegroupBySew_3_25};
  wire [15:0]      dataInMem_hi_hi_29;
  assign dataInMem_hi_hi_29 = _GEN_222;
  wire [15:0]      dataInMem_hi_lo_31;
  assign dataInMem_hi_lo_31 = _GEN_222;
  wire [23:0]      dataInMem_hi_157 = {dataInMem_hi_hi_29, dataRegroupBySew_2_25};
  wire [15:0]      _GEN_223 = {dataRegroupBySew_4_26, dataRegroupBySew_3_26};
  wire [15:0]      dataInMem_hi_hi_30;
  assign dataInMem_hi_hi_30 = _GEN_223;
  wire [15:0]      dataInMem_hi_lo_32;
  assign dataInMem_hi_lo_32 = _GEN_223;
  wire [23:0]      dataInMem_hi_158 = {dataInMem_hi_hi_30, dataRegroupBySew_2_26};
  wire [15:0]      _GEN_224 = {dataRegroupBySew_4_27, dataRegroupBySew_3_27};
  wire [15:0]      dataInMem_hi_hi_31;
  assign dataInMem_hi_hi_31 = _GEN_224;
  wire [15:0]      dataInMem_hi_lo_33;
  assign dataInMem_hi_lo_33 = _GEN_224;
  wire [23:0]      dataInMem_hi_159 = {dataInMem_hi_hi_31, dataRegroupBySew_2_27};
  wire [15:0]      _GEN_225 = {dataRegroupBySew_4_28, dataRegroupBySew_3_28};
  wire [15:0]      dataInMem_hi_hi_32;
  assign dataInMem_hi_hi_32 = _GEN_225;
  wire [15:0]      dataInMem_hi_lo_34;
  assign dataInMem_hi_lo_34 = _GEN_225;
  wire [23:0]      dataInMem_hi_160 = {dataInMem_hi_hi_32, dataRegroupBySew_2_28};
  wire [15:0]      _GEN_226 = {dataRegroupBySew_4_29, dataRegroupBySew_3_29};
  wire [15:0]      dataInMem_hi_hi_33;
  assign dataInMem_hi_hi_33 = _GEN_226;
  wire [15:0]      dataInMem_hi_lo_35;
  assign dataInMem_hi_lo_35 = _GEN_226;
  wire [23:0]      dataInMem_hi_161 = {dataInMem_hi_hi_33, dataRegroupBySew_2_29};
  wire [15:0]      _GEN_227 = {dataRegroupBySew_4_30, dataRegroupBySew_3_30};
  wire [15:0]      dataInMem_hi_hi_34;
  assign dataInMem_hi_hi_34 = _GEN_227;
  wire [15:0]      dataInMem_hi_lo_36;
  assign dataInMem_hi_lo_36 = _GEN_227;
  wire [23:0]      dataInMem_hi_162 = {dataInMem_hi_hi_34, dataRegroupBySew_2_30};
  wire [15:0]      _GEN_228 = {dataRegroupBySew_4_31, dataRegroupBySew_3_31};
  wire [15:0]      dataInMem_hi_hi_35;
  assign dataInMem_hi_hi_35 = _GEN_228;
  wire [15:0]      dataInMem_hi_lo_37;
  assign dataInMem_hi_lo_37 = _GEN_228;
  wire [23:0]      dataInMem_hi_163 = {dataInMem_hi_hi_35, dataRegroupBySew_2_31};
  wire [15:0]      _GEN_229 = {dataRegroupBySew_4_32, dataRegroupBySew_3_32};
  wire [15:0]      dataInMem_hi_hi_36;
  assign dataInMem_hi_hi_36 = _GEN_229;
  wire [15:0]      dataInMem_hi_lo_38;
  assign dataInMem_hi_lo_38 = _GEN_229;
  wire [23:0]      dataInMem_hi_164 = {dataInMem_hi_hi_36, dataRegroupBySew_2_32};
  wire [15:0]      _GEN_230 = {dataRegroupBySew_4_33, dataRegroupBySew_3_33};
  wire [15:0]      dataInMem_hi_hi_37;
  assign dataInMem_hi_hi_37 = _GEN_230;
  wire [15:0]      dataInMem_hi_lo_39;
  assign dataInMem_hi_lo_39 = _GEN_230;
  wire [23:0]      dataInMem_hi_165 = {dataInMem_hi_hi_37, dataRegroupBySew_2_33};
  wire [15:0]      _GEN_231 = {dataRegroupBySew_4_34, dataRegroupBySew_3_34};
  wire [15:0]      dataInMem_hi_hi_38;
  assign dataInMem_hi_hi_38 = _GEN_231;
  wire [15:0]      dataInMem_hi_lo_40;
  assign dataInMem_hi_lo_40 = _GEN_231;
  wire [23:0]      dataInMem_hi_166 = {dataInMem_hi_hi_38, dataRegroupBySew_2_34};
  wire [15:0]      _GEN_232 = {dataRegroupBySew_4_35, dataRegroupBySew_3_35};
  wire [15:0]      dataInMem_hi_hi_39;
  assign dataInMem_hi_hi_39 = _GEN_232;
  wire [15:0]      dataInMem_hi_lo_41;
  assign dataInMem_hi_lo_41 = _GEN_232;
  wire [23:0]      dataInMem_hi_167 = {dataInMem_hi_hi_39, dataRegroupBySew_2_35};
  wire [15:0]      _GEN_233 = {dataRegroupBySew_4_36, dataRegroupBySew_3_36};
  wire [15:0]      dataInMem_hi_hi_40;
  assign dataInMem_hi_hi_40 = _GEN_233;
  wire [15:0]      dataInMem_hi_lo_42;
  assign dataInMem_hi_lo_42 = _GEN_233;
  wire [23:0]      dataInMem_hi_168 = {dataInMem_hi_hi_40, dataRegroupBySew_2_36};
  wire [15:0]      _GEN_234 = {dataRegroupBySew_4_37, dataRegroupBySew_3_37};
  wire [15:0]      dataInMem_hi_hi_41;
  assign dataInMem_hi_hi_41 = _GEN_234;
  wire [15:0]      dataInMem_hi_lo_43;
  assign dataInMem_hi_lo_43 = _GEN_234;
  wire [23:0]      dataInMem_hi_169 = {dataInMem_hi_hi_41, dataRegroupBySew_2_37};
  wire [15:0]      _GEN_235 = {dataRegroupBySew_4_38, dataRegroupBySew_3_38};
  wire [15:0]      dataInMem_hi_hi_42;
  assign dataInMem_hi_hi_42 = _GEN_235;
  wire [15:0]      dataInMem_hi_lo_44;
  assign dataInMem_hi_lo_44 = _GEN_235;
  wire [23:0]      dataInMem_hi_170 = {dataInMem_hi_hi_42, dataRegroupBySew_2_38};
  wire [15:0]      _GEN_236 = {dataRegroupBySew_4_39, dataRegroupBySew_3_39};
  wire [15:0]      dataInMem_hi_hi_43;
  assign dataInMem_hi_hi_43 = _GEN_236;
  wire [15:0]      dataInMem_hi_lo_45;
  assign dataInMem_hi_lo_45 = _GEN_236;
  wire [23:0]      dataInMem_hi_171 = {dataInMem_hi_hi_43, dataRegroupBySew_2_39};
  wire [15:0]      _GEN_237 = {dataRegroupBySew_4_40, dataRegroupBySew_3_40};
  wire [15:0]      dataInMem_hi_hi_44;
  assign dataInMem_hi_hi_44 = _GEN_237;
  wire [15:0]      dataInMem_hi_lo_46;
  assign dataInMem_hi_lo_46 = _GEN_237;
  wire [23:0]      dataInMem_hi_172 = {dataInMem_hi_hi_44, dataRegroupBySew_2_40};
  wire [15:0]      _GEN_238 = {dataRegroupBySew_4_41, dataRegroupBySew_3_41};
  wire [15:0]      dataInMem_hi_hi_45;
  assign dataInMem_hi_hi_45 = _GEN_238;
  wire [15:0]      dataInMem_hi_lo_47;
  assign dataInMem_hi_lo_47 = _GEN_238;
  wire [23:0]      dataInMem_hi_173 = {dataInMem_hi_hi_45, dataRegroupBySew_2_41};
  wire [15:0]      _GEN_239 = {dataRegroupBySew_4_42, dataRegroupBySew_3_42};
  wire [15:0]      dataInMem_hi_hi_46;
  assign dataInMem_hi_hi_46 = _GEN_239;
  wire [15:0]      dataInMem_hi_lo_48;
  assign dataInMem_hi_lo_48 = _GEN_239;
  wire [23:0]      dataInMem_hi_174 = {dataInMem_hi_hi_46, dataRegroupBySew_2_42};
  wire [15:0]      _GEN_240 = {dataRegroupBySew_4_43, dataRegroupBySew_3_43};
  wire [15:0]      dataInMem_hi_hi_47;
  assign dataInMem_hi_hi_47 = _GEN_240;
  wire [15:0]      dataInMem_hi_lo_49;
  assign dataInMem_hi_lo_49 = _GEN_240;
  wire [23:0]      dataInMem_hi_175 = {dataInMem_hi_hi_47, dataRegroupBySew_2_43};
  wire [15:0]      _GEN_241 = {dataRegroupBySew_4_44, dataRegroupBySew_3_44};
  wire [15:0]      dataInMem_hi_hi_48;
  assign dataInMem_hi_hi_48 = _GEN_241;
  wire [15:0]      dataInMem_hi_lo_50;
  assign dataInMem_hi_lo_50 = _GEN_241;
  wire [23:0]      dataInMem_hi_176 = {dataInMem_hi_hi_48, dataRegroupBySew_2_44};
  wire [15:0]      _GEN_242 = {dataRegroupBySew_4_45, dataRegroupBySew_3_45};
  wire [15:0]      dataInMem_hi_hi_49;
  assign dataInMem_hi_hi_49 = _GEN_242;
  wire [15:0]      dataInMem_hi_lo_51;
  assign dataInMem_hi_lo_51 = _GEN_242;
  wire [23:0]      dataInMem_hi_177 = {dataInMem_hi_hi_49, dataRegroupBySew_2_45};
  wire [15:0]      _GEN_243 = {dataRegroupBySew_4_46, dataRegroupBySew_3_46};
  wire [15:0]      dataInMem_hi_hi_50;
  assign dataInMem_hi_hi_50 = _GEN_243;
  wire [15:0]      dataInMem_hi_lo_52;
  assign dataInMem_hi_lo_52 = _GEN_243;
  wire [23:0]      dataInMem_hi_178 = {dataInMem_hi_hi_50, dataRegroupBySew_2_46};
  wire [15:0]      _GEN_244 = {dataRegroupBySew_4_47, dataRegroupBySew_3_47};
  wire [15:0]      dataInMem_hi_hi_51;
  assign dataInMem_hi_hi_51 = _GEN_244;
  wire [15:0]      dataInMem_hi_lo_53;
  assign dataInMem_hi_lo_53 = _GEN_244;
  wire [23:0]      dataInMem_hi_179 = {dataInMem_hi_hi_51, dataRegroupBySew_2_47};
  wire [15:0]      _GEN_245 = {dataRegroupBySew_4_48, dataRegroupBySew_3_48};
  wire [15:0]      dataInMem_hi_hi_52;
  assign dataInMem_hi_hi_52 = _GEN_245;
  wire [15:0]      dataInMem_hi_lo_54;
  assign dataInMem_hi_lo_54 = _GEN_245;
  wire [23:0]      dataInMem_hi_180 = {dataInMem_hi_hi_52, dataRegroupBySew_2_48};
  wire [15:0]      _GEN_246 = {dataRegroupBySew_4_49, dataRegroupBySew_3_49};
  wire [15:0]      dataInMem_hi_hi_53;
  assign dataInMem_hi_hi_53 = _GEN_246;
  wire [15:0]      dataInMem_hi_lo_55;
  assign dataInMem_hi_lo_55 = _GEN_246;
  wire [23:0]      dataInMem_hi_181 = {dataInMem_hi_hi_53, dataRegroupBySew_2_49};
  wire [15:0]      _GEN_247 = {dataRegroupBySew_4_50, dataRegroupBySew_3_50};
  wire [15:0]      dataInMem_hi_hi_54;
  assign dataInMem_hi_hi_54 = _GEN_247;
  wire [15:0]      dataInMem_hi_lo_56;
  assign dataInMem_hi_lo_56 = _GEN_247;
  wire [23:0]      dataInMem_hi_182 = {dataInMem_hi_hi_54, dataRegroupBySew_2_50};
  wire [15:0]      _GEN_248 = {dataRegroupBySew_4_51, dataRegroupBySew_3_51};
  wire [15:0]      dataInMem_hi_hi_55;
  assign dataInMem_hi_hi_55 = _GEN_248;
  wire [15:0]      dataInMem_hi_lo_57;
  assign dataInMem_hi_lo_57 = _GEN_248;
  wire [23:0]      dataInMem_hi_183 = {dataInMem_hi_hi_55, dataRegroupBySew_2_51};
  wire [15:0]      _GEN_249 = {dataRegroupBySew_4_52, dataRegroupBySew_3_52};
  wire [15:0]      dataInMem_hi_hi_56;
  assign dataInMem_hi_hi_56 = _GEN_249;
  wire [15:0]      dataInMem_hi_lo_58;
  assign dataInMem_hi_lo_58 = _GEN_249;
  wire [23:0]      dataInMem_hi_184 = {dataInMem_hi_hi_56, dataRegroupBySew_2_52};
  wire [15:0]      _GEN_250 = {dataRegroupBySew_4_53, dataRegroupBySew_3_53};
  wire [15:0]      dataInMem_hi_hi_57;
  assign dataInMem_hi_hi_57 = _GEN_250;
  wire [15:0]      dataInMem_hi_lo_59;
  assign dataInMem_hi_lo_59 = _GEN_250;
  wire [23:0]      dataInMem_hi_185 = {dataInMem_hi_hi_57, dataRegroupBySew_2_53};
  wire [15:0]      _GEN_251 = {dataRegroupBySew_4_54, dataRegroupBySew_3_54};
  wire [15:0]      dataInMem_hi_hi_58;
  assign dataInMem_hi_hi_58 = _GEN_251;
  wire [15:0]      dataInMem_hi_lo_60;
  assign dataInMem_hi_lo_60 = _GEN_251;
  wire [23:0]      dataInMem_hi_186 = {dataInMem_hi_hi_58, dataRegroupBySew_2_54};
  wire [15:0]      _GEN_252 = {dataRegroupBySew_4_55, dataRegroupBySew_3_55};
  wire [15:0]      dataInMem_hi_hi_59;
  assign dataInMem_hi_hi_59 = _GEN_252;
  wire [15:0]      dataInMem_hi_lo_61;
  assign dataInMem_hi_lo_61 = _GEN_252;
  wire [23:0]      dataInMem_hi_187 = {dataInMem_hi_hi_59, dataRegroupBySew_2_55};
  wire [15:0]      _GEN_253 = {dataRegroupBySew_4_56, dataRegroupBySew_3_56};
  wire [15:0]      dataInMem_hi_hi_60;
  assign dataInMem_hi_hi_60 = _GEN_253;
  wire [15:0]      dataInMem_hi_lo_62;
  assign dataInMem_hi_lo_62 = _GEN_253;
  wire [23:0]      dataInMem_hi_188 = {dataInMem_hi_hi_60, dataRegroupBySew_2_56};
  wire [15:0]      _GEN_254 = {dataRegroupBySew_4_57, dataRegroupBySew_3_57};
  wire [15:0]      dataInMem_hi_hi_61;
  assign dataInMem_hi_hi_61 = _GEN_254;
  wire [15:0]      dataInMem_hi_lo_63;
  assign dataInMem_hi_lo_63 = _GEN_254;
  wire [23:0]      dataInMem_hi_189 = {dataInMem_hi_hi_61, dataRegroupBySew_2_57};
  wire [15:0]      _GEN_255 = {dataRegroupBySew_4_58, dataRegroupBySew_3_58};
  wire [15:0]      dataInMem_hi_hi_62;
  assign dataInMem_hi_hi_62 = _GEN_255;
  wire [15:0]      dataInMem_hi_lo_64;
  assign dataInMem_hi_lo_64 = _GEN_255;
  wire [23:0]      dataInMem_hi_190 = {dataInMem_hi_hi_62, dataRegroupBySew_2_58};
  wire [15:0]      _GEN_256 = {dataRegroupBySew_4_59, dataRegroupBySew_3_59};
  wire [15:0]      dataInMem_hi_hi_63;
  assign dataInMem_hi_hi_63 = _GEN_256;
  wire [15:0]      dataInMem_hi_lo_65;
  assign dataInMem_hi_lo_65 = _GEN_256;
  wire [23:0]      dataInMem_hi_191 = {dataInMem_hi_hi_63, dataRegroupBySew_2_59};
  wire [15:0]      _GEN_257 = {dataRegroupBySew_4_60, dataRegroupBySew_3_60};
  wire [15:0]      dataInMem_hi_hi_64;
  assign dataInMem_hi_hi_64 = _GEN_257;
  wire [15:0]      dataInMem_hi_lo_66;
  assign dataInMem_hi_lo_66 = _GEN_257;
  wire [23:0]      dataInMem_hi_192 = {dataInMem_hi_hi_64, dataRegroupBySew_2_60};
  wire [15:0]      _GEN_258 = {dataRegroupBySew_4_61, dataRegroupBySew_3_61};
  wire [15:0]      dataInMem_hi_hi_65;
  assign dataInMem_hi_hi_65 = _GEN_258;
  wire [15:0]      dataInMem_hi_lo_67;
  assign dataInMem_hi_lo_67 = _GEN_258;
  wire [23:0]      dataInMem_hi_193 = {dataInMem_hi_hi_65, dataRegroupBySew_2_61};
  wire [15:0]      _GEN_259 = {dataRegroupBySew_4_62, dataRegroupBySew_3_62};
  wire [15:0]      dataInMem_hi_hi_66;
  assign dataInMem_hi_hi_66 = _GEN_259;
  wire [15:0]      dataInMem_hi_lo_68;
  assign dataInMem_hi_lo_68 = _GEN_259;
  wire [23:0]      dataInMem_hi_194 = {dataInMem_hi_hi_66, dataRegroupBySew_2_62};
  wire [15:0]      _GEN_260 = {dataRegroupBySew_4_63, dataRegroupBySew_3_63};
  wire [15:0]      dataInMem_hi_hi_67;
  assign dataInMem_hi_hi_67 = _GEN_260;
  wire [15:0]      dataInMem_hi_lo_69;
  assign dataInMem_hi_lo_69 = _GEN_260;
  wire [23:0]      dataInMem_hi_195 = {dataInMem_hi_hi_67, dataRegroupBySew_2_63};
  wire [79:0]      dataInMem_lo_lo_lo_lo_lo_4 = {dataInMem_hi_133, dataInMem_lo_69, dataInMem_hi_132, dataInMem_lo_68};
  wire [79:0]      dataInMem_lo_lo_lo_lo_hi_4 = {dataInMem_hi_135, dataInMem_lo_71, dataInMem_hi_134, dataInMem_lo_70};
  wire [159:0]     dataInMem_lo_lo_lo_lo_4 = {dataInMem_lo_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_lo_lo_hi_lo_4 = {dataInMem_hi_137, dataInMem_lo_73, dataInMem_hi_136, dataInMem_lo_72};
  wire [79:0]      dataInMem_lo_lo_lo_hi_hi_4 = {dataInMem_hi_139, dataInMem_lo_75, dataInMem_hi_138, dataInMem_lo_74};
  wire [159:0]     dataInMem_lo_lo_lo_hi_4 = {dataInMem_lo_lo_lo_hi_hi_4, dataInMem_lo_lo_lo_hi_lo_4};
  wire [319:0]     dataInMem_lo_lo_lo_4 = {dataInMem_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_lo_hi_lo_lo_4 = {dataInMem_hi_141, dataInMem_lo_77, dataInMem_hi_140, dataInMem_lo_76};
  wire [79:0]      dataInMem_lo_lo_hi_lo_hi_4 = {dataInMem_hi_143, dataInMem_lo_79, dataInMem_hi_142, dataInMem_lo_78};
  wire [159:0]     dataInMem_lo_lo_hi_lo_4 = {dataInMem_lo_lo_hi_lo_hi_4, dataInMem_lo_lo_hi_lo_lo_4};
  wire [79:0]      dataInMem_lo_lo_hi_hi_lo_4 = {dataInMem_hi_145, dataInMem_lo_81, dataInMem_hi_144, dataInMem_lo_80};
  wire [79:0]      dataInMem_lo_lo_hi_hi_hi_4 = {dataInMem_hi_147, dataInMem_lo_83, dataInMem_hi_146, dataInMem_lo_82};
  wire [159:0]     dataInMem_lo_lo_hi_hi_4 = {dataInMem_lo_lo_hi_hi_hi_4, dataInMem_lo_lo_hi_hi_lo_4};
  wire [319:0]     dataInMem_lo_lo_hi_4 = {dataInMem_lo_lo_hi_hi_4, dataInMem_lo_lo_hi_lo_4};
  wire [639:0]     dataInMem_lo_lo_4 = {dataInMem_lo_lo_hi_4, dataInMem_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_lo_lo_lo_4 = {dataInMem_hi_149, dataInMem_lo_85, dataInMem_hi_148, dataInMem_lo_84};
  wire [79:0]      dataInMem_lo_hi_lo_lo_hi_4 = {dataInMem_hi_151, dataInMem_lo_87, dataInMem_hi_150, dataInMem_lo_86};
  wire [159:0]     dataInMem_lo_hi_lo_lo_4 = {dataInMem_lo_hi_lo_lo_hi_4, dataInMem_lo_hi_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_lo_hi_lo_4 = {dataInMem_hi_153, dataInMem_lo_89, dataInMem_hi_152, dataInMem_lo_88};
  wire [79:0]      dataInMem_lo_hi_lo_hi_hi_4 = {dataInMem_hi_155, dataInMem_lo_91, dataInMem_hi_154, dataInMem_lo_90};
  wire [159:0]     dataInMem_lo_hi_lo_hi_4 = {dataInMem_lo_hi_lo_hi_hi_4, dataInMem_lo_hi_lo_hi_lo_4};
  wire [319:0]     dataInMem_lo_hi_lo_4 = {dataInMem_lo_hi_lo_hi_4, dataInMem_lo_hi_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_hi_lo_lo_4 = {dataInMem_hi_157, dataInMem_lo_93, dataInMem_hi_156, dataInMem_lo_92};
  wire [79:0]      dataInMem_lo_hi_hi_lo_hi_4 = {dataInMem_hi_159, dataInMem_lo_95, dataInMem_hi_158, dataInMem_lo_94};
  wire [159:0]     dataInMem_lo_hi_hi_lo_4 = {dataInMem_lo_hi_hi_lo_hi_4, dataInMem_lo_hi_hi_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_hi_hi_lo_4 = {dataInMem_hi_161, dataInMem_lo_97, dataInMem_hi_160, dataInMem_lo_96};
  wire [79:0]      dataInMem_lo_hi_hi_hi_hi_4 = {dataInMem_hi_163, dataInMem_lo_99, dataInMem_hi_162, dataInMem_lo_98};
  wire [159:0]     dataInMem_lo_hi_hi_hi_4 = {dataInMem_lo_hi_hi_hi_hi_4, dataInMem_lo_hi_hi_hi_lo_4};
  wire [319:0]     dataInMem_lo_hi_hi_4 = {dataInMem_lo_hi_hi_hi_4, dataInMem_lo_hi_hi_lo_4};
  wire [639:0]     dataInMem_lo_hi_4 = {dataInMem_lo_hi_hi_4, dataInMem_lo_hi_lo_4};
  wire [1279:0]    dataInMem_lo_132 = {dataInMem_lo_hi_4, dataInMem_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_lo_lo_lo_4 = {dataInMem_hi_165, dataInMem_lo_101, dataInMem_hi_164, dataInMem_lo_100};
  wire [79:0]      dataInMem_hi_lo_lo_lo_hi_4 = {dataInMem_hi_167, dataInMem_lo_103, dataInMem_hi_166, dataInMem_lo_102};
  wire [159:0]     dataInMem_hi_lo_lo_lo_4 = {dataInMem_hi_lo_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_lo_hi_lo_4 = {dataInMem_hi_169, dataInMem_lo_105, dataInMem_hi_168, dataInMem_lo_104};
  wire [79:0]      dataInMem_hi_lo_lo_hi_hi_4 = {dataInMem_hi_171, dataInMem_lo_107, dataInMem_hi_170, dataInMem_lo_106};
  wire [159:0]     dataInMem_hi_lo_lo_hi_4 = {dataInMem_hi_lo_lo_hi_hi_4, dataInMem_hi_lo_lo_hi_lo_4};
  wire [319:0]     dataInMem_hi_lo_lo_4 = {dataInMem_hi_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_hi_lo_lo_4 = {dataInMem_hi_173, dataInMem_lo_109, dataInMem_hi_172, dataInMem_lo_108};
  wire [79:0]      dataInMem_hi_lo_hi_lo_hi_4 = {dataInMem_hi_175, dataInMem_lo_111, dataInMem_hi_174, dataInMem_lo_110};
  wire [159:0]     dataInMem_hi_lo_hi_lo_4 = {dataInMem_hi_lo_hi_lo_hi_4, dataInMem_hi_lo_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_hi_hi_lo_4 = {dataInMem_hi_177, dataInMem_lo_113, dataInMem_hi_176, dataInMem_lo_112};
  wire [79:0]      dataInMem_hi_lo_hi_hi_hi_4 = {dataInMem_hi_179, dataInMem_lo_115, dataInMem_hi_178, dataInMem_lo_114};
  wire [159:0]     dataInMem_hi_lo_hi_hi_4 = {dataInMem_hi_lo_hi_hi_hi_4, dataInMem_hi_lo_hi_hi_lo_4};
  wire [319:0]     dataInMem_hi_lo_hi_4 = {dataInMem_hi_lo_hi_hi_4, dataInMem_hi_lo_hi_lo_4};
  wire [639:0]     dataInMem_hi_lo_4 = {dataInMem_hi_lo_hi_4, dataInMem_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_lo_lo_lo_4 = {dataInMem_hi_181, dataInMem_lo_117, dataInMem_hi_180, dataInMem_lo_116};
  wire [79:0]      dataInMem_hi_hi_lo_lo_hi_4 = {dataInMem_hi_183, dataInMem_lo_119, dataInMem_hi_182, dataInMem_lo_118};
  wire [159:0]     dataInMem_hi_hi_lo_lo_4 = {dataInMem_hi_hi_lo_lo_hi_4, dataInMem_hi_hi_lo_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_lo_hi_lo_4 = {dataInMem_hi_185, dataInMem_lo_121, dataInMem_hi_184, dataInMem_lo_120};
  wire [79:0]      dataInMem_hi_hi_lo_hi_hi_4 = {dataInMem_hi_187, dataInMem_lo_123, dataInMem_hi_186, dataInMem_lo_122};
  wire [159:0]     dataInMem_hi_hi_lo_hi_4 = {dataInMem_hi_hi_lo_hi_hi_4, dataInMem_hi_hi_lo_hi_lo_4};
  wire [319:0]     dataInMem_hi_hi_lo_4 = {dataInMem_hi_hi_lo_hi_4, dataInMem_hi_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_hi_lo_lo_4 = {dataInMem_hi_189, dataInMem_lo_125, dataInMem_hi_188, dataInMem_lo_124};
  wire [79:0]      dataInMem_hi_hi_hi_lo_hi_4 = {dataInMem_hi_191, dataInMem_lo_127, dataInMem_hi_190, dataInMem_lo_126};
  wire [159:0]     dataInMem_hi_hi_hi_lo_4 = {dataInMem_hi_hi_hi_lo_hi_4, dataInMem_hi_hi_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_hi_hi_lo_4 = {dataInMem_hi_193, dataInMem_lo_129, dataInMem_hi_192, dataInMem_lo_128};
  wire [79:0]      dataInMem_hi_hi_hi_hi_hi_4 = {dataInMem_hi_195, dataInMem_lo_131, dataInMem_hi_194, dataInMem_lo_130};
  wire [159:0]     dataInMem_hi_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_hi_lo_4};
  wire [319:0]     dataInMem_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_lo_4};
  wire [639:0]     dataInMem_hi_hi_68 = {dataInMem_hi_hi_hi_4, dataInMem_hi_hi_lo_4};
  wire [1279:0]    dataInMem_hi_196 = {dataInMem_hi_hi_68, dataInMem_hi_lo_4};
  wire [2559:0]    dataInMem_4 = {dataInMem_hi_196, dataInMem_lo_132};
  wire [511:0]     regroupCacheLine_4_0 = dataInMem_4[511:0];
  wire [511:0]     regroupCacheLine_4_1 = dataInMem_4[1023:512];
  wire [511:0]     regroupCacheLine_4_2 = dataInMem_4[1535:1024];
  wire [511:0]     regroupCacheLine_4_3 = dataInMem_4[2047:1536];
  wire [511:0]     regroupCacheLine_4_4 = dataInMem_4[2559:2048];
  wire [511:0]     res_32 = regroupCacheLine_4_0;
  wire [511:0]     res_33 = regroupCacheLine_4_1;
  wire [511:0]     res_34 = regroupCacheLine_4_2;
  wire [511:0]     res_35 = regroupCacheLine_4_3;
  wire [511:0]     res_36 = regroupCacheLine_4_4;
  wire [1023:0]    lo_lo_4 = {res_33, res_32};
  wire [1023:0]    lo_hi_4 = {res_35, res_34};
  wire [2047:0]    lo_4 = {lo_hi_4, lo_lo_4};
  wire [1023:0]    hi_lo_4 = {512'h0, res_36};
  wire [2047:0]    hi_4 = {1024'h0, hi_lo_4};
  wire [4095:0]    regroupLoadData_0_4 = {hi_4, lo_4};
  wire [23:0]      dataInMem_lo_133 = {dataInMem_lo_hi_5, dataRegroupBySew_0_0};
  wire [15:0]      _GEN_261 = {dataRegroupBySew_5_0, dataRegroupBySew_4_0};
  wire [15:0]      dataInMem_hi_hi_69;
  assign dataInMem_hi_hi_69 = _GEN_261;
  wire [15:0]      dataInMem_hi_lo_71;
  assign dataInMem_hi_lo_71 = _GEN_261;
  wire [23:0]      dataInMem_hi_197 = {dataInMem_hi_hi_69, dataRegroupBySew_3_0};
  wire [23:0]      dataInMem_lo_134 = {dataInMem_lo_hi_6, dataRegroupBySew_0_1};
  wire [15:0]      _GEN_262 = {dataRegroupBySew_5_1, dataRegroupBySew_4_1};
  wire [15:0]      dataInMem_hi_hi_70;
  assign dataInMem_hi_hi_70 = _GEN_262;
  wire [15:0]      dataInMem_hi_lo_72;
  assign dataInMem_hi_lo_72 = _GEN_262;
  wire [23:0]      dataInMem_hi_198 = {dataInMem_hi_hi_70, dataRegroupBySew_3_1};
  wire [23:0]      dataInMem_lo_135 = {dataInMem_lo_hi_7, dataRegroupBySew_0_2};
  wire [15:0]      _GEN_263 = {dataRegroupBySew_5_2, dataRegroupBySew_4_2};
  wire [15:0]      dataInMem_hi_hi_71;
  assign dataInMem_hi_hi_71 = _GEN_263;
  wire [15:0]      dataInMem_hi_lo_73;
  assign dataInMem_hi_lo_73 = _GEN_263;
  wire [23:0]      dataInMem_hi_199 = {dataInMem_hi_hi_71, dataRegroupBySew_3_2};
  wire [23:0]      dataInMem_lo_136 = {dataInMem_lo_hi_8, dataRegroupBySew_0_3};
  wire [15:0]      _GEN_264 = {dataRegroupBySew_5_3, dataRegroupBySew_4_3};
  wire [15:0]      dataInMem_hi_hi_72;
  assign dataInMem_hi_hi_72 = _GEN_264;
  wire [15:0]      dataInMem_hi_lo_74;
  assign dataInMem_hi_lo_74 = _GEN_264;
  wire [23:0]      dataInMem_hi_200 = {dataInMem_hi_hi_72, dataRegroupBySew_3_3};
  wire [23:0]      dataInMem_lo_137 = {dataInMem_lo_hi_9, dataRegroupBySew_0_4};
  wire [15:0]      _GEN_265 = {dataRegroupBySew_5_4, dataRegroupBySew_4_4};
  wire [15:0]      dataInMem_hi_hi_73;
  assign dataInMem_hi_hi_73 = _GEN_265;
  wire [15:0]      dataInMem_hi_lo_75;
  assign dataInMem_hi_lo_75 = _GEN_265;
  wire [23:0]      dataInMem_hi_201 = {dataInMem_hi_hi_73, dataRegroupBySew_3_4};
  wire [23:0]      dataInMem_lo_138 = {dataInMem_lo_hi_10, dataRegroupBySew_0_5};
  wire [15:0]      _GEN_266 = {dataRegroupBySew_5_5, dataRegroupBySew_4_5};
  wire [15:0]      dataInMem_hi_hi_74;
  assign dataInMem_hi_hi_74 = _GEN_266;
  wire [15:0]      dataInMem_hi_lo_76;
  assign dataInMem_hi_lo_76 = _GEN_266;
  wire [23:0]      dataInMem_hi_202 = {dataInMem_hi_hi_74, dataRegroupBySew_3_5};
  wire [23:0]      dataInMem_lo_139 = {dataInMem_lo_hi_11, dataRegroupBySew_0_6};
  wire [15:0]      _GEN_267 = {dataRegroupBySew_5_6, dataRegroupBySew_4_6};
  wire [15:0]      dataInMem_hi_hi_75;
  assign dataInMem_hi_hi_75 = _GEN_267;
  wire [15:0]      dataInMem_hi_lo_77;
  assign dataInMem_hi_lo_77 = _GEN_267;
  wire [23:0]      dataInMem_hi_203 = {dataInMem_hi_hi_75, dataRegroupBySew_3_6};
  wire [23:0]      dataInMem_lo_140 = {dataInMem_lo_hi_12, dataRegroupBySew_0_7};
  wire [15:0]      _GEN_268 = {dataRegroupBySew_5_7, dataRegroupBySew_4_7};
  wire [15:0]      dataInMem_hi_hi_76;
  assign dataInMem_hi_hi_76 = _GEN_268;
  wire [15:0]      dataInMem_hi_lo_78;
  assign dataInMem_hi_lo_78 = _GEN_268;
  wire [23:0]      dataInMem_hi_204 = {dataInMem_hi_hi_76, dataRegroupBySew_3_7};
  wire [23:0]      dataInMem_lo_141 = {dataInMem_lo_hi_13, dataRegroupBySew_0_8};
  wire [15:0]      _GEN_269 = {dataRegroupBySew_5_8, dataRegroupBySew_4_8};
  wire [15:0]      dataInMem_hi_hi_77;
  assign dataInMem_hi_hi_77 = _GEN_269;
  wire [15:0]      dataInMem_hi_lo_79;
  assign dataInMem_hi_lo_79 = _GEN_269;
  wire [23:0]      dataInMem_hi_205 = {dataInMem_hi_hi_77, dataRegroupBySew_3_8};
  wire [23:0]      dataInMem_lo_142 = {dataInMem_lo_hi_14, dataRegroupBySew_0_9};
  wire [15:0]      _GEN_270 = {dataRegroupBySew_5_9, dataRegroupBySew_4_9};
  wire [15:0]      dataInMem_hi_hi_78;
  assign dataInMem_hi_hi_78 = _GEN_270;
  wire [15:0]      dataInMem_hi_lo_80;
  assign dataInMem_hi_lo_80 = _GEN_270;
  wire [23:0]      dataInMem_hi_206 = {dataInMem_hi_hi_78, dataRegroupBySew_3_9};
  wire [23:0]      dataInMem_lo_143 = {dataInMem_lo_hi_15, dataRegroupBySew_0_10};
  wire [15:0]      _GEN_271 = {dataRegroupBySew_5_10, dataRegroupBySew_4_10};
  wire [15:0]      dataInMem_hi_hi_79;
  assign dataInMem_hi_hi_79 = _GEN_271;
  wire [15:0]      dataInMem_hi_lo_81;
  assign dataInMem_hi_lo_81 = _GEN_271;
  wire [23:0]      dataInMem_hi_207 = {dataInMem_hi_hi_79, dataRegroupBySew_3_10};
  wire [23:0]      dataInMem_lo_144 = {dataInMem_lo_hi_16, dataRegroupBySew_0_11};
  wire [15:0]      _GEN_272 = {dataRegroupBySew_5_11, dataRegroupBySew_4_11};
  wire [15:0]      dataInMem_hi_hi_80;
  assign dataInMem_hi_hi_80 = _GEN_272;
  wire [15:0]      dataInMem_hi_lo_82;
  assign dataInMem_hi_lo_82 = _GEN_272;
  wire [23:0]      dataInMem_hi_208 = {dataInMem_hi_hi_80, dataRegroupBySew_3_11};
  wire [23:0]      dataInMem_lo_145 = {dataInMem_lo_hi_17, dataRegroupBySew_0_12};
  wire [15:0]      _GEN_273 = {dataRegroupBySew_5_12, dataRegroupBySew_4_12};
  wire [15:0]      dataInMem_hi_hi_81;
  assign dataInMem_hi_hi_81 = _GEN_273;
  wire [15:0]      dataInMem_hi_lo_83;
  assign dataInMem_hi_lo_83 = _GEN_273;
  wire [23:0]      dataInMem_hi_209 = {dataInMem_hi_hi_81, dataRegroupBySew_3_12};
  wire [23:0]      dataInMem_lo_146 = {dataInMem_lo_hi_18, dataRegroupBySew_0_13};
  wire [15:0]      _GEN_274 = {dataRegroupBySew_5_13, dataRegroupBySew_4_13};
  wire [15:0]      dataInMem_hi_hi_82;
  assign dataInMem_hi_hi_82 = _GEN_274;
  wire [15:0]      dataInMem_hi_lo_84;
  assign dataInMem_hi_lo_84 = _GEN_274;
  wire [23:0]      dataInMem_hi_210 = {dataInMem_hi_hi_82, dataRegroupBySew_3_13};
  wire [23:0]      dataInMem_lo_147 = {dataInMem_lo_hi_19, dataRegroupBySew_0_14};
  wire [15:0]      _GEN_275 = {dataRegroupBySew_5_14, dataRegroupBySew_4_14};
  wire [15:0]      dataInMem_hi_hi_83;
  assign dataInMem_hi_hi_83 = _GEN_275;
  wire [15:0]      dataInMem_hi_lo_85;
  assign dataInMem_hi_lo_85 = _GEN_275;
  wire [23:0]      dataInMem_hi_211 = {dataInMem_hi_hi_83, dataRegroupBySew_3_14};
  wire [23:0]      dataInMem_lo_148 = {dataInMem_lo_hi_20, dataRegroupBySew_0_15};
  wire [15:0]      _GEN_276 = {dataRegroupBySew_5_15, dataRegroupBySew_4_15};
  wire [15:0]      dataInMem_hi_hi_84;
  assign dataInMem_hi_hi_84 = _GEN_276;
  wire [15:0]      dataInMem_hi_lo_86;
  assign dataInMem_hi_lo_86 = _GEN_276;
  wire [23:0]      dataInMem_hi_212 = {dataInMem_hi_hi_84, dataRegroupBySew_3_15};
  wire [23:0]      dataInMem_lo_149 = {dataInMem_lo_hi_21, dataRegroupBySew_0_16};
  wire [15:0]      _GEN_277 = {dataRegroupBySew_5_16, dataRegroupBySew_4_16};
  wire [15:0]      dataInMem_hi_hi_85;
  assign dataInMem_hi_hi_85 = _GEN_277;
  wire [15:0]      dataInMem_hi_lo_87;
  assign dataInMem_hi_lo_87 = _GEN_277;
  wire [23:0]      dataInMem_hi_213 = {dataInMem_hi_hi_85, dataRegroupBySew_3_16};
  wire [23:0]      dataInMem_lo_150 = {dataInMem_lo_hi_22, dataRegroupBySew_0_17};
  wire [15:0]      _GEN_278 = {dataRegroupBySew_5_17, dataRegroupBySew_4_17};
  wire [15:0]      dataInMem_hi_hi_86;
  assign dataInMem_hi_hi_86 = _GEN_278;
  wire [15:0]      dataInMem_hi_lo_88;
  assign dataInMem_hi_lo_88 = _GEN_278;
  wire [23:0]      dataInMem_hi_214 = {dataInMem_hi_hi_86, dataRegroupBySew_3_17};
  wire [23:0]      dataInMem_lo_151 = {dataInMem_lo_hi_23, dataRegroupBySew_0_18};
  wire [15:0]      _GEN_279 = {dataRegroupBySew_5_18, dataRegroupBySew_4_18};
  wire [15:0]      dataInMem_hi_hi_87;
  assign dataInMem_hi_hi_87 = _GEN_279;
  wire [15:0]      dataInMem_hi_lo_89;
  assign dataInMem_hi_lo_89 = _GEN_279;
  wire [23:0]      dataInMem_hi_215 = {dataInMem_hi_hi_87, dataRegroupBySew_3_18};
  wire [23:0]      dataInMem_lo_152 = {dataInMem_lo_hi_24, dataRegroupBySew_0_19};
  wire [15:0]      _GEN_280 = {dataRegroupBySew_5_19, dataRegroupBySew_4_19};
  wire [15:0]      dataInMem_hi_hi_88;
  assign dataInMem_hi_hi_88 = _GEN_280;
  wire [15:0]      dataInMem_hi_lo_90;
  assign dataInMem_hi_lo_90 = _GEN_280;
  wire [23:0]      dataInMem_hi_216 = {dataInMem_hi_hi_88, dataRegroupBySew_3_19};
  wire [23:0]      dataInMem_lo_153 = {dataInMem_lo_hi_25, dataRegroupBySew_0_20};
  wire [15:0]      _GEN_281 = {dataRegroupBySew_5_20, dataRegroupBySew_4_20};
  wire [15:0]      dataInMem_hi_hi_89;
  assign dataInMem_hi_hi_89 = _GEN_281;
  wire [15:0]      dataInMem_hi_lo_91;
  assign dataInMem_hi_lo_91 = _GEN_281;
  wire [23:0]      dataInMem_hi_217 = {dataInMem_hi_hi_89, dataRegroupBySew_3_20};
  wire [23:0]      dataInMem_lo_154 = {dataInMem_lo_hi_26, dataRegroupBySew_0_21};
  wire [15:0]      _GEN_282 = {dataRegroupBySew_5_21, dataRegroupBySew_4_21};
  wire [15:0]      dataInMem_hi_hi_90;
  assign dataInMem_hi_hi_90 = _GEN_282;
  wire [15:0]      dataInMem_hi_lo_92;
  assign dataInMem_hi_lo_92 = _GEN_282;
  wire [23:0]      dataInMem_hi_218 = {dataInMem_hi_hi_90, dataRegroupBySew_3_21};
  wire [23:0]      dataInMem_lo_155 = {dataInMem_lo_hi_27, dataRegroupBySew_0_22};
  wire [15:0]      _GEN_283 = {dataRegroupBySew_5_22, dataRegroupBySew_4_22};
  wire [15:0]      dataInMem_hi_hi_91;
  assign dataInMem_hi_hi_91 = _GEN_283;
  wire [15:0]      dataInMem_hi_lo_93;
  assign dataInMem_hi_lo_93 = _GEN_283;
  wire [23:0]      dataInMem_hi_219 = {dataInMem_hi_hi_91, dataRegroupBySew_3_22};
  wire [23:0]      dataInMem_lo_156 = {dataInMem_lo_hi_28, dataRegroupBySew_0_23};
  wire [15:0]      _GEN_284 = {dataRegroupBySew_5_23, dataRegroupBySew_4_23};
  wire [15:0]      dataInMem_hi_hi_92;
  assign dataInMem_hi_hi_92 = _GEN_284;
  wire [15:0]      dataInMem_hi_lo_94;
  assign dataInMem_hi_lo_94 = _GEN_284;
  wire [23:0]      dataInMem_hi_220 = {dataInMem_hi_hi_92, dataRegroupBySew_3_23};
  wire [23:0]      dataInMem_lo_157 = {dataInMem_lo_hi_29, dataRegroupBySew_0_24};
  wire [15:0]      _GEN_285 = {dataRegroupBySew_5_24, dataRegroupBySew_4_24};
  wire [15:0]      dataInMem_hi_hi_93;
  assign dataInMem_hi_hi_93 = _GEN_285;
  wire [15:0]      dataInMem_hi_lo_95;
  assign dataInMem_hi_lo_95 = _GEN_285;
  wire [23:0]      dataInMem_hi_221 = {dataInMem_hi_hi_93, dataRegroupBySew_3_24};
  wire [23:0]      dataInMem_lo_158 = {dataInMem_lo_hi_30, dataRegroupBySew_0_25};
  wire [15:0]      _GEN_286 = {dataRegroupBySew_5_25, dataRegroupBySew_4_25};
  wire [15:0]      dataInMem_hi_hi_94;
  assign dataInMem_hi_hi_94 = _GEN_286;
  wire [15:0]      dataInMem_hi_lo_96;
  assign dataInMem_hi_lo_96 = _GEN_286;
  wire [23:0]      dataInMem_hi_222 = {dataInMem_hi_hi_94, dataRegroupBySew_3_25};
  wire [23:0]      dataInMem_lo_159 = {dataInMem_lo_hi_31, dataRegroupBySew_0_26};
  wire [15:0]      _GEN_287 = {dataRegroupBySew_5_26, dataRegroupBySew_4_26};
  wire [15:0]      dataInMem_hi_hi_95;
  assign dataInMem_hi_hi_95 = _GEN_287;
  wire [15:0]      dataInMem_hi_lo_97;
  assign dataInMem_hi_lo_97 = _GEN_287;
  wire [23:0]      dataInMem_hi_223 = {dataInMem_hi_hi_95, dataRegroupBySew_3_26};
  wire [23:0]      dataInMem_lo_160 = {dataInMem_lo_hi_32, dataRegroupBySew_0_27};
  wire [15:0]      _GEN_288 = {dataRegroupBySew_5_27, dataRegroupBySew_4_27};
  wire [15:0]      dataInMem_hi_hi_96;
  assign dataInMem_hi_hi_96 = _GEN_288;
  wire [15:0]      dataInMem_hi_lo_98;
  assign dataInMem_hi_lo_98 = _GEN_288;
  wire [23:0]      dataInMem_hi_224 = {dataInMem_hi_hi_96, dataRegroupBySew_3_27};
  wire [23:0]      dataInMem_lo_161 = {dataInMem_lo_hi_33, dataRegroupBySew_0_28};
  wire [15:0]      _GEN_289 = {dataRegroupBySew_5_28, dataRegroupBySew_4_28};
  wire [15:0]      dataInMem_hi_hi_97;
  assign dataInMem_hi_hi_97 = _GEN_289;
  wire [15:0]      dataInMem_hi_lo_99;
  assign dataInMem_hi_lo_99 = _GEN_289;
  wire [23:0]      dataInMem_hi_225 = {dataInMem_hi_hi_97, dataRegroupBySew_3_28};
  wire [23:0]      dataInMem_lo_162 = {dataInMem_lo_hi_34, dataRegroupBySew_0_29};
  wire [15:0]      _GEN_290 = {dataRegroupBySew_5_29, dataRegroupBySew_4_29};
  wire [15:0]      dataInMem_hi_hi_98;
  assign dataInMem_hi_hi_98 = _GEN_290;
  wire [15:0]      dataInMem_hi_lo_100;
  assign dataInMem_hi_lo_100 = _GEN_290;
  wire [23:0]      dataInMem_hi_226 = {dataInMem_hi_hi_98, dataRegroupBySew_3_29};
  wire [23:0]      dataInMem_lo_163 = {dataInMem_lo_hi_35, dataRegroupBySew_0_30};
  wire [15:0]      _GEN_291 = {dataRegroupBySew_5_30, dataRegroupBySew_4_30};
  wire [15:0]      dataInMem_hi_hi_99;
  assign dataInMem_hi_hi_99 = _GEN_291;
  wire [15:0]      dataInMem_hi_lo_101;
  assign dataInMem_hi_lo_101 = _GEN_291;
  wire [23:0]      dataInMem_hi_227 = {dataInMem_hi_hi_99, dataRegroupBySew_3_30};
  wire [23:0]      dataInMem_lo_164 = {dataInMem_lo_hi_36, dataRegroupBySew_0_31};
  wire [15:0]      _GEN_292 = {dataRegroupBySew_5_31, dataRegroupBySew_4_31};
  wire [15:0]      dataInMem_hi_hi_100;
  assign dataInMem_hi_hi_100 = _GEN_292;
  wire [15:0]      dataInMem_hi_lo_102;
  assign dataInMem_hi_lo_102 = _GEN_292;
  wire [23:0]      dataInMem_hi_228 = {dataInMem_hi_hi_100, dataRegroupBySew_3_31};
  wire [23:0]      dataInMem_lo_165 = {dataInMem_lo_hi_37, dataRegroupBySew_0_32};
  wire [15:0]      _GEN_293 = {dataRegroupBySew_5_32, dataRegroupBySew_4_32};
  wire [15:0]      dataInMem_hi_hi_101;
  assign dataInMem_hi_hi_101 = _GEN_293;
  wire [15:0]      dataInMem_hi_lo_103;
  assign dataInMem_hi_lo_103 = _GEN_293;
  wire [23:0]      dataInMem_hi_229 = {dataInMem_hi_hi_101, dataRegroupBySew_3_32};
  wire [23:0]      dataInMem_lo_166 = {dataInMem_lo_hi_38, dataRegroupBySew_0_33};
  wire [15:0]      _GEN_294 = {dataRegroupBySew_5_33, dataRegroupBySew_4_33};
  wire [15:0]      dataInMem_hi_hi_102;
  assign dataInMem_hi_hi_102 = _GEN_294;
  wire [15:0]      dataInMem_hi_lo_104;
  assign dataInMem_hi_lo_104 = _GEN_294;
  wire [23:0]      dataInMem_hi_230 = {dataInMem_hi_hi_102, dataRegroupBySew_3_33};
  wire [23:0]      dataInMem_lo_167 = {dataInMem_lo_hi_39, dataRegroupBySew_0_34};
  wire [15:0]      _GEN_295 = {dataRegroupBySew_5_34, dataRegroupBySew_4_34};
  wire [15:0]      dataInMem_hi_hi_103;
  assign dataInMem_hi_hi_103 = _GEN_295;
  wire [15:0]      dataInMem_hi_lo_105;
  assign dataInMem_hi_lo_105 = _GEN_295;
  wire [23:0]      dataInMem_hi_231 = {dataInMem_hi_hi_103, dataRegroupBySew_3_34};
  wire [23:0]      dataInMem_lo_168 = {dataInMem_lo_hi_40, dataRegroupBySew_0_35};
  wire [15:0]      _GEN_296 = {dataRegroupBySew_5_35, dataRegroupBySew_4_35};
  wire [15:0]      dataInMem_hi_hi_104;
  assign dataInMem_hi_hi_104 = _GEN_296;
  wire [15:0]      dataInMem_hi_lo_106;
  assign dataInMem_hi_lo_106 = _GEN_296;
  wire [23:0]      dataInMem_hi_232 = {dataInMem_hi_hi_104, dataRegroupBySew_3_35};
  wire [23:0]      dataInMem_lo_169 = {dataInMem_lo_hi_41, dataRegroupBySew_0_36};
  wire [15:0]      _GEN_297 = {dataRegroupBySew_5_36, dataRegroupBySew_4_36};
  wire [15:0]      dataInMem_hi_hi_105;
  assign dataInMem_hi_hi_105 = _GEN_297;
  wire [15:0]      dataInMem_hi_lo_107;
  assign dataInMem_hi_lo_107 = _GEN_297;
  wire [23:0]      dataInMem_hi_233 = {dataInMem_hi_hi_105, dataRegroupBySew_3_36};
  wire [23:0]      dataInMem_lo_170 = {dataInMem_lo_hi_42, dataRegroupBySew_0_37};
  wire [15:0]      _GEN_298 = {dataRegroupBySew_5_37, dataRegroupBySew_4_37};
  wire [15:0]      dataInMem_hi_hi_106;
  assign dataInMem_hi_hi_106 = _GEN_298;
  wire [15:0]      dataInMem_hi_lo_108;
  assign dataInMem_hi_lo_108 = _GEN_298;
  wire [23:0]      dataInMem_hi_234 = {dataInMem_hi_hi_106, dataRegroupBySew_3_37};
  wire [23:0]      dataInMem_lo_171 = {dataInMem_lo_hi_43, dataRegroupBySew_0_38};
  wire [15:0]      _GEN_299 = {dataRegroupBySew_5_38, dataRegroupBySew_4_38};
  wire [15:0]      dataInMem_hi_hi_107;
  assign dataInMem_hi_hi_107 = _GEN_299;
  wire [15:0]      dataInMem_hi_lo_109;
  assign dataInMem_hi_lo_109 = _GEN_299;
  wire [23:0]      dataInMem_hi_235 = {dataInMem_hi_hi_107, dataRegroupBySew_3_38};
  wire [23:0]      dataInMem_lo_172 = {dataInMem_lo_hi_44, dataRegroupBySew_0_39};
  wire [15:0]      _GEN_300 = {dataRegroupBySew_5_39, dataRegroupBySew_4_39};
  wire [15:0]      dataInMem_hi_hi_108;
  assign dataInMem_hi_hi_108 = _GEN_300;
  wire [15:0]      dataInMem_hi_lo_110;
  assign dataInMem_hi_lo_110 = _GEN_300;
  wire [23:0]      dataInMem_hi_236 = {dataInMem_hi_hi_108, dataRegroupBySew_3_39};
  wire [23:0]      dataInMem_lo_173 = {dataInMem_lo_hi_45, dataRegroupBySew_0_40};
  wire [15:0]      _GEN_301 = {dataRegroupBySew_5_40, dataRegroupBySew_4_40};
  wire [15:0]      dataInMem_hi_hi_109;
  assign dataInMem_hi_hi_109 = _GEN_301;
  wire [15:0]      dataInMem_hi_lo_111;
  assign dataInMem_hi_lo_111 = _GEN_301;
  wire [23:0]      dataInMem_hi_237 = {dataInMem_hi_hi_109, dataRegroupBySew_3_40};
  wire [23:0]      dataInMem_lo_174 = {dataInMem_lo_hi_46, dataRegroupBySew_0_41};
  wire [15:0]      _GEN_302 = {dataRegroupBySew_5_41, dataRegroupBySew_4_41};
  wire [15:0]      dataInMem_hi_hi_110;
  assign dataInMem_hi_hi_110 = _GEN_302;
  wire [15:0]      dataInMem_hi_lo_112;
  assign dataInMem_hi_lo_112 = _GEN_302;
  wire [23:0]      dataInMem_hi_238 = {dataInMem_hi_hi_110, dataRegroupBySew_3_41};
  wire [23:0]      dataInMem_lo_175 = {dataInMem_lo_hi_47, dataRegroupBySew_0_42};
  wire [15:0]      _GEN_303 = {dataRegroupBySew_5_42, dataRegroupBySew_4_42};
  wire [15:0]      dataInMem_hi_hi_111;
  assign dataInMem_hi_hi_111 = _GEN_303;
  wire [15:0]      dataInMem_hi_lo_113;
  assign dataInMem_hi_lo_113 = _GEN_303;
  wire [23:0]      dataInMem_hi_239 = {dataInMem_hi_hi_111, dataRegroupBySew_3_42};
  wire [23:0]      dataInMem_lo_176 = {dataInMem_lo_hi_48, dataRegroupBySew_0_43};
  wire [15:0]      _GEN_304 = {dataRegroupBySew_5_43, dataRegroupBySew_4_43};
  wire [15:0]      dataInMem_hi_hi_112;
  assign dataInMem_hi_hi_112 = _GEN_304;
  wire [15:0]      dataInMem_hi_lo_114;
  assign dataInMem_hi_lo_114 = _GEN_304;
  wire [23:0]      dataInMem_hi_240 = {dataInMem_hi_hi_112, dataRegroupBySew_3_43};
  wire [23:0]      dataInMem_lo_177 = {dataInMem_lo_hi_49, dataRegroupBySew_0_44};
  wire [15:0]      _GEN_305 = {dataRegroupBySew_5_44, dataRegroupBySew_4_44};
  wire [15:0]      dataInMem_hi_hi_113;
  assign dataInMem_hi_hi_113 = _GEN_305;
  wire [15:0]      dataInMem_hi_lo_115;
  assign dataInMem_hi_lo_115 = _GEN_305;
  wire [23:0]      dataInMem_hi_241 = {dataInMem_hi_hi_113, dataRegroupBySew_3_44};
  wire [23:0]      dataInMem_lo_178 = {dataInMem_lo_hi_50, dataRegroupBySew_0_45};
  wire [15:0]      _GEN_306 = {dataRegroupBySew_5_45, dataRegroupBySew_4_45};
  wire [15:0]      dataInMem_hi_hi_114;
  assign dataInMem_hi_hi_114 = _GEN_306;
  wire [15:0]      dataInMem_hi_lo_116;
  assign dataInMem_hi_lo_116 = _GEN_306;
  wire [23:0]      dataInMem_hi_242 = {dataInMem_hi_hi_114, dataRegroupBySew_3_45};
  wire [23:0]      dataInMem_lo_179 = {dataInMem_lo_hi_51, dataRegroupBySew_0_46};
  wire [15:0]      _GEN_307 = {dataRegroupBySew_5_46, dataRegroupBySew_4_46};
  wire [15:0]      dataInMem_hi_hi_115;
  assign dataInMem_hi_hi_115 = _GEN_307;
  wire [15:0]      dataInMem_hi_lo_117;
  assign dataInMem_hi_lo_117 = _GEN_307;
  wire [23:0]      dataInMem_hi_243 = {dataInMem_hi_hi_115, dataRegroupBySew_3_46};
  wire [23:0]      dataInMem_lo_180 = {dataInMem_lo_hi_52, dataRegroupBySew_0_47};
  wire [15:0]      _GEN_308 = {dataRegroupBySew_5_47, dataRegroupBySew_4_47};
  wire [15:0]      dataInMem_hi_hi_116;
  assign dataInMem_hi_hi_116 = _GEN_308;
  wire [15:0]      dataInMem_hi_lo_118;
  assign dataInMem_hi_lo_118 = _GEN_308;
  wire [23:0]      dataInMem_hi_244 = {dataInMem_hi_hi_116, dataRegroupBySew_3_47};
  wire [23:0]      dataInMem_lo_181 = {dataInMem_lo_hi_53, dataRegroupBySew_0_48};
  wire [15:0]      _GEN_309 = {dataRegroupBySew_5_48, dataRegroupBySew_4_48};
  wire [15:0]      dataInMem_hi_hi_117;
  assign dataInMem_hi_hi_117 = _GEN_309;
  wire [15:0]      dataInMem_hi_lo_119;
  assign dataInMem_hi_lo_119 = _GEN_309;
  wire [23:0]      dataInMem_hi_245 = {dataInMem_hi_hi_117, dataRegroupBySew_3_48};
  wire [23:0]      dataInMem_lo_182 = {dataInMem_lo_hi_54, dataRegroupBySew_0_49};
  wire [15:0]      _GEN_310 = {dataRegroupBySew_5_49, dataRegroupBySew_4_49};
  wire [15:0]      dataInMem_hi_hi_118;
  assign dataInMem_hi_hi_118 = _GEN_310;
  wire [15:0]      dataInMem_hi_lo_120;
  assign dataInMem_hi_lo_120 = _GEN_310;
  wire [23:0]      dataInMem_hi_246 = {dataInMem_hi_hi_118, dataRegroupBySew_3_49};
  wire [23:0]      dataInMem_lo_183 = {dataInMem_lo_hi_55, dataRegroupBySew_0_50};
  wire [15:0]      _GEN_311 = {dataRegroupBySew_5_50, dataRegroupBySew_4_50};
  wire [15:0]      dataInMem_hi_hi_119;
  assign dataInMem_hi_hi_119 = _GEN_311;
  wire [15:0]      dataInMem_hi_lo_121;
  assign dataInMem_hi_lo_121 = _GEN_311;
  wire [23:0]      dataInMem_hi_247 = {dataInMem_hi_hi_119, dataRegroupBySew_3_50};
  wire [23:0]      dataInMem_lo_184 = {dataInMem_lo_hi_56, dataRegroupBySew_0_51};
  wire [15:0]      _GEN_312 = {dataRegroupBySew_5_51, dataRegroupBySew_4_51};
  wire [15:0]      dataInMem_hi_hi_120;
  assign dataInMem_hi_hi_120 = _GEN_312;
  wire [15:0]      dataInMem_hi_lo_122;
  assign dataInMem_hi_lo_122 = _GEN_312;
  wire [23:0]      dataInMem_hi_248 = {dataInMem_hi_hi_120, dataRegroupBySew_3_51};
  wire [23:0]      dataInMem_lo_185 = {dataInMem_lo_hi_57, dataRegroupBySew_0_52};
  wire [15:0]      _GEN_313 = {dataRegroupBySew_5_52, dataRegroupBySew_4_52};
  wire [15:0]      dataInMem_hi_hi_121;
  assign dataInMem_hi_hi_121 = _GEN_313;
  wire [15:0]      dataInMem_hi_lo_123;
  assign dataInMem_hi_lo_123 = _GEN_313;
  wire [23:0]      dataInMem_hi_249 = {dataInMem_hi_hi_121, dataRegroupBySew_3_52};
  wire [23:0]      dataInMem_lo_186 = {dataInMem_lo_hi_58, dataRegroupBySew_0_53};
  wire [15:0]      _GEN_314 = {dataRegroupBySew_5_53, dataRegroupBySew_4_53};
  wire [15:0]      dataInMem_hi_hi_122;
  assign dataInMem_hi_hi_122 = _GEN_314;
  wire [15:0]      dataInMem_hi_lo_124;
  assign dataInMem_hi_lo_124 = _GEN_314;
  wire [23:0]      dataInMem_hi_250 = {dataInMem_hi_hi_122, dataRegroupBySew_3_53};
  wire [23:0]      dataInMem_lo_187 = {dataInMem_lo_hi_59, dataRegroupBySew_0_54};
  wire [15:0]      _GEN_315 = {dataRegroupBySew_5_54, dataRegroupBySew_4_54};
  wire [15:0]      dataInMem_hi_hi_123;
  assign dataInMem_hi_hi_123 = _GEN_315;
  wire [15:0]      dataInMem_hi_lo_125;
  assign dataInMem_hi_lo_125 = _GEN_315;
  wire [23:0]      dataInMem_hi_251 = {dataInMem_hi_hi_123, dataRegroupBySew_3_54};
  wire [23:0]      dataInMem_lo_188 = {dataInMem_lo_hi_60, dataRegroupBySew_0_55};
  wire [15:0]      _GEN_316 = {dataRegroupBySew_5_55, dataRegroupBySew_4_55};
  wire [15:0]      dataInMem_hi_hi_124;
  assign dataInMem_hi_hi_124 = _GEN_316;
  wire [15:0]      dataInMem_hi_lo_126;
  assign dataInMem_hi_lo_126 = _GEN_316;
  wire [23:0]      dataInMem_hi_252 = {dataInMem_hi_hi_124, dataRegroupBySew_3_55};
  wire [23:0]      dataInMem_lo_189 = {dataInMem_lo_hi_61, dataRegroupBySew_0_56};
  wire [15:0]      _GEN_317 = {dataRegroupBySew_5_56, dataRegroupBySew_4_56};
  wire [15:0]      dataInMem_hi_hi_125;
  assign dataInMem_hi_hi_125 = _GEN_317;
  wire [15:0]      dataInMem_hi_lo_127;
  assign dataInMem_hi_lo_127 = _GEN_317;
  wire [23:0]      dataInMem_hi_253 = {dataInMem_hi_hi_125, dataRegroupBySew_3_56};
  wire [23:0]      dataInMem_lo_190 = {dataInMem_lo_hi_62, dataRegroupBySew_0_57};
  wire [15:0]      _GEN_318 = {dataRegroupBySew_5_57, dataRegroupBySew_4_57};
  wire [15:0]      dataInMem_hi_hi_126;
  assign dataInMem_hi_hi_126 = _GEN_318;
  wire [15:0]      dataInMem_hi_lo_128;
  assign dataInMem_hi_lo_128 = _GEN_318;
  wire [23:0]      dataInMem_hi_254 = {dataInMem_hi_hi_126, dataRegroupBySew_3_57};
  wire [23:0]      dataInMem_lo_191 = {dataInMem_lo_hi_63, dataRegroupBySew_0_58};
  wire [15:0]      _GEN_319 = {dataRegroupBySew_5_58, dataRegroupBySew_4_58};
  wire [15:0]      dataInMem_hi_hi_127;
  assign dataInMem_hi_hi_127 = _GEN_319;
  wire [15:0]      dataInMem_hi_lo_129;
  assign dataInMem_hi_lo_129 = _GEN_319;
  wire [23:0]      dataInMem_hi_255 = {dataInMem_hi_hi_127, dataRegroupBySew_3_58};
  wire [23:0]      dataInMem_lo_192 = {dataInMem_lo_hi_64, dataRegroupBySew_0_59};
  wire [15:0]      _GEN_320 = {dataRegroupBySew_5_59, dataRegroupBySew_4_59};
  wire [15:0]      dataInMem_hi_hi_128;
  assign dataInMem_hi_hi_128 = _GEN_320;
  wire [15:0]      dataInMem_hi_lo_130;
  assign dataInMem_hi_lo_130 = _GEN_320;
  wire [23:0]      dataInMem_hi_256 = {dataInMem_hi_hi_128, dataRegroupBySew_3_59};
  wire [23:0]      dataInMem_lo_193 = {dataInMem_lo_hi_65, dataRegroupBySew_0_60};
  wire [15:0]      _GEN_321 = {dataRegroupBySew_5_60, dataRegroupBySew_4_60};
  wire [15:0]      dataInMem_hi_hi_129;
  assign dataInMem_hi_hi_129 = _GEN_321;
  wire [15:0]      dataInMem_hi_lo_131;
  assign dataInMem_hi_lo_131 = _GEN_321;
  wire [23:0]      dataInMem_hi_257 = {dataInMem_hi_hi_129, dataRegroupBySew_3_60};
  wire [23:0]      dataInMem_lo_194 = {dataInMem_lo_hi_66, dataRegroupBySew_0_61};
  wire [15:0]      _GEN_322 = {dataRegroupBySew_5_61, dataRegroupBySew_4_61};
  wire [15:0]      dataInMem_hi_hi_130;
  assign dataInMem_hi_hi_130 = _GEN_322;
  wire [15:0]      dataInMem_hi_lo_132;
  assign dataInMem_hi_lo_132 = _GEN_322;
  wire [23:0]      dataInMem_hi_258 = {dataInMem_hi_hi_130, dataRegroupBySew_3_61};
  wire [23:0]      dataInMem_lo_195 = {dataInMem_lo_hi_67, dataRegroupBySew_0_62};
  wire [15:0]      _GEN_323 = {dataRegroupBySew_5_62, dataRegroupBySew_4_62};
  wire [15:0]      dataInMem_hi_hi_131;
  assign dataInMem_hi_hi_131 = _GEN_323;
  wire [15:0]      dataInMem_hi_lo_133;
  assign dataInMem_hi_lo_133 = _GEN_323;
  wire [23:0]      dataInMem_hi_259 = {dataInMem_hi_hi_131, dataRegroupBySew_3_62};
  wire [23:0]      dataInMem_lo_196 = {dataInMem_lo_hi_68, dataRegroupBySew_0_63};
  wire [15:0]      _GEN_324 = {dataRegroupBySew_5_63, dataRegroupBySew_4_63};
  wire [15:0]      dataInMem_hi_hi_132;
  assign dataInMem_hi_hi_132 = _GEN_324;
  wire [15:0]      dataInMem_hi_lo_134;
  assign dataInMem_hi_lo_134 = _GEN_324;
  wire [23:0]      dataInMem_hi_260 = {dataInMem_hi_hi_132, dataRegroupBySew_3_63};
  wire [95:0]      dataInMem_lo_lo_lo_lo_lo_5 = {dataInMem_hi_198, dataInMem_lo_134, dataInMem_hi_197, dataInMem_lo_133};
  wire [95:0]      dataInMem_lo_lo_lo_lo_hi_5 = {dataInMem_hi_200, dataInMem_lo_136, dataInMem_hi_199, dataInMem_lo_135};
  wire [191:0]     dataInMem_lo_lo_lo_lo_5 = {dataInMem_lo_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_lo_lo_hi_lo_5 = {dataInMem_hi_202, dataInMem_lo_138, dataInMem_hi_201, dataInMem_lo_137};
  wire [95:0]      dataInMem_lo_lo_lo_hi_hi_5 = {dataInMem_hi_204, dataInMem_lo_140, dataInMem_hi_203, dataInMem_lo_139};
  wire [191:0]     dataInMem_lo_lo_lo_hi_5 = {dataInMem_lo_lo_lo_hi_hi_5, dataInMem_lo_lo_lo_hi_lo_5};
  wire [383:0]     dataInMem_lo_lo_lo_5 = {dataInMem_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_lo_hi_lo_lo_5 = {dataInMem_hi_206, dataInMem_lo_142, dataInMem_hi_205, dataInMem_lo_141};
  wire [95:0]      dataInMem_lo_lo_hi_lo_hi_5 = {dataInMem_hi_208, dataInMem_lo_144, dataInMem_hi_207, dataInMem_lo_143};
  wire [191:0]     dataInMem_lo_lo_hi_lo_5 = {dataInMem_lo_lo_hi_lo_hi_5, dataInMem_lo_lo_hi_lo_lo_5};
  wire [95:0]      dataInMem_lo_lo_hi_hi_lo_5 = {dataInMem_hi_210, dataInMem_lo_146, dataInMem_hi_209, dataInMem_lo_145};
  wire [95:0]      dataInMem_lo_lo_hi_hi_hi_5 = {dataInMem_hi_212, dataInMem_lo_148, dataInMem_hi_211, dataInMem_lo_147};
  wire [191:0]     dataInMem_lo_lo_hi_hi_5 = {dataInMem_lo_lo_hi_hi_hi_5, dataInMem_lo_lo_hi_hi_lo_5};
  wire [383:0]     dataInMem_lo_lo_hi_5 = {dataInMem_lo_lo_hi_hi_5, dataInMem_lo_lo_hi_lo_5};
  wire [767:0]     dataInMem_lo_lo_5 = {dataInMem_lo_lo_hi_5, dataInMem_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_lo_lo_lo_5 = {dataInMem_hi_214, dataInMem_lo_150, dataInMem_hi_213, dataInMem_lo_149};
  wire [95:0]      dataInMem_lo_hi_lo_lo_hi_5 = {dataInMem_hi_216, dataInMem_lo_152, dataInMem_hi_215, dataInMem_lo_151};
  wire [191:0]     dataInMem_lo_hi_lo_lo_5 = {dataInMem_lo_hi_lo_lo_hi_5, dataInMem_lo_hi_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_lo_hi_lo_5 = {dataInMem_hi_218, dataInMem_lo_154, dataInMem_hi_217, dataInMem_lo_153};
  wire [95:0]      dataInMem_lo_hi_lo_hi_hi_5 = {dataInMem_hi_220, dataInMem_lo_156, dataInMem_hi_219, dataInMem_lo_155};
  wire [191:0]     dataInMem_lo_hi_lo_hi_5 = {dataInMem_lo_hi_lo_hi_hi_5, dataInMem_lo_hi_lo_hi_lo_5};
  wire [383:0]     dataInMem_lo_hi_lo_5 = {dataInMem_lo_hi_lo_hi_5, dataInMem_lo_hi_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_hi_lo_lo_5 = {dataInMem_hi_222, dataInMem_lo_158, dataInMem_hi_221, dataInMem_lo_157};
  wire [95:0]      dataInMem_lo_hi_hi_lo_hi_5 = {dataInMem_hi_224, dataInMem_lo_160, dataInMem_hi_223, dataInMem_lo_159};
  wire [191:0]     dataInMem_lo_hi_hi_lo_5 = {dataInMem_lo_hi_hi_lo_hi_5, dataInMem_lo_hi_hi_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_hi_hi_lo_5 = {dataInMem_hi_226, dataInMem_lo_162, dataInMem_hi_225, dataInMem_lo_161};
  wire [95:0]      dataInMem_lo_hi_hi_hi_hi_5 = {dataInMem_hi_228, dataInMem_lo_164, dataInMem_hi_227, dataInMem_lo_163};
  wire [191:0]     dataInMem_lo_hi_hi_hi_5 = {dataInMem_lo_hi_hi_hi_hi_5, dataInMem_lo_hi_hi_hi_lo_5};
  wire [383:0]     dataInMem_lo_hi_hi_5 = {dataInMem_lo_hi_hi_hi_5, dataInMem_lo_hi_hi_lo_5};
  wire [767:0]     dataInMem_lo_hi_69 = {dataInMem_lo_hi_hi_5, dataInMem_lo_hi_lo_5};
  wire [1535:0]    dataInMem_lo_197 = {dataInMem_lo_hi_69, dataInMem_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_lo_lo_lo_5 = {dataInMem_hi_230, dataInMem_lo_166, dataInMem_hi_229, dataInMem_lo_165};
  wire [95:0]      dataInMem_hi_lo_lo_lo_hi_5 = {dataInMem_hi_232, dataInMem_lo_168, dataInMem_hi_231, dataInMem_lo_167};
  wire [191:0]     dataInMem_hi_lo_lo_lo_5 = {dataInMem_hi_lo_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_lo_hi_lo_5 = {dataInMem_hi_234, dataInMem_lo_170, dataInMem_hi_233, dataInMem_lo_169};
  wire [95:0]      dataInMem_hi_lo_lo_hi_hi_5 = {dataInMem_hi_236, dataInMem_lo_172, dataInMem_hi_235, dataInMem_lo_171};
  wire [191:0]     dataInMem_hi_lo_lo_hi_5 = {dataInMem_hi_lo_lo_hi_hi_5, dataInMem_hi_lo_lo_hi_lo_5};
  wire [383:0]     dataInMem_hi_lo_lo_5 = {dataInMem_hi_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_hi_lo_lo_5 = {dataInMem_hi_238, dataInMem_lo_174, dataInMem_hi_237, dataInMem_lo_173};
  wire [95:0]      dataInMem_hi_lo_hi_lo_hi_5 = {dataInMem_hi_240, dataInMem_lo_176, dataInMem_hi_239, dataInMem_lo_175};
  wire [191:0]     dataInMem_hi_lo_hi_lo_5 = {dataInMem_hi_lo_hi_lo_hi_5, dataInMem_hi_lo_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_hi_hi_lo_5 = {dataInMem_hi_242, dataInMem_lo_178, dataInMem_hi_241, dataInMem_lo_177};
  wire [95:0]      dataInMem_hi_lo_hi_hi_hi_5 = {dataInMem_hi_244, dataInMem_lo_180, dataInMem_hi_243, dataInMem_lo_179};
  wire [191:0]     dataInMem_hi_lo_hi_hi_5 = {dataInMem_hi_lo_hi_hi_hi_5, dataInMem_hi_lo_hi_hi_lo_5};
  wire [383:0]     dataInMem_hi_lo_hi_5 = {dataInMem_hi_lo_hi_hi_5, dataInMem_hi_lo_hi_lo_5};
  wire [767:0]     dataInMem_hi_lo_5 = {dataInMem_hi_lo_hi_5, dataInMem_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_lo_lo_lo_5 = {dataInMem_hi_246, dataInMem_lo_182, dataInMem_hi_245, dataInMem_lo_181};
  wire [95:0]      dataInMem_hi_hi_lo_lo_hi_5 = {dataInMem_hi_248, dataInMem_lo_184, dataInMem_hi_247, dataInMem_lo_183};
  wire [191:0]     dataInMem_hi_hi_lo_lo_5 = {dataInMem_hi_hi_lo_lo_hi_5, dataInMem_hi_hi_lo_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_lo_hi_lo_5 = {dataInMem_hi_250, dataInMem_lo_186, dataInMem_hi_249, dataInMem_lo_185};
  wire [95:0]      dataInMem_hi_hi_lo_hi_hi_5 = {dataInMem_hi_252, dataInMem_lo_188, dataInMem_hi_251, dataInMem_lo_187};
  wire [191:0]     dataInMem_hi_hi_lo_hi_5 = {dataInMem_hi_hi_lo_hi_hi_5, dataInMem_hi_hi_lo_hi_lo_5};
  wire [383:0]     dataInMem_hi_hi_lo_5 = {dataInMem_hi_hi_lo_hi_5, dataInMem_hi_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_hi_lo_lo_5 = {dataInMem_hi_254, dataInMem_lo_190, dataInMem_hi_253, dataInMem_lo_189};
  wire [95:0]      dataInMem_hi_hi_hi_lo_hi_5 = {dataInMem_hi_256, dataInMem_lo_192, dataInMem_hi_255, dataInMem_lo_191};
  wire [191:0]     dataInMem_hi_hi_hi_lo_5 = {dataInMem_hi_hi_hi_lo_hi_5, dataInMem_hi_hi_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_hi_hi_lo_5 = {dataInMem_hi_258, dataInMem_lo_194, dataInMem_hi_257, dataInMem_lo_193};
  wire [95:0]      dataInMem_hi_hi_hi_hi_hi_5 = {dataInMem_hi_260, dataInMem_lo_196, dataInMem_hi_259, dataInMem_lo_195};
  wire [191:0]     dataInMem_hi_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_hi_lo_5};
  wire [383:0]     dataInMem_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_lo_5};
  wire [767:0]     dataInMem_hi_hi_133 = {dataInMem_hi_hi_hi_5, dataInMem_hi_hi_lo_5};
  wire [1535:0]    dataInMem_hi_261 = {dataInMem_hi_hi_133, dataInMem_hi_lo_5};
  wire [3071:0]    dataInMem_5 = {dataInMem_hi_261, dataInMem_lo_197};
  wire [511:0]     regroupCacheLine_5_0 = dataInMem_5[511:0];
  wire [511:0]     regroupCacheLine_5_1 = dataInMem_5[1023:512];
  wire [511:0]     regroupCacheLine_5_2 = dataInMem_5[1535:1024];
  wire [511:0]     regroupCacheLine_5_3 = dataInMem_5[2047:1536];
  wire [511:0]     regroupCacheLine_5_4 = dataInMem_5[2559:2048];
  wire [511:0]     regroupCacheLine_5_5 = dataInMem_5[3071:2560];
  wire [511:0]     res_40 = regroupCacheLine_5_0;
  wire [511:0]     res_41 = regroupCacheLine_5_1;
  wire [511:0]     res_42 = regroupCacheLine_5_2;
  wire [511:0]     res_43 = regroupCacheLine_5_3;
  wire [511:0]     res_44 = regroupCacheLine_5_4;
  wire [511:0]     res_45 = regroupCacheLine_5_5;
  wire [1023:0]    lo_lo_5 = {res_41, res_40};
  wire [1023:0]    lo_hi_5 = {res_43, res_42};
  wire [2047:0]    lo_5 = {lo_hi_5, lo_lo_5};
  wire [1023:0]    hi_lo_5 = {res_45, res_44};
  wire [2047:0]    hi_5 = {1024'h0, hi_lo_5};
  wire [4095:0]    regroupLoadData_0_5 = {hi_5, lo_5};
  wire [23:0]      dataInMem_lo_198 = {dataInMem_lo_hi_70, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_hi_hi_134 = {dataRegroupBySew_6_0, dataRegroupBySew_5_0};
  wire [31:0]      dataInMem_hi_262 = {dataInMem_hi_hi_134, dataInMem_hi_lo_6};
  wire [23:0]      dataInMem_lo_199 = {dataInMem_lo_hi_71, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_hi_hi_135 = {dataRegroupBySew_6_1, dataRegroupBySew_5_1};
  wire [31:0]      dataInMem_hi_263 = {dataInMem_hi_hi_135, dataInMem_hi_lo_7};
  wire [23:0]      dataInMem_lo_200 = {dataInMem_lo_hi_72, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_hi_hi_136 = {dataRegroupBySew_6_2, dataRegroupBySew_5_2};
  wire [31:0]      dataInMem_hi_264 = {dataInMem_hi_hi_136, dataInMem_hi_lo_8};
  wire [23:0]      dataInMem_lo_201 = {dataInMem_lo_hi_73, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_hi_hi_137 = {dataRegroupBySew_6_3, dataRegroupBySew_5_3};
  wire [31:0]      dataInMem_hi_265 = {dataInMem_hi_hi_137, dataInMem_hi_lo_9};
  wire [23:0]      dataInMem_lo_202 = {dataInMem_lo_hi_74, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_hi_hi_138 = {dataRegroupBySew_6_4, dataRegroupBySew_5_4};
  wire [31:0]      dataInMem_hi_266 = {dataInMem_hi_hi_138, dataInMem_hi_lo_10};
  wire [23:0]      dataInMem_lo_203 = {dataInMem_lo_hi_75, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_hi_hi_139 = {dataRegroupBySew_6_5, dataRegroupBySew_5_5};
  wire [31:0]      dataInMem_hi_267 = {dataInMem_hi_hi_139, dataInMem_hi_lo_11};
  wire [23:0]      dataInMem_lo_204 = {dataInMem_lo_hi_76, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_hi_hi_140 = {dataRegroupBySew_6_6, dataRegroupBySew_5_6};
  wire [31:0]      dataInMem_hi_268 = {dataInMem_hi_hi_140, dataInMem_hi_lo_12};
  wire [23:0]      dataInMem_lo_205 = {dataInMem_lo_hi_77, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_hi_hi_141 = {dataRegroupBySew_6_7, dataRegroupBySew_5_7};
  wire [31:0]      dataInMem_hi_269 = {dataInMem_hi_hi_141, dataInMem_hi_lo_13};
  wire [23:0]      dataInMem_lo_206 = {dataInMem_lo_hi_78, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_hi_hi_142 = {dataRegroupBySew_6_8, dataRegroupBySew_5_8};
  wire [31:0]      dataInMem_hi_270 = {dataInMem_hi_hi_142, dataInMem_hi_lo_14};
  wire [23:0]      dataInMem_lo_207 = {dataInMem_lo_hi_79, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_hi_hi_143 = {dataRegroupBySew_6_9, dataRegroupBySew_5_9};
  wire [31:0]      dataInMem_hi_271 = {dataInMem_hi_hi_143, dataInMem_hi_lo_15};
  wire [23:0]      dataInMem_lo_208 = {dataInMem_lo_hi_80, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_hi_hi_144 = {dataRegroupBySew_6_10, dataRegroupBySew_5_10};
  wire [31:0]      dataInMem_hi_272 = {dataInMem_hi_hi_144, dataInMem_hi_lo_16};
  wire [23:0]      dataInMem_lo_209 = {dataInMem_lo_hi_81, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_hi_hi_145 = {dataRegroupBySew_6_11, dataRegroupBySew_5_11};
  wire [31:0]      dataInMem_hi_273 = {dataInMem_hi_hi_145, dataInMem_hi_lo_17};
  wire [23:0]      dataInMem_lo_210 = {dataInMem_lo_hi_82, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_hi_hi_146 = {dataRegroupBySew_6_12, dataRegroupBySew_5_12};
  wire [31:0]      dataInMem_hi_274 = {dataInMem_hi_hi_146, dataInMem_hi_lo_18};
  wire [23:0]      dataInMem_lo_211 = {dataInMem_lo_hi_83, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_hi_hi_147 = {dataRegroupBySew_6_13, dataRegroupBySew_5_13};
  wire [31:0]      dataInMem_hi_275 = {dataInMem_hi_hi_147, dataInMem_hi_lo_19};
  wire [23:0]      dataInMem_lo_212 = {dataInMem_lo_hi_84, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_hi_hi_148 = {dataRegroupBySew_6_14, dataRegroupBySew_5_14};
  wire [31:0]      dataInMem_hi_276 = {dataInMem_hi_hi_148, dataInMem_hi_lo_20};
  wire [23:0]      dataInMem_lo_213 = {dataInMem_lo_hi_85, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_hi_hi_149 = {dataRegroupBySew_6_15, dataRegroupBySew_5_15};
  wire [31:0]      dataInMem_hi_277 = {dataInMem_hi_hi_149, dataInMem_hi_lo_21};
  wire [23:0]      dataInMem_lo_214 = {dataInMem_lo_hi_86, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_hi_hi_150 = {dataRegroupBySew_6_16, dataRegroupBySew_5_16};
  wire [31:0]      dataInMem_hi_278 = {dataInMem_hi_hi_150, dataInMem_hi_lo_22};
  wire [23:0]      dataInMem_lo_215 = {dataInMem_lo_hi_87, dataRegroupBySew_0_17};
  wire [15:0]      dataInMem_hi_hi_151 = {dataRegroupBySew_6_17, dataRegroupBySew_5_17};
  wire [31:0]      dataInMem_hi_279 = {dataInMem_hi_hi_151, dataInMem_hi_lo_23};
  wire [23:0]      dataInMem_lo_216 = {dataInMem_lo_hi_88, dataRegroupBySew_0_18};
  wire [15:0]      dataInMem_hi_hi_152 = {dataRegroupBySew_6_18, dataRegroupBySew_5_18};
  wire [31:0]      dataInMem_hi_280 = {dataInMem_hi_hi_152, dataInMem_hi_lo_24};
  wire [23:0]      dataInMem_lo_217 = {dataInMem_lo_hi_89, dataRegroupBySew_0_19};
  wire [15:0]      dataInMem_hi_hi_153 = {dataRegroupBySew_6_19, dataRegroupBySew_5_19};
  wire [31:0]      dataInMem_hi_281 = {dataInMem_hi_hi_153, dataInMem_hi_lo_25};
  wire [23:0]      dataInMem_lo_218 = {dataInMem_lo_hi_90, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_hi_hi_154 = {dataRegroupBySew_6_20, dataRegroupBySew_5_20};
  wire [31:0]      dataInMem_hi_282 = {dataInMem_hi_hi_154, dataInMem_hi_lo_26};
  wire [23:0]      dataInMem_lo_219 = {dataInMem_lo_hi_91, dataRegroupBySew_0_21};
  wire [15:0]      dataInMem_hi_hi_155 = {dataRegroupBySew_6_21, dataRegroupBySew_5_21};
  wire [31:0]      dataInMem_hi_283 = {dataInMem_hi_hi_155, dataInMem_hi_lo_27};
  wire [23:0]      dataInMem_lo_220 = {dataInMem_lo_hi_92, dataRegroupBySew_0_22};
  wire [15:0]      dataInMem_hi_hi_156 = {dataRegroupBySew_6_22, dataRegroupBySew_5_22};
  wire [31:0]      dataInMem_hi_284 = {dataInMem_hi_hi_156, dataInMem_hi_lo_28};
  wire [23:0]      dataInMem_lo_221 = {dataInMem_lo_hi_93, dataRegroupBySew_0_23};
  wire [15:0]      dataInMem_hi_hi_157 = {dataRegroupBySew_6_23, dataRegroupBySew_5_23};
  wire [31:0]      dataInMem_hi_285 = {dataInMem_hi_hi_157, dataInMem_hi_lo_29};
  wire [23:0]      dataInMem_lo_222 = {dataInMem_lo_hi_94, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_hi_hi_158 = {dataRegroupBySew_6_24, dataRegroupBySew_5_24};
  wire [31:0]      dataInMem_hi_286 = {dataInMem_hi_hi_158, dataInMem_hi_lo_30};
  wire [23:0]      dataInMem_lo_223 = {dataInMem_lo_hi_95, dataRegroupBySew_0_25};
  wire [15:0]      dataInMem_hi_hi_159 = {dataRegroupBySew_6_25, dataRegroupBySew_5_25};
  wire [31:0]      dataInMem_hi_287 = {dataInMem_hi_hi_159, dataInMem_hi_lo_31};
  wire [23:0]      dataInMem_lo_224 = {dataInMem_lo_hi_96, dataRegroupBySew_0_26};
  wire [15:0]      dataInMem_hi_hi_160 = {dataRegroupBySew_6_26, dataRegroupBySew_5_26};
  wire [31:0]      dataInMem_hi_288 = {dataInMem_hi_hi_160, dataInMem_hi_lo_32};
  wire [23:0]      dataInMem_lo_225 = {dataInMem_lo_hi_97, dataRegroupBySew_0_27};
  wire [15:0]      dataInMem_hi_hi_161 = {dataRegroupBySew_6_27, dataRegroupBySew_5_27};
  wire [31:0]      dataInMem_hi_289 = {dataInMem_hi_hi_161, dataInMem_hi_lo_33};
  wire [23:0]      dataInMem_lo_226 = {dataInMem_lo_hi_98, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_hi_hi_162 = {dataRegroupBySew_6_28, dataRegroupBySew_5_28};
  wire [31:0]      dataInMem_hi_290 = {dataInMem_hi_hi_162, dataInMem_hi_lo_34};
  wire [23:0]      dataInMem_lo_227 = {dataInMem_lo_hi_99, dataRegroupBySew_0_29};
  wire [15:0]      dataInMem_hi_hi_163 = {dataRegroupBySew_6_29, dataRegroupBySew_5_29};
  wire [31:0]      dataInMem_hi_291 = {dataInMem_hi_hi_163, dataInMem_hi_lo_35};
  wire [23:0]      dataInMem_lo_228 = {dataInMem_lo_hi_100, dataRegroupBySew_0_30};
  wire [15:0]      dataInMem_hi_hi_164 = {dataRegroupBySew_6_30, dataRegroupBySew_5_30};
  wire [31:0]      dataInMem_hi_292 = {dataInMem_hi_hi_164, dataInMem_hi_lo_36};
  wire [23:0]      dataInMem_lo_229 = {dataInMem_lo_hi_101, dataRegroupBySew_0_31};
  wire [15:0]      dataInMem_hi_hi_165 = {dataRegroupBySew_6_31, dataRegroupBySew_5_31};
  wire [31:0]      dataInMem_hi_293 = {dataInMem_hi_hi_165, dataInMem_hi_lo_37};
  wire [23:0]      dataInMem_lo_230 = {dataInMem_lo_hi_102, dataRegroupBySew_0_32};
  wire [15:0]      dataInMem_hi_hi_166 = {dataRegroupBySew_6_32, dataRegroupBySew_5_32};
  wire [31:0]      dataInMem_hi_294 = {dataInMem_hi_hi_166, dataInMem_hi_lo_38};
  wire [23:0]      dataInMem_lo_231 = {dataInMem_lo_hi_103, dataRegroupBySew_0_33};
  wire [15:0]      dataInMem_hi_hi_167 = {dataRegroupBySew_6_33, dataRegroupBySew_5_33};
  wire [31:0]      dataInMem_hi_295 = {dataInMem_hi_hi_167, dataInMem_hi_lo_39};
  wire [23:0]      dataInMem_lo_232 = {dataInMem_lo_hi_104, dataRegroupBySew_0_34};
  wire [15:0]      dataInMem_hi_hi_168 = {dataRegroupBySew_6_34, dataRegroupBySew_5_34};
  wire [31:0]      dataInMem_hi_296 = {dataInMem_hi_hi_168, dataInMem_hi_lo_40};
  wire [23:0]      dataInMem_lo_233 = {dataInMem_lo_hi_105, dataRegroupBySew_0_35};
  wire [15:0]      dataInMem_hi_hi_169 = {dataRegroupBySew_6_35, dataRegroupBySew_5_35};
  wire [31:0]      dataInMem_hi_297 = {dataInMem_hi_hi_169, dataInMem_hi_lo_41};
  wire [23:0]      dataInMem_lo_234 = {dataInMem_lo_hi_106, dataRegroupBySew_0_36};
  wire [15:0]      dataInMem_hi_hi_170 = {dataRegroupBySew_6_36, dataRegroupBySew_5_36};
  wire [31:0]      dataInMem_hi_298 = {dataInMem_hi_hi_170, dataInMem_hi_lo_42};
  wire [23:0]      dataInMem_lo_235 = {dataInMem_lo_hi_107, dataRegroupBySew_0_37};
  wire [15:0]      dataInMem_hi_hi_171 = {dataRegroupBySew_6_37, dataRegroupBySew_5_37};
  wire [31:0]      dataInMem_hi_299 = {dataInMem_hi_hi_171, dataInMem_hi_lo_43};
  wire [23:0]      dataInMem_lo_236 = {dataInMem_lo_hi_108, dataRegroupBySew_0_38};
  wire [15:0]      dataInMem_hi_hi_172 = {dataRegroupBySew_6_38, dataRegroupBySew_5_38};
  wire [31:0]      dataInMem_hi_300 = {dataInMem_hi_hi_172, dataInMem_hi_lo_44};
  wire [23:0]      dataInMem_lo_237 = {dataInMem_lo_hi_109, dataRegroupBySew_0_39};
  wire [15:0]      dataInMem_hi_hi_173 = {dataRegroupBySew_6_39, dataRegroupBySew_5_39};
  wire [31:0]      dataInMem_hi_301 = {dataInMem_hi_hi_173, dataInMem_hi_lo_45};
  wire [23:0]      dataInMem_lo_238 = {dataInMem_lo_hi_110, dataRegroupBySew_0_40};
  wire [15:0]      dataInMem_hi_hi_174 = {dataRegroupBySew_6_40, dataRegroupBySew_5_40};
  wire [31:0]      dataInMem_hi_302 = {dataInMem_hi_hi_174, dataInMem_hi_lo_46};
  wire [23:0]      dataInMem_lo_239 = {dataInMem_lo_hi_111, dataRegroupBySew_0_41};
  wire [15:0]      dataInMem_hi_hi_175 = {dataRegroupBySew_6_41, dataRegroupBySew_5_41};
  wire [31:0]      dataInMem_hi_303 = {dataInMem_hi_hi_175, dataInMem_hi_lo_47};
  wire [23:0]      dataInMem_lo_240 = {dataInMem_lo_hi_112, dataRegroupBySew_0_42};
  wire [15:0]      dataInMem_hi_hi_176 = {dataRegroupBySew_6_42, dataRegroupBySew_5_42};
  wire [31:0]      dataInMem_hi_304 = {dataInMem_hi_hi_176, dataInMem_hi_lo_48};
  wire [23:0]      dataInMem_lo_241 = {dataInMem_lo_hi_113, dataRegroupBySew_0_43};
  wire [15:0]      dataInMem_hi_hi_177 = {dataRegroupBySew_6_43, dataRegroupBySew_5_43};
  wire [31:0]      dataInMem_hi_305 = {dataInMem_hi_hi_177, dataInMem_hi_lo_49};
  wire [23:0]      dataInMem_lo_242 = {dataInMem_lo_hi_114, dataRegroupBySew_0_44};
  wire [15:0]      dataInMem_hi_hi_178 = {dataRegroupBySew_6_44, dataRegroupBySew_5_44};
  wire [31:0]      dataInMem_hi_306 = {dataInMem_hi_hi_178, dataInMem_hi_lo_50};
  wire [23:0]      dataInMem_lo_243 = {dataInMem_lo_hi_115, dataRegroupBySew_0_45};
  wire [15:0]      dataInMem_hi_hi_179 = {dataRegroupBySew_6_45, dataRegroupBySew_5_45};
  wire [31:0]      dataInMem_hi_307 = {dataInMem_hi_hi_179, dataInMem_hi_lo_51};
  wire [23:0]      dataInMem_lo_244 = {dataInMem_lo_hi_116, dataRegroupBySew_0_46};
  wire [15:0]      dataInMem_hi_hi_180 = {dataRegroupBySew_6_46, dataRegroupBySew_5_46};
  wire [31:0]      dataInMem_hi_308 = {dataInMem_hi_hi_180, dataInMem_hi_lo_52};
  wire [23:0]      dataInMem_lo_245 = {dataInMem_lo_hi_117, dataRegroupBySew_0_47};
  wire [15:0]      dataInMem_hi_hi_181 = {dataRegroupBySew_6_47, dataRegroupBySew_5_47};
  wire [31:0]      dataInMem_hi_309 = {dataInMem_hi_hi_181, dataInMem_hi_lo_53};
  wire [23:0]      dataInMem_lo_246 = {dataInMem_lo_hi_118, dataRegroupBySew_0_48};
  wire [15:0]      dataInMem_hi_hi_182 = {dataRegroupBySew_6_48, dataRegroupBySew_5_48};
  wire [31:0]      dataInMem_hi_310 = {dataInMem_hi_hi_182, dataInMem_hi_lo_54};
  wire [23:0]      dataInMem_lo_247 = {dataInMem_lo_hi_119, dataRegroupBySew_0_49};
  wire [15:0]      dataInMem_hi_hi_183 = {dataRegroupBySew_6_49, dataRegroupBySew_5_49};
  wire [31:0]      dataInMem_hi_311 = {dataInMem_hi_hi_183, dataInMem_hi_lo_55};
  wire [23:0]      dataInMem_lo_248 = {dataInMem_lo_hi_120, dataRegroupBySew_0_50};
  wire [15:0]      dataInMem_hi_hi_184 = {dataRegroupBySew_6_50, dataRegroupBySew_5_50};
  wire [31:0]      dataInMem_hi_312 = {dataInMem_hi_hi_184, dataInMem_hi_lo_56};
  wire [23:0]      dataInMem_lo_249 = {dataInMem_lo_hi_121, dataRegroupBySew_0_51};
  wire [15:0]      dataInMem_hi_hi_185 = {dataRegroupBySew_6_51, dataRegroupBySew_5_51};
  wire [31:0]      dataInMem_hi_313 = {dataInMem_hi_hi_185, dataInMem_hi_lo_57};
  wire [23:0]      dataInMem_lo_250 = {dataInMem_lo_hi_122, dataRegroupBySew_0_52};
  wire [15:0]      dataInMem_hi_hi_186 = {dataRegroupBySew_6_52, dataRegroupBySew_5_52};
  wire [31:0]      dataInMem_hi_314 = {dataInMem_hi_hi_186, dataInMem_hi_lo_58};
  wire [23:0]      dataInMem_lo_251 = {dataInMem_lo_hi_123, dataRegroupBySew_0_53};
  wire [15:0]      dataInMem_hi_hi_187 = {dataRegroupBySew_6_53, dataRegroupBySew_5_53};
  wire [31:0]      dataInMem_hi_315 = {dataInMem_hi_hi_187, dataInMem_hi_lo_59};
  wire [23:0]      dataInMem_lo_252 = {dataInMem_lo_hi_124, dataRegroupBySew_0_54};
  wire [15:0]      dataInMem_hi_hi_188 = {dataRegroupBySew_6_54, dataRegroupBySew_5_54};
  wire [31:0]      dataInMem_hi_316 = {dataInMem_hi_hi_188, dataInMem_hi_lo_60};
  wire [23:0]      dataInMem_lo_253 = {dataInMem_lo_hi_125, dataRegroupBySew_0_55};
  wire [15:0]      dataInMem_hi_hi_189 = {dataRegroupBySew_6_55, dataRegroupBySew_5_55};
  wire [31:0]      dataInMem_hi_317 = {dataInMem_hi_hi_189, dataInMem_hi_lo_61};
  wire [23:0]      dataInMem_lo_254 = {dataInMem_lo_hi_126, dataRegroupBySew_0_56};
  wire [15:0]      dataInMem_hi_hi_190 = {dataRegroupBySew_6_56, dataRegroupBySew_5_56};
  wire [31:0]      dataInMem_hi_318 = {dataInMem_hi_hi_190, dataInMem_hi_lo_62};
  wire [23:0]      dataInMem_lo_255 = {dataInMem_lo_hi_127, dataRegroupBySew_0_57};
  wire [15:0]      dataInMem_hi_hi_191 = {dataRegroupBySew_6_57, dataRegroupBySew_5_57};
  wire [31:0]      dataInMem_hi_319 = {dataInMem_hi_hi_191, dataInMem_hi_lo_63};
  wire [23:0]      dataInMem_lo_256 = {dataInMem_lo_hi_128, dataRegroupBySew_0_58};
  wire [15:0]      dataInMem_hi_hi_192 = {dataRegroupBySew_6_58, dataRegroupBySew_5_58};
  wire [31:0]      dataInMem_hi_320 = {dataInMem_hi_hi_192, dataInMem_hi_lo_64};
  wire [23:0]      dataInMem_lo_257 = {dataInMem_lo_hi_129, dataRegroupBySew_0_59};
  wire [15:0]      dataInMem_hi_hi_193 = {dataRegroupBySew_6_59, dataRegroupBySew_5_59};
  wire [31:0]      dataInMem_hi_321 = {dataInMem_hi_hi_193, dataInMem_hi_lo_65};
  wire [23:0]      dataInMem_lo_258 = {dataInMem_lo_hi_130, dataRegroupBySew_0_60};
  wire [15:0]      dataInMem_hi_hi_194 = {dataRegroupBySew_6_60, dataRegroupBySew_5_60};
  wire [31:0]      dataInMem_hi_322 = {dataInMem_hi_hi_194, dataInMem_hi_lo_66};
  wire [23:0]      dataInMem_lo_259 = {dataInMem_lo_hi_131, dataRegroupBySew_0_61};
  wire [15:0]      dataInMem_hi_hi_195 = {dataRegroupBySew_6_61, dataRegroupBySew_5_61};
  wire [31:0]      dataInMem_hi_323 = {dataInMem_hi_hi_195, dataInMem_hi_lo_67};
  wire [23:0]      dataInMem_lo_260 = {dataInMem_lo_hi_132, dataRegroupBySew_0_62};
  wire [15:0]      dataInMem_hi_hi_196 = {dataRegroupBySew_6_62, dataRegroupBySew_5_62};
  wire [31:0]      dataInMem_hi_324 = {dataInMem_hi_hi_196, dataInMem_hi_lo_68};
  wire [23:0]      dataInMem_lo_261 = {dataInMem_lo_hi_133, dataRegroupBySew_0_63};
  wire [15:0]      dataInMem_hi_hi_197 = {dataRegroupBySew_6_63, dataRegroupBySew_5_63};
  wire [31:0]      dataInMem_hi_325 = {dataInMem_hi_hi_197, dataInMem_hi_lo_69};
  wire [111:0]     dataInMem_lo_lo_lo_lo_lo_6 = {dataInMem_hi_263, dataInMem_lo_199, dataInMem_hi_262, dataInMem_lo_198};
  wire [111:0]     dataInMem_lo_lo_lo_lo_hi_6 = {dataInMem_hi_265, dataInMem_lo_201, dataInMem_hi_264, dataInMem_lo_200};
  wire [223:0]     dataInMem_lo_lo_lo_lo_6 = {dataInMem_lo_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_lo_lo_hi_lo_6 = {dataInMem_hi_267, dataInMem_lo_203, dataInMem_hi_266, dataInMem_lo_202};
  wire [111:0]     dataInMem_lo_lo_lo_hi_hi_6 = {dataInMem_hi_269, dataInMem_lo_205, dataInMem_hi_268, dataInMem_lo_204};
  wire [223:0]     dataInMem_lo_lo_lo_hi_6 = {dataInMem_lo_lo_lo_hi_hi_6, dataInMem_lo_lo_lo_hi_lo_6};
  wire [447:0]     dataInMem_lo_lo_lo_6 = {dataInMem_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_lo_hi_lo_lo_6 = {dataInMem_hi_271, dataInMem_lo_207, dataInMem_hi_270, dataInMem_lo_206};
  wire [111:0]     dataInMem_lo_lo_hi_lo_hi_6 = {dataInMem_hi_273, dataInMem_lo_209, dataInMem_hi_272, dataInMem_lo_208};
  wire [223:0]     dataInMem_lo_lo_hi_lo_6 = {dataInMem_lo_lo_hi_lo_hi_6, dataInMem_lo_lo_hi_lo_lo_6};
  wire [111:0]     dataInMem_lo_lo_hi_hi_lo_6 = {dataInMem_hi_275, dataInMem_lo_211, dataInMem_hi_274, dataInMem_lo_210};
  wire [111:0]     dataInMem_lo_lo_hi_hi_hi_6 = {dataInMem_hi_277, dataInMem_lo_213, dataInMem_hi_276, dataInMem_lo_212};
  wire [223:0]     dataInMem_lo_lo_hi_hi_6 = {dataInMem_lo_lo_hi_hi_hi_6, dataInMem_lo_lo_hi_hi_lo_6};
  wire [447:0]     dataInMem_lo_lo_hi_6 = {dataInMem_lo_lo_hi_hi_6, dataInMem_lo_lo_hi_lo_6};
  wire [895:0]     dataInMem_lo_lo_6 = {dataInMem_lo_lo_hi_6, dataInMem_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_lo_lo_lo_6 = {dataInMem_hi_279, dataInMem_lo_215, dataInMem_hi_278, dataInMem_lo_214};
  wire [111:0]     dataInMem_lo_hi_lo_lo_hi_6 = {dataInMem_hi_281, dataInMem_lo_217, dataInMem_hi_280, dataInMem_lo_216};
  wire [223:0]     dataInMem_lo_hi_lo_lo_6 = {dataInMem_lo_hi_lo_lo_hi_6, dataInMem_lo_hi_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_lo_hi_lo_6 = {dataInMem_hi_283, dataInMem_lo_219, dataInMem_hi_282, dataInMem_lo_218};
  wire [111:0]     dataInMem_lo_hi_lo_hi_hi_6 = {dataInMem_hi_285, dataInMem_lo_221, dataInMem_hi_284, dataInMem_lo_220};
  wire [223:0]     dataInMem_lo_hi_lo_hi_6 = {dataInMem_lo_hi_lo_hi_hi_6, dataInMem_lo_hi_lo_hi_lo_6};
  wire [447:0]     dataInMem_lo_hi_lo_6 = {dataInMem_lo_hi_lo_hi_6, dataInMem_lo_hi_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_hi_lo_lo_6 = {dataInMem_hi_287, dataInMem_lo_223, dataInMem_hi_286, dataInMem_lo_222};
  wire [111:0]     dataInMem_lo_hi_hi_lo_hi_6 = {dataInMem_hi_289, dataInMem_lo_225, dataInMem_hi_288, dataInMem_lo_224};
  wire [223:0]     dataInMem_lo_hi_hi_lo_6 = {dataInMem_lo_hi_hi_lo_hi_6, dataInMem_lo_hi_hi_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_hi_hi_lo_6 = {dataInMem_hi_291, dataInMem_lo_227, dataInMem_hi_290, dataInMem_lo_226};
  wire [111:0]     dataInMem_lo_hi_hi_hi_hi_6 = {dataInMem_hi_293, dataInMem_lo_229, dataInMem_hi_292, dataInMem_lo_228};
  wire [223:0]     dataInMem_lo_hi_hi_hi_6 = {dataInMem_lo_hi_hi_hi_hi_6, dataInMem_lo_hi_hi_hi_lo_6};
  wire [447:0]     dataInMem_lo_hi_hi_6 = {dataInMem_lo_hi_hi_hi_6, dataInMem_lo_hi_hi_lo_6};
  wire [895:0]     dataInMem_lo_hi_134 = {dataInMem_lo_hi_hi_6, dataInMem_lo_hi_lo_6};
  wire [1791:0]    dataInMem_lo_262 = {dataInMem_lo_hi_134, dataInMem_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_lo_lo_lo_6 = {dataInMem_hi_295, dataInMem_lo_231, dataInMem_hi_294, dataInMem_lo_230};
  wire [111:0]     dataInMem_hi_lo_lo_lo_hi_6 = {dataInMem_hi_297, dataInMem_lo_233, dataInMem_hi_296, dataInMem_lo_232};
  wire [223:0]     dataInMem_hi_lo_lo_lo_6 = {dataInMem_hi_lo_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_lo_hi_lo_6 = {dataInMem_hi_299, dataInMem_lo_235, dataInMem_hi_298, dataInMem_lo_234};
  wire [111:0]     dataInMem_hi_lo_lo_hi_hi_6 = {dataInMem_hi_301, dataInMem_lo_237, dataInMem_hi_300, dataInMem_lo_236};
  wire [223:0]     dataInMem_hi_lo_lo_hi_6 = {dataInMem_hi_lo_lo_hi_hi_6, dataInMem_hi_lo_lo_hi_lo_6};
  wire [447:0]     dataInMem_hi_lo_lo_6 = {dataInMem_hi_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_hi_lo_lo_6 = {dataInMem_hi_303, dataInMem_lo_239, dataInMem_hi_302, dataInMem_lo_238};
  wire [111:0]     dataInMem_hi_lo_hi_lo_hi_6 = {dataInMem_hi_305, dataInMem_lo_241, dataInMem_hi_304, dataInMem_lo_240};
  wire [223:0]     dataInMem_hi_lo_hi_lo_6 = {dataInMem_hi_lo_hi_lo_hi_6, dataInMem_hi_lo_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_hi_hi_lo_6 = {dataInMem_hi_307, dataInMem_lo_243, dataInMem_hi_306, dataInMem_lo_242};
  wire [111:0]     dataInMem_hi_lo_hi_hi_hi_6 = {dataInMem_hi_309, dataInMem_lo_245, dataInMem_hi_308, dataInMem_lo_244};
  wire [223:0]     dataInMem_hi_lo_hi_hi_6 = {dataInMem_hi_lo_hi_hi_hi_6, dataInMem_hi_lo_hi_hi_lo_6};
  wire [447:0]     dataInMem_hi_lo_hi_6 = {dataInMem_hi_lo_hi_hi_6, dataInMem_hi_lo_hi_lo_6};
  wire [895:0]     dataInMem_hi_lo_70 = {dataInMem_hi_lo_hi_6, dataInMem_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_lo_lo_lo_6 = {dataInMem_hi_311, dataInMem_lo_247, dataInMem_hi_310, dataInMem_lo_246};
  wire [111:0]     dataInMem_hi_hi_lo_lo_hi_6 = {dataInMem_hi_313, dataInMem_lo_249, dataInMem_hi_312, dataInMem_lo_248};
  wire [223:0]     dataInMem_hi_hi_lo_lo_6 = {dataInMem_hi_hi_lo_lo_hi_6, dataInMem_hi_hi_lo_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_lo_hi_lo_6 = {dataInMem_hi_315, dataInMem_lo_251, dataInMem_hi_314, dataInMem_lo_250};
  wire [111:0]     dataInMem_hi_hi_lo_hi_hi_6 = {dataInMem_hi_317, dataInMem_lo_253, dataInMem_hi_316, dataInMem_lo_252};
  wire [223:0]     dataInMem_hi_hi_lo_hi_6 = {dataInMem_hi_hi_lo_hi_hi_6, dataInMem_hi_hi_lo_hi_lo_6};
  wire [447:0]     dataInMem_hi_hi_lo_6 = {dataInMem_hi_hi_lo_hi_6, dataInMem_hi_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_hi_lo_lo_6 = {dataInMem_hi_319, dataInMem_lo_255, dataInMem_hi_318, dataInMem_lo_254};
  wire [111:0]     dataInMem_hi_hi_hi_lo_hi_6 = {dataInMem_hi_321, dataInMem_lo_257, dataInMem_hi_320, dataInMem_lo_256};
  wire [223:0]     dataInMem_hi_hi_hi_lo_6 = {dataInMem_hi_hi_hi_lo_hi_6, dataInMem_hi_hi_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_hi_hi_lo_6 = {dataInMem_hi_323, dataInMem_lo_259, dataInMem_hi_322, dataInMem_lo_258};
  wire [111:0]     dataInMem_hi_hi_hi_hi_hi_6 = {dataInMem_hi_325, dataInMem_lo_261, dataInMem_hi_324, dataInMem_lo_260};
  wire [223:0]     dataInMem_hi_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_hi_lo_6};
  wire [447:0]     dataInMem_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_lo_6};
  wire [895:0]     dataInMem_hi_hi_198 = {dataInMem_hi_hi_hi_6, dataInMem_hi_hi_lo_6};
  wire [1791:0]    dataInMem_hi_326 = {dataInMem_hi_hi_198, dataInMem_hi_lo_70};
  wire [3583:0]    dataInMem_6 = {dataInMem_hi_326, dataInMem_lo_262};
  wire [511:0]     regroupCacheLine_6_0 = dataInMem_6[511:0];
  wire [511:0]     regroupCacheLine_6_1 = dataInMem_6[1023:512];
  wire [511:0]     regroupCacheLine_6_2 = dataInMem_6[1535:1024];
  wire [511:0]     regroupCacheLine_6_3 = dataInMem_6[2047:1536];
  wire [511:0]     regroupCacheLine_6_4 = dataInMem_6[2559:2048];
  wire [511:0]     regroupCacheLine_6_5 = dataInMem_6[3071:2560];
  wire [511:0]     regroupCacheLine_6_6 = dataInMem_6[3583:3072];
  wire [511:0]     res_48 = regroupCacheLine_6_0;
  wire [511:0]     res_49 = regroupCacheLine_6_1;
  wire [511:0]     res_50 = regroupCacheLine_6_2;
  wire [511:0]     res_51 = regroupCacheLine_6_3;
  wire [511:0]     res_52 = regroupCacheLine_6_4;
  wire [511:0]     res_53 = regroupCacheLine_6_5;
  wire [511:0]     res_54 = regroupCacheLine_6_6;
  wire [1023:0]    lo_lo_6 = {res_49, res_48};
  wire [1023:0]    lo_hi_6 = {res_51, res_50};
  wire [2047:0]    lo_6 = {lo_hi_6, lo_lo_6};
  wire [1023:0]    hi_lo_6 = {res_53, res_52};
  wire [1023:0]    hi_hi_6 = {512'h0, res_54};
  wire [2047:0]    hi_6 = {hi_hi_6, hi_lo_6};
  wire [4095:0]    regroupLoadData_0_6 = {hi_6, lo_6};
  wire [31:0]      dataInMem_lo_263 = {dataInMem_lo_hi_135, dataInMem_lo_lo_7};
  wire [15:0]      dataInMem_hi_hi_199 = {dataRegroupBySew_7_0, dataRegroupBySew_6_0};
  wire [31:0]      dataInMem_hi_327 = {dataInMem_hi_hi_199, dataInMem_hi_lo_71};
  wire [31:0]      dataInMem_lo_264 = {dataInMem_lo_hi_136, dataInMem_lo_lo_8};
  wire [15:0]      dataInMem_hi_hi_200 = {dataRegroupBySew_7_1, dataRegroupBySew_6_1};
  wire [31:0]      dataInMem_hi_328 = {dataInMem_hi_hi_200, dataInMem_hi_lo_72};
  wire [31:0]      dataInMem_lo_265 = {dataInMem_lo_hi_137, dataInMem_lo_lo_9};
  wire [15:0]      dataInMem_hi_hi_201 = {dataRegroupBySew_7_2, dataRegroupBySew_6_2};
  wire [31:0]      dataInMem_hi_329 = {dataInMem_hi_hi_201, dataInMem_hi_lo_73};
  wire [31:0]      dataInMem_lo_266 = {dataInMem_lo_hi_138, dataInMem_lo_lo_10};
  wire [15:0]      dataInMem_hi_hi_202 = {dataRegroupBySew_7_3, dataRegroupBySew_6_3};
  wire [31:0]      dataInMem_hi_330 = {dataInMem_hi_hi_202, dataInMem_hi_lo_74};
  wire [31:0]      dataInMem_lo_267 = {dataInMem_lo_hi_139, dataInMem_lo_lo_11};
  wire [15:0]      dataInMem_hi_hi_203 = {dataRegroupBySew_7_4, dataRegroupBySew_6_4};
  wire [31:0]      dataInMem_hi_331 = {dataInMem_hi_hi_203, dataInMem_hi_lo_75};
  wire [31:0]      dataInMem_lo_268 = {dataInMem_lo_hi_140, dataInMem_lo_lo_12};
  wire [15:0]      dataInMem_hi_hi_204 = {dataRegroupBySew_7_5, dataRegroupBySew_6_5};
  wire [31:0]      dataInMem_hi_332 = {dataInMem_hi_hi_204, dataInMem_hi_lo_76};
  wire [31:0]      dataInMem_lo_269 = {dataInMem_lo_hi_141, dataInMem_lo_lo_13};
  wire [15:0]      dataInMem_hi_hi_205 = {dataRegroupBySew_7_6, dataRegroupBySew_6_6};
  wire [31:0]      dataInMem_hi_333 = {dataInMem_hi_hi_205, dataInMem_hi_lo_77};
  wire [31:0]      dataInMem_lo_270 = {dataInMem_lo_hi_142, dataInMem_lo_lo_14};
  wire [15:0]      dataInMem_hi_hi_206 = {dataRegroupBySew_7_7, dataRegroupBySew_6_7};
  wire [31:0]      dataInMem_hi_334 = {dataInMem_hi_hi_206, dataInMem_hi_lo_78};
  wire [31:0]      dataInMem_lo_271 = {dataInMem_lo_hi_143, dataInMem_lo_lo_15};
  wire [15:0]      dataInMem_hi_hi_207 = {dataRegroupBySew_7_8, dataRegroupBySew_6_8};
  wire [31:0]      dataInMem_hi_335 = {dataInMem_hi_hi_207, dataInMem_hi_lo_79};
  wire [31:0]      dataInMem_lo_272 = {dataInMem_lo_hi_144, dataInMem_lo_lo_16};
  wire [15:0]      dataInMem_hi_hi_208 = {dataRegroupBySew_7_9, dataRegroupBySew_6_9};
  wire [31:0]      dataInMem_hi_336 = {dataInMem_hi_hi_208, dataInMem_hi_lo_80};
  wire [31:0]      dataInMem_lo_273 = {dataInMem_lo_hi_145, dataInMem_lo_lo_17};
  wire [15:0]      dataInMem_hi_hi_209 = {dataRegroupBySew_7_10, dataRegroupBySew_6_10};
  wire [31:0]      dataInMem_hi_337 = {dataInMem_hi_hi_209, dataInMem_hi_lo_81};
  wire [31:0]      dataInMem_lo_274 = {dataInMem_lo_hi_146, dataInMem_lo_lo_18};
  wire [15:0]      dataInMem_hi_hi_210 = {dataRegroupBySew_7_11, dataRegroupBySew_6_11};
  wire [31:0]      dataInMem_hi_338 = {dataInMem_hi_hi_210, dataInMem_hi_lo_82};
  wire [31:0]      dataInMem_lo_275 = {dataInMem_lo_hi_147, dataInMem_lo_lo_19};
  wire [15:0]      dataInMem_hi_hi_211 = {dataRegroupBySew_7_12, dataRegroupBySew_6_12};
  wire [31:0]      dataInMem_hi_339 = {dataInMem_hi_hi_211, dataInMem_hi_lo_83};
  wire [31:0]      dataInMem_lo_276 = {dataInMem_lo_hi_148, dataInMem_lo_lo_20};
  wire [15:0]      dataInMem_hi_hi_212 = {dataRegroupBySew_7_13, dataRegroupBySew_6_13};
  wire [31:0]      dataInMem_hi_340 = {dataInMem_hi_hi_212, dataInMem_hi_lo_84};
  wire [31:0]      dataInMem_lo_277 = {dataInMem_lo_hi_149, dataInMem_lo_lo_21};
  wire [15:0]      dataInMem_hi_hi_213 = {dataRegroupBySew_7_14, dataRegroupBySew_6_14};
  wire [31:0]      dataInMem_hi_341 = {dataInMem_hi_hi_213, dataInMem_hi_lo_85};
  wire [31:0]      dataInMem_lo_278 = {dataInMem_lo_hi_150, dataInMem_lo_lo_22};
  wire [15:0]      dataInMem_hi_hi_214 = {dataRegroupBySew_7_15, dataRegroupBySew_6_15};
  wire [31:0]      dataInMem_hi_342 = {dataInMem_hi_hi_214, dataInMem_hi_lo_86};
  wire [31:0]      dataInMem_lo_279 = {dataInMem_lo_hi_151, dataInMem_lo_lo_23};
  wire [15:0]      dataInMem_hi_hi_215 = {dataRegroupBySew_7_16, dataRegroupBySew_6_16};
  wire [31:0]      dataInMem_hi_343 = {dataInMem_hi_hi_215, dataInMem_hi_lo_87};
  wire [31:0]      dataInMem_lo_280 = {dataInMem_lo_hi_152, dataInMem_lo_lo_24};
  wire [15:0]      dataInMem_hi_hi_216 = {dataRegroupBySew_7_17, dataRegroupBySew_6_17};
  wire [31:0]      dataInMem_hi_344 = {dataInMem_hi_hi_216, dataInMem_hi_lo_88};
  wire [31:0]      dataInMem_lo_281 = {dataInMem_lo_hi_153, dataInMem_lo_lo_25};
  wire [15:0]      dataInMem_hi_hi_217 = {dataRegroupBySew_7_18, dataRegroupBySew_6_18};
  wire [31:0]      dataInMem_hi_345 = {dataInMem_hi_hi_217, dataInMem_hi_lo_89};
  wire [31:0]      dataInMem_lo_282 = {dataInMem_lo_hi_154, dataInMem_lo_lo_26};
  wire [15:0]      dataInMem_hi_hi_218 = {dataRegroupBySew_7_19, dataRegroupBySew_6_19};
  wire [31:0]      dataInMem_hi_346 = {dataInMem_hi_hi_218, dataInMem_hi_lo_90};
  wire [31:0]      dataInMem_lo_283 = {dataInMem_lo_hi_155, dataInMem_lo_lo_27};
  wire [15:0]      dataInMem_hi_hi_219 = {dataRegroupBySew_7_20, dataRegroupBySew_6_20};
  wire [31:0]      dataInMem_hi_347 = {dataInMem_hi_hi_219, dataInMem_hi_lo_91};
  wire [31:0]      dataInMem_lo_284 = {dataInMem_lo_hi_156, dataInMem_lo_lo_28};
  wire [15:0]      dataInMem_hi_hi_220 = {dataRegroupBySew_7_21, dataRegroupBySew_6_21};
  wire [31:0]      dataInMem_hi_348 = {dataInMem_hi_hi_220, dataInMem_hi_lo_92};
  wire [31:0]      dataInMem_lo_285 = {dataInMem_lo_hi_157, dataInMem_lo_lo_29};
  wire [15:0]      dataInMem_hi_hi_221 = {dataRegroupBySew_7_22, dataRegroupBySew_6_22};
  wire [31:0]      dataInMem_hi_349 = {dataInMem_hi_hi_221, dataInMem_hi_lo_93};
  wire [31:0]      dataInMem_lo_286 = {dataInMem_lo_hi_158, dataInMem_lo_lo_30};
  wire [15:0]      dataInMem_hi_hi_222 = {dataRegroupBySew_7_23, dataRegroupBySew_6_23};
  wire [31:0]      dataInMem_hi_350 = {dataInMem_hi_hi_222, dataInMem_hi_lo_94};
  wire [31:0]      dataInMem_lo_287 = {dataInMem_lo_hi_159, dataInMem_lo_lo_31};
  wire [15:0]      dataInMem_hi_hi_223 = {dataRegroupBySew_7_24, dataRegroupBySew_6_24};
  wire [31:0]      dataInMem_hi_351 = {dataInMem_hi_hi_223, dataInMem_hi_lo_95};
  wire [31:0]      dataInMem_lo_288 = {dataInMem_lo_hi_160, dataInMem_lo_lo_32};
  wire [15:0]      dataInMem_hi_hi_224 = {dataRegroupBySew_7_25, dataRegroupBySew_6_25};
  wire [31:0]      dataInMem_hi_352 = {dataInMem_hi_hi_224, dataInMem_hi_lo_96};
  wire [31:0]      dataInMem_lo_289 = {dataInMem_lo_hi_161, dataInMem_lo_lo_33};
  wire [15:0]      dataInMem_hi_hi_225 = {dataRegroupBySew_7_26, dataRegroupBySew_6_26};
  wire [31:0]      dataInMem_hi_353 = {dataInMem_hi_hi_225, dataInMem_hi_lo_97};
  wire [31:0]      dataInMem_lo_290 = {dataInMem_lo_hi_162, dataInMem_lo_lo_34};
  wire [15:0]      dataInMem_hi_hi_226 = {dataRegroupBySew_7_27, dataRegroupBySew_6_27};
  wire [31:0]      dataInMem_hi_354 = {dataInMem_hi_hi_226, dataInMem_hi_lo_98};
  wire [31:0]      dataInMem_lo_291 = {dataInMem_lo_hi_163, dataInMem_lo_lo_35};
  wire [15:0]      dataInMem_hi_hi_227 = {dataRegroupBySew_7_28, dataRegroupBySew_6_28};
  wire [31:0]      dataInMem_hi_355 = {dataInMem_hi_hi_227, dataInMem_hi_lo_99};
  wire [31:0]      dataInMem_lo_292 = {dataInMem_lo_hi_164, dataInMem_lo_lo_36};
  wire [15:0]      dataInMem_hi_hi_228 = {dataRegroupBySew_7_29, dataRegroupBySew_6_29};
  wire [31:0]      dataInMem_hi_356 = {dataInMem_hi_hi_228, dataInMem_hi_lo_100};
  wire [31:0]      dataInMem_lo_293 = {dataInMem_lo_hi_165, dataInMem_lo_lo_37};
  wire [15:0]      dataInMem_hi_hi_229 = {dataRegroupBySew_7_30, dataRegroupBySew_6_30};
  wire [31:0]      dataInMem_hi_357 = {dataInMem_hi_hi_229, dataInMem_hi_lo_101};
  wire [31:0]      dataInMem_lo_294 = {dataInMem_lo_hi_166, dataInMem_lo_lo_38};
  wire [15:0]      dataInMem_hi_hi_230 = {dataRegroupBySew_7_31, dataRegroupBySew_6_31};
  wire [31:0]      dataInMem_hi_358 = {dataInMem_hi_hi_230, dataInMem_hi_lo_102};
  wire [31:0]      dataInMem_lo_295 = {dataInMem_lo_hi_167, dataInMem_lo_lo_39};
  wire [15:0]      dataInMem_hi_hi_231 = {dataRegroupBySew_7_32, dataRegroupBySew_6_32};
  wire [31:0]      dataInMem_hi_359 = {dataInMem_hi_hi_231, dataInMem_hi_lo_103};
  wire [31:0]      dataInMem_lo_296 = {dataInMem_lo_hi_168, dataInMem_lo_lo_40};
  wire [15:0]      dataInMem_hi_hi_232 = {dataRegroupBySew_7_33, dataRegroupBySew_6_33};
  wire [31:0]      dataInMem_hi_360 = {dataInMem_hi_hi_232, dataInMem_hi_lo_104};
  wire [31:0]      dataInMem_lo_297 = {dataInMem_lo_hi_169, dataInMem_lo_lo_41};
  wire [15:0]      dataInMem_hi_hi_233 = {dataRegroupBySew_7_34, dataRegroupBySew_6_34};
  wire [31:0]      dataInMem_hi_361 = {dataInMem_hi_hi_233, dataInMem_hi_lo_105};
  wire [31:0]      dataInMem_lo_298 = {dataInMem_lo_hi_170, dataInMem_lo_lo_42};
  wire [15:0]      dataInMem_hi_hi_234 = {dataRegroupBySew_7_35, dataRegroupBySew_6_35};
  wire [31:0]      dataInMem_hi_362 = {dataInMem_hi_hi_234, dataInMem_hi_lo_106};
  wire [31:0]      dataInMem_lo_299 = {dataInMem_lo_hi_171, dataInMem_lo_lo_43};
  wire [15:0]      dataInMem_hi_hi_235 = {dataRegroupBySew_7_36, dataRegroupBySew_6_36};
  wire [31:0]      dataInMem_hi_363 = {dataInMem_hi_hi_235, dataInMem_hi_lo_107};
  wire [31:0]      dataInMem_lo_300 = {dataInMem_lo_hi_172, dataInMem_lo_lo_44};
  wire [15:0]      dataInMem_hi_hi_236 = {dataRegroupBySew_7_37, dataRegroupBySew_6_37};
  wire [31:0]      dataInMem_hi_364 = {dataInMem_hi_hi_236, dataInMem_hi_lo_108};
  wire [31:0]      dataInMem_lo_301 = {dataInMem_lo_hi_173, dataInMem_lo_lo_45};
  wire [15:0]      dataInMem_hi_hi_237 = {dataRegroupBySew_7_38, dataRegroupBySew_6_38};
  wire [31:0]      dataInMem_hi_365 = {dataInMem_hi_hi_237, dataInMem_hi_lo_109};
  wire [31:0]      dataInMem_lo_302 = {dataInMem_lo_hi_174, dataInMem_lo_lo_46};
  wire [15:0]      dataInMem_hi_hi_238 = {dataRegroupBySew_7_39, dataRegroupBySew_6_39};
  wire [31:0]      dataInMem_hi_366 = {dataInMem_hi_hi_238, dataInMem_hi_lo_110};
  wire [31:0]      dataInMem_lo_303 = {dataInMem_lo_hi_175, dataInMem_lo_lo_47};
  wire [15:0]      dataInMem_hi_hi_239 = {dataRegroupBySew_7_40, dataRegroupBySew_6_40};
  wire [31:0]      dataInMem_hi_367 = {dataInMem_hi_hi_239, dataInMem_hi_lo_111};
  wire [31:0]      dataInMem_lo_304 = {dataInMem_lo_hi_176, dataInMem_lo_lo_48};
  wire [15:0]      dataInMem_hi_hi_240 = {dataRegroupBySew_7_41, dataRegroupBySew_6_41};
  wire [31:0]      dataInMem_hi_368 = {dataInMem_hi_hi_240, dataInMem_hi_lo_112};
  wire [31:0]      dataInMem_lo_305 = {dataInMem_lo_hi_177, dataInMem_lo_lo_49};
  wire [15:0]      dataInMem_hi_hi_241 = {dataRegroupBySew_7_42, dataRegroupBySew_6_42};
  wire [31:0]      dataInMem_hi_369 = {dataInMem_hi_hi_241, dataInMem_hi_lo_113};
  wire [31:0]      dataInMem_lo_306 = {dataInMem_lo_hi_178, dataInMem_lo_lo_50};
  wire [15:0]      dataInMem_hi_hi_242 = {dataRegroupBySew_7_43, dataRegroupBySew_6_43};
  wire [31:0]      dataInMem_hi_370 = {dataInMem_hi_hi_242, dataInMem_hi_lo_114};
  wire [31:0]      dataInMem_lo_307 = {dataInMem_lo_hi_179, dataInMem_lo_lo_51};
  wire [15:0]      dataInMem_hi_hi_243 = {dataRegroupBySew_7_44, dataRegroupBySew_6_44};
  wire [31:0]      dataInMem_hi_371 = {dataInMem_hi_hi_243, dataInMem_hi_lo_115};
  wire [31:0]      dataInMem_lo_308 = {dataInMem_lo_hi_180, dataInMem_lo_lo_52};
  wire [15:0]      dataInMem_hi_hi_244 = {dataRegroupBySew_7_45, dataRegroupBySew_6_45};
  wire [31:0]      dataInMem_hi_372 = {dataInMem_hi_hi_244, dataInMem_hi_lo_116};
  wire [31:0]      dataInMem_lo_309 = {dataInMem_lo_hi_181, dataInMem_lo_lo_53};
  wire [15:0]      dataInMem_hi_hi_245 = {dataRegroupBySew_7_46, dataRegroupBySew_6_46};
  wire [31:0]      dataInMem_hi_373 = {dataInMem_hi_hi_245, dataInMem_hi_lo_117};
  wire [31:0]      dataInMem_lo_310 = {dataInMem_lo_hi_182, dataInMem_lo_lo_54};
  wire [15:0]      dataInMem_hi_hi_246 = {dataRegroupBySew_7_47, dataRegroupBySew_6_47};
  wire [31:0]      dataInMem_hi_374 = {dataInMem_hi_hi_246, dataInMem_hi_lo_118};
  wire [31:0]      dataInMem_lo_311 = {dataInMem_lo_hi_183, dataInMem_lo_lo_55};
  wire [15:0]      dataInMem_hi_hi_247 = {dataRegroupBySew_7_48, dataRegroupBySew_6_48};
  wire [31:0]      dataInMem_hi_375 = {dataInMem_hi_hi_247, dataInMem_hi_lo_119};
  wire [31:0]      dataInMem_lo_312 = {dataInMem_lo_hi_184, dataInMem_lo_lo_56};
  wire [15:0]      dataInMem_hi_hi_248 = {dataRegroupBySew_7_49, dataRegroupBySew_6_49};
  wire [31:0]      dataInMem_hi_376 = {dataInMem_hi_hi_248, dataInMem_hi_lo_120};
  wire [31:0]      dataInMem_lo_313 = {dataInMem_lo_hi_185, dataInMem_lo_lo_57};
  wire [15:0]      dataInMem_hi_hi_249 = {dataRegroupBySew_7_50, dataRegroupBySew_6_50};
  wire [31:0]      dataInMem_hi_377 = {dataInMem_hi_hi_249, dataInMem_hi_lo_121};
  wire [31:0]      dataInMem_lo_314 = {dataInMem_lo_hi_186, dataInMem_lo_lo_58};
  wire [15:0]      dataInMem_hi_hi_250 = {dataRegroupBySew_7_51, dataRegroupBySew_6_51};
  wire [31:0]      dataInMem_hi_378 = {dataInMem_hi_hi_250, dataInMem_hi_lo_122};
  wire [31:0]      dataInMem_lo_315 = {dataInMem_lo_hi_187, dataInMem_lo_lo_59};
  wire [15:0]      dataInMem_hi_hi_251 = {dataRegroupBySew_7_52, dataRegroupBySew_6_52};
  wire [31:0]      dataInMem_hi_379 = {dataInMem_hi_hi_251, dataInMem_hi_lo_123};
  wire [31:0]      dataInMem_lo_316 = {dataInMem_lo_hi_188, dataInMem_lo_lo_60};
  wire [15:0]      dataInMem_hi_hi_252 = {dataRegroupBySew_7_53, dataRegroupBySew_6_53};
  wire [31:0]      dataInMem_hi_380 = {dataInMem_hi_hi_252, dataInMem_hi_lo_124};
  wire [31:0]      dataInMem_lo_317 = {dataInMem_lo_hi_189, dataInMem_lo_lo_61};
  wire [15:0]      dataInMem_hi_hi_253 = {dataRegroupBySew_7_54, dataRegroupBySew_6_54};
  wire [31:0]      dataInMem_hi_381 = {dataInMem_hi_hi_253, dataInMem_hi_lo_125};
  wire [31:0]      dataInMem_lo_318 = {dataInMem_lo_hi_190, dataInMem_lo_lo_62};
  wire [15:0]      dataInMem_hi_hi_254 = {dataRegroupBySew_7_55, dataRegroupBySew_6_55};
  wire [31:0]      dataInMem_hi_382 = {dataInMem_hi_hi_254, dataInMem_hi_lo_126};
  wire [31:0]      dataInMem_lo_319 = {dataInMem_lo_hi_191, dataInMem_lo_lo_63};
  wire [15:0]      dataInMem_hi_hi_255 = {dataRegroupBySew_7_56, dataRegroupBySew_6_56};
  wire [31:0]      dataInMem_hi_383 = {dataInMem_hi_hi_255, dataInMem_hi_lo_127};
  wire [31:0]      dataInMem_lo_320 = {dataInMem_lo_hi_192, dataInMem_lo_lo_64};
  wire [15:0]      dataInMem_hi_hi_256 = {dataRegroupBySew_7_57, dataRegroupBySew_6_57};
  wire [31:0]      dataInMem_hi_384 = {dataInMem_hi_hi_256, dataInMem_hi_lo_128};
  wire [31:0]      dataInMem_lo_321 = {dataInMem_lo_hi_193, dataInMem_lo_lo_65};
  wire [15:0]      dataInMem_hi_hi_257 = {dataRegroupBySew_7_58, dataRegroupBySew_6_58};
  wire [31:0]      dataInMem_hi_385 = {dataInMem_hi_hi_257, dataInMem_hi_lo_129};
  wire [31:0]      dataInMem_lo_322 = {dataInMem_lo_hi_194, dataInMem_lo_lo_66};
  wire [15:0]      dataInMem_hi_hi_258 = {dataRegroupBySew_7_59, dataRegroupBySew_6_59};
  wire [31:0]      dataInMem_hi_386 = {dataInMem_hi_hi_258, dataInMem_hi_lo_130};
  wire [31:0]      dataInMem_lo_323 = {dataInMem_lo_hi_195, dataInMem_lo_lo_67};
  wire [15:0]      dataInMem_hi_hi_259 = {dataRegroupBySew_7_60, dataRegroupBySew_6_60};
  wire [31:0]      dataInMem_hi_387 = {dataInMem_hi_hi_259, dataInMem_hi_lo_131};
  wire [31:0]      dataInMem_lo_324 = {dataInMem_lo_hi_196, dataInMem_lo_lo_68};
  wire [15:0]      dataInMem_hi_hi_260 = {dataRegroupBySew_7_61, dataRegroupBySew_6_61};
  wire [31:0]      dataInMem_hi_388 = {dataInMem_hi_hi_260, dataInMem_hi_lo_132};
  wire [31:0]      dataInMem_lo_325 = {dataInMem_lo_hi_197, dataInMem_lo_lo_69};
  wire [15:0]      dataInMem_hi_hi_261 = {dataRegroupBySew_7_62, dataRegroupBySew_6_62};
  wire [31:0]      dataInMem_hi_389 = {dataInMem_hi_hi_261, dataInMem_hi_lo_133};
  wire [31:0]      dataInMem_lo_326 = {dataInMem_lo_hi_198, dataInMem_lo_lo_70};
  wire [15:0]      dataInMem_hi_hi_262 = {dataRegroupBySew_7_63, dataRegroupBySew_6_63};
  wire [31:0]      dataInMem_hi_390 = {dataInMem_hi_hi_262, dataInMem_hi_lo_134};
  wire [127:0]     dataInMem_lo_lo_lo_lo_lo_7 = {dataInMem_hi_328, dataInMem_lo_264, dataInMem_hi_327, dataInMem_lo_263};
  wire [127:0]     dataInMem_lo_lo_lo_lo_hi_7 = {dataInMem_hi_330, dataInMem_lo_266, dataInMem_hi_329, dataInMem_lo_265};
  wire [255:0]     dataInMem_lo_lo_lo_lo_7 = {dataInMem_lo_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_lo_lo_hi_lo_7 = {dataInMem_hi_332, dataInMem_lo_268, dataInMem_hi_331, dataInMem_lo_267};
  wire [127:0]     dataInMem_lo_lo_lo_hi_hi_7 = {dataInMem_hi_334, dataInMem_lo_270, dataInMem_hi_333, dataInMem_lo_269};
  wire [255:0]     dataInMem_lo_lo_lo_hi_7 = {dataInMem_lo_lo_lo_hi_hi_7, dataInMem_lo_lo_lo_hi_lo_7};
  wire [511:0]     dataInMem_lo_lo_lo_7 = {dataInMem_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_lo_hi_lo_lo_7 = {dataInMem_hi_336, dataInMem_lo_272, dataInMem_hi_335, dataInMem_lo_271};
  wire [127:0]     dataInMem_lo_lo_hi_lo_hi_7 = {dataInMem_hi_338, dataInMem_lo_274, dataInMem_hi_337, dataInMem_lo_273};
  wire [255:0]     dataInMem_lo_lo_hi_lo_7 = {dataInMem_lo_lo_hi_lo_hi_7, dataInMem_lo_lo_hi_lo_lo_7};
  wire [127:0]     dataInMem_lo_lo_hi_hi_lo_7 = {dataInMem_hi_340, dataInMem_lo_276, dataInMem_hi_339, dataInMem_lo_275};
  wire [127:0]     dataInMem_lo_lo_hi_hi_hi_7 = {dataInMem_hi_342, dataInMem_lo_278, dataInMem_hi_341, dataInMem_lo_277};
  wire [255:0]     dataInMem_lo_lo_hi_hi_7 = {dataInMem_lo_lo_hi_hi_hi_7, dataInMem_lo_lo_hi_hi_lo_7};
  wire [511:0]     dataInMem_lo_lo_hi_7 = {dataInMem_lo_lo_hi_hi_7, dataInMem_lo_lo_hi_lo_7};
  wire [1023:0]    dataInMem_lo_lo_71 = {dataInMem_lo_lo_hi_7, dataInMem_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_lo_lo_lo_7 = {dataInMem_hi_344, dataInMem_lo_280, dataInMem_hi_343, dataInMem_lo_279};
  wire [127:0]     dataInMem_lo_hi_lo_lo_hi_7 = {dataInMem_hi_346, dataInMem_lo_282, dataInMem_hi_345, dataInMem_lo_281};
  wire [255:0]     dataInMem_lo_hi_lo_lo_7 = {dataInMem_lo_hi_lo_lo_hi_7, dataInMem_lo_hi_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_lo_hi_lo_7 = {dataInMem_hi_348, dataInMem_lo_284, dataInMem_hi_347, dataInMem_lo_283};
  wire [127:0]     dataInMem_lo_hi_lo_hi_hi_7 = {dataInMem_hi_350, dataInMem_lo_286, dataInMem_hi_349, dataInMem_lo_285};
  wire [255:0]     dataInMem_lo_hi_lo_hi_7 = {dataInMem_lo_hi_lo_hi_hi_7, dataInMem_lo_hi_lo_hi_lo_7};
  wire [511:0]     dataInMem_lo_hi_lo_7 = {dataInMem_lo_hi_lo_hi_7, dataInMem_lo_hi_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_hi_lo_lo_7 = {dataInMem_hi_352, dataInMem_lo_288, dataInMem_hi_351, dataInMem_lo_287};
  wire [127:0]     dataInMem_lo_hi_hi_lo_hi_7 = {dataInMem_hi_354, dataInMem_lo_290, dataInMem_hi_353, dataInMem_lo_289};
  wire [255:0]     dataInMem_lo_hi_hi_lo_7 = {dataInMem_lo_hi_hi_lo_hi_7, dataInMem_lo_hi_hi_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_hi_hi_lo_7 = {dataInMem_hi_356, dataInMem_lo_292, dataInMem_hi_355, dataInMem_lo_291};
  wire [127:0]     dataInMem_lo_hi_hi_hi_hi_7 = {dataInMem_hi_358, dataInMem_lo_294, dataInMem_hi_357, dataInMem_lo_293};
  wire [255:0]     dataInMem_lo_hi_hi_hi_7 = {dataInMem_lo_hi_hi_hi_hi_7, dataInMem_lo_hi_hi_hi_lo_7};
  wire [511:0]     dataInMem_lo_hi_hi_7 = {dataInMem_lo_hi_hi_hi_7, dataInMem_lo_hi_hi_lo_7};
  wire [1023:0]    dataInMem_lo_hi_199 = {dataInMem_lo_hi_hi_7, dataInMem_lo_hi_lo_7};
  wire [2047:0]    dataInMem_lo_327 = {dataInMem_lo_hi_199, dataInMem_lo_lo_71};
  wire [127:0]     dataInMem_hi_lo_lo_lo_lo_7 = {dataInMem_hi_360, dataInMem_lo_296, dataInMem_hi_359, dataInMem_lo_295};
  wire [127:0]     dataInMem_hi_lo_lo_lo_hi_7 = {dataInMem_hi_362, dataInMem_lo_298, dataInMem_hi_361, dataInMem_lo_297};
  wire [255:0]     dataInMem_hi_lo_lo_lo_7 = {dataInMem_hi_lo_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_lo_7};
  wire [127:0]     dataInMem_hi_lo_lo_hi_lo_7 = {dataInMem_hi_364, dataInMem_lo_300, dataInMem_hi_363, dataInMem_lo_299};
  wire [127:0]     dataInMem_hi_lo_lo_hi_hi_7 = {dataInMem_hi_366, dataInMem_lo_302, dataInMem_hi_365, dataInMem_lo_301};
  wire [255:0]     dataInMem_hi_lo_lo_hi_7 = {dataInMem_hi_lo_lo_hi_hi_7, dataInMem_hi_lo_lo_hi_lo_7};
  wire [511:0]     dataInMem_hi_lo_lo_7 = {dataInMem_hi_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_7};
  wire [127:0]     dataInMem_hi_lo_hi_lo_lo_7 = {dataInMem_hi_368, dataInMem_lo_304, dataInMem_hi_367, dataInMem_lo_303};
  wire [127:0]     dataInMem_hi_lo_hi_lo_hi_7 = {dataInMem_hi_370, dataInMem_lo_306, dataInMem_hi_369, dataInMem_lo_305};
  wire [255:0]     dataInMem_hi_lo_hi_lo_7 = {dataInMem_hi_lo_hi_lo_hi_7, dataInMem_hi_lo_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_lo_hi_hi_lo_7 = {dataInMem_hi_372, dataInMem_lo_308, dataInMem_hi_371, dataInMem_lo_307};
  wire [127:0]     dataInMem_hi_lo_hi_hi_hi_7 = {dataInMem_hi_374, dataInMem_lo_310, dataInMem_hi_373, dataInMem_lo_309};
  wire [255:0]     dataInMem_hi_lo_hi_hi_7 = {dataInMem_hi_lo_hi_hi_hi_7, dataInMem_hi_lo_hi_hi_lo_7};
  wire [511:0]     dataInMem_hi_lo_hi_7 = {dataInMem_hi_lo_hi_hi_7, dataInMem_hi_lo_hi_lo_7};
  wire [1023:0]    dataInMem_hi_lo_135 = {dataInMem_hi_lo_hi_7, dataInMem_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_lo_lo_lo_7 = {dataInMem_hi_376, dataInMem_lo_312, dataInMem_hi_375, dataInMem_lo_311};
  wire [127:0]     dataInMem_hi_hi_lo_lo_hi_7 = {dataInMem_hi_378, dataInMem_lo_314, dataInMem_hi_377, dataInMem_lo_313};
  wire [255:0]     dataInMem_hi_hi_lo_lo_7 = {dataInMem_hi_hi_lo_lo_hi_7, dataInMem_hi_hi_lo_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_lo_hi_lo_7 = {dataInMem_hi_380, dataInMem_lo_316, dataInMem_hi_379, dataInMem_lo_315};
  wire [127:0]     dataInMem_hi_hi_lo_hi_hi_7 = {dataInMem_hi_382, dataInMem_lo_318, dataInMem_hi_381, dataInMem_lo_317};
  wire [255:0]     dataInMem_hi_hi_lo_hi_7 = {dataInMem_hi_hi_lo_hi_hi_7, dataInMem_hi_hi_lo_hi_lo_7};
  wire [511:0]     dataInMem_hi_hi_lo_7 = {dataInMem_hi_hi_lo_hi_7, dataInMem_hi_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_hi_lo_lo_7 = {dataInMem_hi_384, dataInMem_lo_320, dataInMem_hi_383, dataInMem_lo_319};
  wire [127:0]     dataInMem_hi_hi_hi_lo_hi_7 = {dataInMem_hi_386, dataInMem_lo_322, dataInMem_hi_385, dataInMem_lo_321};
  wire [255:0]     dataInMem_hi_hi_hi_lo_7 = {dataInMem_hi_hi_hi_lo_hi_7, dataInMem_hi_hi_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_hi_hi_lo_7 = {dataInMem_hi_388, dataInMem_lo_324, dataInMem_hi_387, dataInMem_lo_323};
  wire [127:0]     dataInMem_hi_hi_hi_hi_hi_7 = {dataInMem_hi_390, dataInMem_lo_326, dataInMem_hi_389, dataInMem_lo_325};
  wire [255:0]     dataInMem_hi_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_hi_lo_7};
  wire [511:0]     dataInMem_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_lo_7};
  wire [1023:0]    dataInMem_hi_hi_263 = {dataInMem_hi_hi_hi_7, dataInMem_hi_hi_lo_7};
  wire [2047:0]    dataInMem_hi_391 = {dataInMem_hi_hi_263, dataInMem_hi_lo_135};
  wire [4095:0]    dataInMem_7 = {dataInMem_hi_391, dataInMem_lo_327};
  wire [511:0]     regroupCacheLine_7_0 = dataInMem_7[511:0];
  wire [511:0]     regroupCacheLine_7_1 = dataInMem_7[1023:512];
  wire [511:0]     regroupCacheLine_7_2 = dataInMem_7[1535:1024];
  wire [511:0]     regroupCacheLine_7_3 = dataInMem_7[2047:1536];
  wire [511:0]     regroupCacheLine_7_4 = dataInMem_7[2559:2048];
  wire [511:0]     regroupCacheLine_7_5 = dataInMem_7[3071:2560];
  wire [511:0]     regroupCacheLine_7_6 = dataInMem_7[3583:3072];
  wire [511:0]     regroupCacheLine_7_7 = dataInMem_7[4095:3584];
  wire [511:0]     res_56 = regroupCacheLine_7_0;
  wire [511:0]     res_57 = regroupCacheLine_7_1;
  wire [511:0]     res_58 = regroupCacheLine_7_2;
  wire [511:0]     res_59 = regroupCacheLine_7_3;
  wire [511:0]     res_60 = regroupCacheLine_7_4;
  wire [511:0]     res_61 = regroupCacheLine_7_5;
  wire [511:0]     res_62 = regroupCacheLine_7_6;
  wire [511:0]     res_63 = regroupCacheLine_7_7;
  wire [1023:0]    lo_lo_7 = {res_57, res_56};
  wire [1023:0]    lo_hi_7 = {res_59, res_58};
  wire [2047:0]    lo_7 = {lo_hi_7, lo_lo_7};
  wire [1023:0]    hi_lo_7 = {res_61, res_60};
  wire [1023:0]    hi_hi_7 = {res_63, res_62};
  wire [2047:0]    hi_7 = {hi_hi_7, hi_lo_7};
  wire [4095:0]    regroupLoadData_0_7 = {hi_7, lo_7};
  wire [15:0]      dataRegroupBySew_0_1_0 = bufferStageEnqueueData_0[15:0];
  wire [15:0]      dataRegroupBySew_0_1_1 = bufferStageEnqueueData_0[31:16];
  wire [15:0]      dataRegroupBySew_0_1_2 = bufferStageEnqueueData_0[47:32];
  wire [15:0]      dataRegroupBySew_0_1_3 = bufferStageEnqueueData_0[63:48];
  wire [15:0]      dataRegroupBySew_0_1_4 = bufferStageEnqueueData_0[79:64];
  wire [15:0]      dataRegroupBySew_0_1_5 = bufferStageEnqueueData_0[95:80];
  wire [15:0]      dataRegroupBySew_0_1_6 = bufferStageEnqueueData_0[111:96];
  wire [15:0]      dataRegroupBySew_0_1_7 = bufferStageEnqueueData_0[127:112];
  wire [15:0]      dataRegroupBySew_0_1_8 = bufferStageEnqueueData_0[143:128];
  wire [15:0]      dataRegroupBySew_0_1_9 = bufferStageEnqueueData_0[159:144];
  wire [15:0]      dataRegroupBySew_0_1_10 = bufferStageEnqueueData_0[175:160];
  wire [15:0]      dataRegroupBySew_0_1_11 = bufferStageEnqueueData_0[191:176];
  wire [15:0]      dataRegroupBySew_0_1_12 = bufferStageEnqueueData_0[207:192];
  wire [15:0]      dataRegroupBySew_0_1_13 = bufferStageEnqueueData_0[223:208];
  wire [15:0]      dataRegroupBySew_0_1_14 = bufferStageEnqueueData_0[239:224];
  wire [15:0]      dataRegroupBySew_0_1_15 = bufferStageEnqueueData_0[255:240];
  wire [15:0]      dataRegroupBySew_0_1_16 = bufferStageEnqueueData_0[271:256];
  wire [15:0]      dataRegroupBySew_0_1_17 = bufferStageEnqueueData_0[287:272];
  wire [15:0]      dataRegroupBySew_0_1_18 = bufferStageEnqueueData_0[303:288];
  wire [15:0]      dataRegroupBySew_0_1_19 = bufferStageEnqueueData_0[319:304];
  wire [15:0]      dataRegroupBySew_0_1_20 = bufferStageEnqueueData_0[335:320];
  wire [15:0]      dataRegroupBySew_0_1_21 = bufferStageEnqueueData_0[351:336];
  wire [15:0]      dataRegroupBySew_0_1_22 = bufferStageEnqueueData_0[367:352];
  wire [15:0]      dataRegroupBySew_0_1_23 = bufferStageEnqueueData_0[383:368];
  wire [15:0]      dataRegroupBySew_0_1_24 = bufferStageEnqueueData_0[399:384];
  wire [15:0]      dataRegroupBySew_0_1_25 = bufferStageEnqueueData_0[415:400];
  wire [15:0]      dataRegroupBySew_0_1_26 = bufferStageEnqueueData_0[431:416];
  wire [15:0]      dataRegroupBySew_0_1_27 = bufferStageEnqueueData_0[447:432];
  wire [15:0]      dataRegroupBySew_0_1_28 = bufferStageEnqueueData_0[463:448];
  wire [15:0]      dataRegroupBySew_0_1_29 = bufferStageEnqueueData_0[479:464];
  wire [15:0]      dataRegroupBySew_0_1_30 = bufferStageEnqueueData_0[495:480];
  wire [15:0]      dataRegroupBySew_0_1_31 = bufferStageEnqueueData_0[511:496];
  wire [15:0]      dataRegroupBySew_1_1_0 = bufferStageEnqueueData_1[15:0];
  wire [15:0]      dataRegroupBySew_1_1_1 = bufferStageEnqueueData_1[31:16];
  wire [15:0]      dataRegroupBySew_1_1_2 = bufferStageEnqueueData_1[47:32];
  wire [15:0]      dataRegroupBySew_1_1_3 = bufferStageEnqueueData_1[63:48];
  wire [15:0]      dataRegroupBySew_1_1_4 = bufferStageEnqueueData_1[79:64];
  wire [15:0]      dataRegroupBySew_1_1_5 = bufferStageEnqueueData_1[95:80];
  wire [15:0]      dataRegroupBySew_1_1_6 = bufferStageEnqueueData_1[111:96];
  wire [15:0]      dataRegroupBySew_1_1_7 = bufferStageEnqueueData_1[127:112];
  wire [15:0]      dataRegroupBySew_1_1_8 = bufferStageEnqueueData_1[143:128];
  wire [15:0]      dataRegroupBySew_1_1_9 = bufferStageEnqueueData_1[159:144];
  wire [15:0]      dataRegroupBySew_1_1_10 = bufferStageEnqueueData_1[175:160];
  wire [15:0]      dataRegroupBySew_1_1_11 = bufferStageEnqueueData_1[191:176];
  wire [15:0]      dataRegroupBySew_1_1_12 = bufferStageEnqueueData_1[207:192];
  wire [15:0]      dataRegroupBySew_1_1_13 = bufferStageEnqueueData_1[223:208];
  wire [15:0]      dataRegroupBySew_1_1_14 = bufferStageEnqueueData_1[239:224];
  wire [15:0]      dataRegroupBySew_1_1_15 = bufferStageEnqueueData_1[255:240];
  wire [15:0]      dataRegroupBySew_1_1_16 = bufferStageEnqueueData_1[271:256];
  wire [15:0]      dataRegroupBySew_1_1_17 = bufferStageEnqueueData_1[287:272];
  wire [15:0]      dataRegroupBySew_1_1_18 = bufferStageEnqueueData_1[303:288];
  wire [15:0]      dataRegroupBySew_1_1_19 = bufferStageEnqueueData_1[319:304];
  wire [15:0]      dataRegroupBySew_1_1_20 = bufferStageEnqueueData_1[335:320];
  wire [15:0]      dataRegroupBySew_1_1_21 = bufferStageEnqueueData_1[351:336];
  wire [15:0]      dataRegroupBySew_1_1_22 = bufferStageEnqueueData_1[367:352];
  wire [15:0]      dataRegroupBySew_1_1_23 = bufferStageEnqueueData_1[383:368];
  wire [15:0]      dataRegroupBySew_1_1_24 = bufferStageEnqueueData_1[399:384];
  wire [15:0]      dataRegroupBySew_1_1_25 = bufferStageEnqueueData_1[415:400];
  wire [15:0]      dataRegroupBySew_1_1_26 = bufferStageEnqueueData_1[431:416];
  wire [15:0]      dataRegroupBySew_1_1_27 = bufferStageEnqueueData_1[447:432];
  wire [15:0]      dataRegroupBySew_1_1_28 = bufferStageEnqueueData_1[463:448];
  wire [15:0]      dataRegroupBySew_1_1_29 = bufferStageEnqueueData_1[479:464];
  wire [15:0]      dataRegroupBySew_1_1_30 = bufferStageEnqueueData_1[495:480];
  wire [15:0]      dataRegroupBySew_1_1_31 = bufferStageEnqueueData_1[511:496];
  wire [15:0]      dataRegroupBySew_2_1_0 = bufferStageEnqueueData_2[15:0];
  wire [15:0]      dataRegroupBySew_2_1_1 = bufferStageEnqueueData_2[31:16];
  wire [15:0]      dataRegroupBySew_2_1_2 = bufferStageEnqueueData_2[47:32];
  wire [15:0]      dataRegroupBySew_2_1_3 = bufferStageEnqueueData_2[63:48];
  wire [15:0]      dataRegroupBySew_2_1_4 = bufferStageEnqueueData_2[79:64];
  wire [15:0]      dataRegroupBySew_2_1_5 = bufferStageEnqueueData_2[95:80];
  wire [15:0]      dataRegroupBySew_2_1_6 = bufferStageEnqueueData_2[111:96];
  wire [15:0]      dataRegroupBySew_2_1_7 = bufferStageEnqueueData_2[127:112];
  wire [15:0]      dataRegroupBySew_2_1_8 = bufferStageEnqueueData_2[143:128];
  wire [15:0]      dataRegroupBySew_2_1_9 = bufferStageEnqueueData_2[159:144];
  wire [15:0]      dataRegroupBySew_2_1_10 = bufferStageEnqueueData_2[175:160];
  wire [15:0]      dataRegroupBySew_2_1_11 = bufferStageEnqueueData_2[191:176];
  wire [15:0]      dataRegroupBySew_2_1_12 = bufferStageEnqueueData_2[207:192];
  wire [15:0]      dataRegroupBySew_2_1_13 = bufferStageEnqueueData_2[223:208];
  wire [15:0]      dataRegroupBySew_2_1_14 = bufferStageEnqueueData_2[239:224];
  wire [15:0]      dataRegroupBySew_2_1_15 = bufferStageEnqueueData_2[255:240];
  wire [15:0]      dataRegroupBySew_2_1_16 = bufferStageEnqueueData_2[271:256];
  wire [15:0]      dataRegroupBySew_2_1_17 = bufferStageEnqueueData_2[287:272];
  wire [15:0]      dataRegroupBySew_2_1_18 = bufferStageEnqueueData_2[303:288];
  wire [15:0]      dataRegroupBySew_2_1_19 = bufferStageEnqueueData_2[319:304];
  wire [15:0]      dataRegroupBySew_2_1_20 = bufferStageEnqueueData_2[335:320];
  wire [15:0]      dataRegroupBySew_2_1_21 = bufferStageEnqueueData_2[351:336];
  wire [15:0]      dataRegroupBySew_2_1_22 = bufferStageEnqueueData_2[367:352];
  wire [15:0]      dataRegroupBySew_2_1_23 = bufferStageEnqueueData_2[383:368];
  wire [15:0]      dataRegroupBySew_2_1_24 = bufferStageEnqueueData_2[399:384];
  wire [15:0]      dataRegroupBySew_2_1_25 = bufferStageEnqueueData_2[415:400];
  wire [15:0]      dataRegroupBySew_2_1_26 = bufferStageEnqueueData_2[431:416];
  wire [15:0]      dataRegroupBySew_2_1_27 = bufferStageEnqueueData_2[447:432];
  wire [15:0]      dataRegroupBySew_2_1_28 = bufferStageEnqueueData_2[463:448];
  wire [15:0]      dataRegroupBySew_2_1_29 = bufferStageEnqueueData_2[479:464];
  wire [15:0]      dataRegroupBySew_2_1_30 = bufferStageEnqueueData_2[495:480];
  wire [15:0]      dataRegroupBySew_2_1_31 = bufferStageEnqueueData_2[511:496];
  wire [15:0]      dataRegroupBySew_3_1_0 = bufferStageEnqueueData_3[15:0];
  wire [15:0]      dataRegroupBySew_3_1_1 = bufferStageEnqueueData_3[31:16];
  wire [15:0]      dataRegroupBySew_3_1_2 = bufferStageEnqueueData_3[47:32];
  wire [15:0]      dataRegroupBySew_3_1_3 = bufferStageEnqueueData_3[63:48];
  wire [15:0]      dataRegroupBySew_3_1_4 = bufferStageEnqueueData_3[79:64];
  wire [15:0]      dataRegroupBySew_3_1_5 = bufferStageEnqueueData_3[95:80];
  wire [15:0]      dataRegroupBySew_3_1_6 = bufferStageEnqueueData_3[111:96];
  wire [15:0]      dataRegroupBySew_3_1_7 = bufferStageEnqueueData_3[127:112];
  wire [15:0]      dataRegroupBySew_3_1_8 = bufferStageEnqueueData_3[143:128];
  wire [15:0]      dataRegroupBySew_3_1_9 = bufferStageEnqueueData_3[159:144];
  wire [15:0]      dataRegroupBySew_3_1_10 = bufferStageEnqueueData_3[175:160];
  wire [15:0]      dataRegroupBySew_3_1_11 = bufferStageEnqueueData_3[191:176];
  wire [15:0]      dataRegroupBySew_3_1_12 = bufferStageEnqueueData_3[207:192];
  wire [15:0]      dataRegroupBySew_3_1_13 = bufferStageEnqueueData_3[223:208];
  wire [15:0]      dataRegroupBySew_3_1_14 = bufferStageEnqueueData_3[239:224];
  wire [15:0]      dataRegroupBySew_3_1_15 = bufferStageEnqueueData_3[255:240];
  wire [15:0]      dataRegroupBySew_3_1_16 = bufferStageEnqueueData_3[271:256];
  wire [15:0]      dataRegroupBySew_3_1_17 = bufferStageEnqueueData_3[287:272];
  wire [15:0]      dataRegroupBySew_3_1_18 = bufferStageEnqueueData_3[303:288];
  wire [15:0]      dataRegroupBySew_3_1_19 = bufferStageEnqueueData_3[319:304];
  wire [15:0]      dataRegroupBySew_3_1_20 = bufferStageEnqueueData_3[335:320];
  wire [15:0]      dataRegroupBySew_3_1_21 = bufferStageEnqueueData_3[351:336];
  wire [15:0]      dataRegroupBySew_3_1_22 = bufferStageEnqueueData_3[367:352];
  wire [15:0]      dataRegroupBySew_3_1_23 = bufferStageEnqueueData_3[383:368];
  wire [15:0]      dataRegroupBySew_3_1_24 = bufferStageEnqueueData_3[399:384];
  wire [15:0]      dataRegroupBySew_3_1_25 = bufferStageEnqueueData_3[415:400];
  wire [15:0]      dataRegroupBySew_3_1_26 = bufferStageEnqueueData_3[431:416];
  wire [15:0]      dataRegroupBySew_3_1_27 = bufferStageEnqueueData_3[447:432];
  wire [15:0]      dataRegroupBySew_3_1_28 = bufferStageEnqueueData_3[463:448];
  wire [15:0]      dataRegroupBySew_3_1_29 = bufferStageEnqueueData_3[479:464];
  wire [15:0]      dataRegroupBySew_3_1_30 = bufferStageEnqueueData_3[495:480];
  wire [15:0]      dataRegroupBySew_3_1_31 = bufferStageEnqueueData_3[511:496];
  wire [15:0]      dataRegroupBySew_4_1_0 = bufferStageEnqueueData_4[15:0];
  wire [15:0]      dataRegroupBySew_4_1_1 = bufferStageEnqueueData_4[31:16];
  wire [15:0]      dataRegroupBySew_4_1_2 = bufferStageEnqueueData_4[47:32];
  wire [15:0]      dataRegroupBySew_4_1_3 = bufferStageEnqueueData_4[63:48];
  wire [15:0]      dataRegroupBySew_4_1_4 = bufferStageEnqueueData_4[79:64];
  wire [15:0]      dataRegroupBySew_4_1_5 = bufferStageEnqueueData_4[95:80];
  wire [15:0]      dataRegroupBySew_4_1_6 = bufferStageEnqueueData_4[111:96];
  wire [15:0]      dataRegroupBySew_4_1_7 = bufferStageEnqueueData_4[127:112];
  wire [15:0]      dataRegroupBySew_4_1_8 = bufferStageEnqueueData_4[143:128];
  wire [15:0]      dataRegroupBySew_4_1_9 = bufferStageEnqueueData_4[159:144];
  wire [15:0]      dataRegroupBySew_4_1_10 = bufferStageEnqueueData_4[175:160];
  wire [15:0]      dataRegroupBySew_4_1_11 = bufferStageEnqueueData_4[191:176];
  wire [15:0]      dataRegroupBySew_4_1_12 = bufferStageEnqueueData_4[207:192];
  wire [15:0]      dataRegroupBySew_4_1_13 = bufferStageEnqueueData_4[223:208];
  wire [15:0]      dataRegroupBySew_4_1_14 = bufferStageEnqueueData_4[239:224];
  wire [15:0]      dataRegroupBySew_4_1_15 = bufferStageEnqueueData_4[255:240];
  wire [15:0]      dataRegroupBySew_4_1_16 = bufferStageEnqueueData_4[271:256];
  wire [15:0]      dataRegroupBySew_4_1_17 = bufferStageEnqueueData_4[287:272];
  wire [15:0]      dataRegroupBySew_4_1_18 = bufferStageEnqueueData_4[303:288];
  wire [15:0]      dataRegroupBySew_4_1_19 = bufferStageEnqueueData_4[319:304];
  wire [15:0]      dataRegroupBySew_4_1_20 = bufferStageEnqueueData_4[335:320];
  wire [15:0]      dataRegroupBySew_4_1_21 = bufferStageEnqueueData_4[351:336];
  wire [15:0]      dataRegroupBySew_4_1_22 = bufferStageEnqueueData_4[367:352];
  wire [15:0]      dataRegroupBySew_4_1_23 = bufferStageEnqueueData_4[383:368];
  wire [15:0]      dataRegroupBySew_4_1_24 = bufferStageEnqueueData_4[399:384];
  wire [15:0]      dataRegroupBySew_4_1_25 = bufferStageEnqueueData_4[415:400];
  wire [15:0]      dataRegroupBySew_4_1_26 = bufferStageEnqueueData_4[431:416];
  wire [15:0]      dataRegroupBySew_4_1_27 = bufferStageEnqueueData_4[447:432];
  wire [15:0]      dataRegroupBySew_4_1_28 = bufferStageEnqueueData_4[463:448];
  wire [15:0]      dataRegroupBySew_4_1_29 = bufferStageEnqueueData_4[479:464];
  wire [15:0]      dataRegroupBySew_4_1_30 = bufferStageEnqueueData_4[495:480];
  wire [15:0]      dataRegroupBySew_4_1_31 = bufferStageEnqueueData_4[511:496];
  wire [15:0]      dataRegroupBySew_5_1_0 = bufferStageEnqueueData_5[15:0];
  wire [15:0]      dataRegroupBySew_5_1_1 = bufferStageEnqueueData_5[31:16];
  wire [15:0]      dataRegroupBySew_5_1_2 = bufferStageEnqueueData_5[47:32];
  wire [15:0]      dataRegroupBySew_5_1_3 = bufferStageEnqueueData_5[63:48];
  wire [15:0]      dataRegroupBySew_5_1_4 = bufferStageEnqueueData_5[79:64];
  wire [15:0]      dataRegroupBySew_5_1_5 = bufferStageEnqueueData_5[95:80];
  wire [15:0]      dataRegroupBySew_5_1_6 = bufferStageEnqueueData_5[111:96];
  wire [15:0]      dataRegroupBySew_5_1_7 = bufferStageEnqueueData_5[127:112];
  wire [15:0]      dataRegroupBySew_5_1_8 = bufferStageEnqueueData_5[143:128];
  wire [15:0]      dataRegroupBySew_5_1_9 = bufferStageEnqueueData_5[159:144];
  wire [15:0]      dataRegroupBySew_5_1_10 = bufferStageEnqueueData_5[175:160];
  wire [15:0]      dataRegroupBySew_5_1_11 = bufferStageEnqueueData_5[191:176];
  wire [15:0]      dataRegroupBySew_5_1_12 = bufferStageEnqueueData_5[207:192];
  wire [15:0]      dataRegroupBySew_5_1_13 = bufferStageEnqueueData_5[223:208];
  wire [15:0]      dataRegroupBySew_5_1_14 = bufferStageEnqueueData_5[239:224];
  wire [15:0]      dataRegroupBySew_5_1_15 = bufferStageEnqueueData_5[255:240];
  wire [15:0]      dataRegroupBySew_5_1_16 = bufferStageEnqueueData_5[271:256];
  wire [15:0]      dataRegroupBySew_5_1_17 = bufferStageEnqueueData_5[287:272];
  wire [15:0]      dataRegroupBySew_5_1_18 = bufferStageEnqueueData_5[303:288];
  wire [15:0]      dataRegroupBySew_5_1_19 = bufferStageEnqueueData_5[319:304];
  wire [15:0]      dataRegroupBySew_5_1_20 = bufferStageEnqueueData_5[335:320];
  wire [15:0]      dataRegroupBySew_5_1_21 = bufferStageEnqueueData_5[351:336];
  wire [15:0]      dataRegroupBySew_5_1_22 = bufferStageEnqueueData_5[367:352];
  wire [15:0]      dataRegroupBySew_5_1_23 = bufferStageEnqueueData_5[383:368];
  wire [15:0]      dataRegroupBySew_5_1_24 = bufferStageEnqueueData_5[399:384];
  wire [15:0]      dataRegroupBySew_5_1_25 = bufferStageEnqueueData_5[415:400];
  wire [15:0]      dataRegroupBySew_5_1_26 = bufferStageEnqueueData_5[431:416];
  wire [15:0]      dataRegroupBySew_5_1_27 = bufferStageEnqueueData_5[447:432];
  wire [15:0]      dataRegroupBySew_5_1_28 = bufferStageEnqueueData_5[463:448];
  wire [15:0]      dataRegroupBySew_5_1_29 = bufferStageEnqueueData_5[479:464];
  wire [15:0]      dataRegroupBySew_5_1_30 = bufferStageEnqueueData_5[495:480];
  wire [15:0]      dataRegroupBySew_5_1_31 = bufferStageEnqueueData_5[511:496];
  wire [15:0]      dataRegroupBySew_6_1_0 = bufferStageEnqueueData_6[15:0];
  wire [15:0]      dataRegroupBySew_6_1_1 = bufferStageEnqueueData_6[31:16];
  wire [15:0]      dataRegroupBySew_6_1_2 = bufferStageEnqueueData_6[47:32];
  wire [15:0]      dataRegroupBySew_6_1_3 = bufferStageEnqueueData_6[63:48];
  wire [15:0]      dataRegroupBySew_6_1_4 = bufferStageEnqueueData_6[79:64];
  wire [15:0]      dataRegroupBySew_6_1_5 = bufferStageEnqueueData_6[95:80];
  wire [15:0]      dataRegroupBySew_6_1_6 = bufferStageEnqueueData_6[111:96];
  wire [15:0]      dataRegroupBySew_6_1_7 = bufferStageEnqueueData_6[127:112];
  wire [15:0]      dataRegroupBySew_6_1_8 = bufferStageEnqueueData_6[143:128];
  wire [15:0]      dataRegroupBySew_6_1_9 = bufferStageEnqueueData_6[159:144];
  wire [15:0]      dataRegroupBySew_6_1_10 = bufferStageEnqueueData_6[175:160];
  wire [15:0]      dataRegroupBySew_6_1_11 = bufferStageEnqueueData_6[191:176];
  wire [15:0]      dataRegroupBySew_6_1_12 = bufferStageEnqueueData_6[207:192];
  wire [15:0]      dataRegroupBySew_6_1_13 = bufferStageEnqueueData_6[223:208];
  wire [15:0]      dataRegroupBySew_6_1_14 = bufferStageEnqueueData_6[239:224];
  wire [15:0]      dataRegroupBySew_6_1_15 = bufferStageEnqueueData_6[255:240];
  wire [15:0]      dataRegroupBySew_6_1_16 = bufferStageEnqueueData_6[271:256];
  wire [15:0]      dataRegroupBySew_6_1_17 = bufferStageEnqueueData_6[287:272];
  wire [15:0]      dataRegroupBySew_6_1_18 = bufferStageEnqueueData_6[303:288];
  wire [15:0]      dataRegroupBySew_6_1_19 = bufferStageEnqueueData_6[319:304];
  wire [15:0]      dataRegroupBySew_6_1_20 = bufferStageEnqueueData_6[335:320];
  wire [15:0]      dataRegroupBySew_6_1_21 = bufferStageEnqueueData_6[351:336];
  wire [15:0]      dataRegroupBySew_6_1_22 = bufferStageEnqueueData_6[367:352];
  wire [15:0]      dataRegroupBySew_6_1_23 = bufferStageEnqueueData_6[383:368];
  wire [15:0]      dataRegroupBySew_6_1_24 = bufferStageEnqueueData_6[399:384];
  wire [15:0]      dataRegroupBySew_6_1_25 = bufferStageEnqueueData_6[415:400];
  wire [15:0]      dataRegroupBySew_6_1_26 = bufferStageEnqueueData_6[431:416];
  wire [15:0]      dataRegroupBySew_6_1_27 = bufferStageEnqueueData_6[447:432];
  wire [15:0]      dataRegroupBySew_6_1_28 = bufferStageEnqueueData_6[463:448];
  wire [15:0]      dataRegroupBySew_6_1_29 = bufferStageEnqueueData_6[479:464];
  wire [15:0]      dataRegroupBySew_6_1_30 = bufferStageEnqueueData_6[495:480];
  wire [15:0]      dataRegroupBySew_6_1_31 = bufferStageEnqueueData_6[511:496];
  wire [15:0]      dataRegroupBySew_7_1_0 = bufferStageEnqueueData_7[15:0];
  wire [15:0]      dataRegroupBySew_7_1_1 = bufferStageEnqueueData_7[31:16];
  wire [15:0]      dataRegroupBySew_7_1_2 = bufferStageEnqueueData_7[47:32];
  wire [15:0]      dataRegroupBySew_7_1_3 = bufferStageEnqueueData_7[63:48];
  wire [15:0]      dataRegroupBySew_7_1_4 = bufferStageEnqueueData_7[79:64];
  wire [15:0]      dataRegroupBySew_7_1_5 = bufferStageEnqueueData_7[95:80];
  wire [15:0]      dataRegroupBySew_7_1_6 = bufferStageEnqueueData_7[111:96];
  wire [15:0]      dataRegroupBySew_7_1_7 = bufferStageEnqueueData_7[127:112];
  wire [15:0]      dataRegroupBySew_7_1_8 = bufferStageEnqueueData_7[143:128];
  wire [15:0]      dataRegroupBySew_7_1_9 = bufferStageEnqueueData_7[159:144];
  wire [15:0]      dataRegroupBySew_7_1_10 = bufferStageEnqueueData_7[175:160];
  wire [15:0]      dataRegroupBySew_7_1_11 = bufferStageEnqueueData_7[191:176];
  wire [15:0]      dataRegroupBySew_7_1_12 = bufferStageEnqueueData_7[207:192];
  wire [15:0]      dataRegroupBySew_7_1_13 = bufferStageEnqueueData_7[223:208];
  wire [15:0]      dataRegroupBySew_7_1_14 = bufferStageEnqueueData_7[239:224];
  wire [15:0]      dataRegroupBySew_7_1_15 = bufferStageEnqueueData_7[255:240];
  wire [15:0]      dataRegroupBySew_7_1_16 = bufferStageEnqueueData_7[271:256];
  wire [15:0]      dataRegroupBySew_7_1_17 = bufferStageEnqueueData_7[287:272];
  wire [15:0]      dataRegroupBySew_7_1_18 = bufferStageEnqueueData_7[303:288];
  wire [15:0]      dataRegroupBySew_7_1_19 = bufferStageEnqueueData_7[319:304];
  wire [15:0]      dataRegroupBySew_7_1_20 = bufferStageEnqueueData_7[335:320];
  wire [15:0]      dataRegroupBySew_7_1_21 = bufferStageEnqueueData_7[351:336];
  wire [15:0]      dataRegroupBySew_7_1_22 = bufferStageEnqueueData_7[367:352];
  wire [15:0]      dataRegroupBySew_7_1_23 = bufferStageEnqueueData_7[383:368];
  wire [15:0]      dataRegroupBySew_7_1_24 = bufferStageEnqueueData_7[399:384];
  wire [15:0]      dataRegroupBySew_7_1_25 = bufferStageEnqueueData_7[415:400];
  wire [15:0]      dataRegroupBySew_7_1_26 = bufferStageEnqueueData_7[431:416];
  wire [15:0]      dataRegroupBySew_7_1_27 = bufferStageEnqueueData_7[447:432];
  wire [15:0]      dataRegroupBySew_7_1_28 = bufferStageEnqueueData_7[463:448];
  wire [15:0]      dataRegroupBySew_7_1_29 = bufferStageEnqueueData_7[479:464];
  wire [15:0]      dataRegroupBySew_7_1_30 = bufferStageEnqueueData_7[495:480];
  wire [15:0]      dataRegroupBySew_7_1_31 = bufferStageEnqueueData_7[511:496];
  wire [31:0]      dataInMem_lo_lo_lo_lo_8 = {dataRegroupBySew_0_1_1, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_lo_lo_hi_8 = {dataRegroupBySew_0_1_3, dataRegroupBySew_0_1_2};
  wire [63:0]      dataInMem_lo_lo_lo_8 = {dataInMem_lo_lo_lo_hi_8, dataInMem_lo_lo_lo_lo_8};
  wire [31:0]      dataInMem_lo_lo_hi_lo_8 = {dataRegroupBySew_0_1_5, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_lo_lo_hi_hi_8 = {dataRegroupBySew_0_1_7, dataRegroupBySew_0_1_6};
  wire [63:0]      dataInMem_lo_lo_hi_8 = {dataInMem_lo_lo_hi_hi_8, dataInMem_lo_lo_hi_lo_8};
  wire [127:0]     dataInMem_lo_lo_72 = {dataInMem_lo_lo_hi_8, dataInMem_lo_lo_lo_8};
  wire [31:0]      dataInMem_lo_hi_lo_lo_8 = {dataRegroupBySew_0_1_9, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_lo_hi_lo_hi_8 = {dataRegroupBySew_0_1_11, dataRegroupBySew_0_1_10};
  wire [63:0]      dataInMem_lo_hi_lo_8 = {dataInMem_lo_hi_lo_hi_8, dataInMem_lo_hi_lo_lo_8};
  wire [31:0]      dataInMem_lo_hi_hi_lo_8 = {dataRegroupBySew_0_1_13, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_lo_hi_hi_hi_8 = {dataRegroupBySew_0_1_15, dataRegroupBySew_0_1_14};
  wire [63:0]      dataInMem_lo_hi_hi_8 = {dataInMem_lo_hi_hi_hi_8, dataInMem_lo_hi_hi_lo_8};
  wire [127:0]     dataInMem_lo_hi_200 = {dataInMem_lo_hi_hi_8, dataInMem_lo_hi_lo_8};
  wire [255:0]     dataInMem_lo_328 = {dataInMem_lo_hi_200, dataInMem_lo_lo_72};
  wire [31:0]      dataInMem_hi_lo_lo_lo_8 = {dataRegroupBySew_0_1_17, dataRegroupBySew_0_1_16};
  wire [31:0]      dataInMem_hi_lo_lo_hi_8 = {dataRegroupBySew_0_1_19, dataRegroupBySew_0_1_18};
  wire [63:0]      dataInMem_hi_lo_lo_8 = {dataInMem_hi_lo_lo_hi_8, dataInMem_hi_lo_lo_lo_8};
  wire [31:0]      dataInMem_hi_lo_hi_lo_8 = {dataRegroupBySew_0_1_21, dataRegroupBySew_0_1_20};
  wire [31:0]      dataInMem_hi_lo_hi_hi_8 = {dataRegroupBySew_0_1_23, dataRegroupBySew_0_1_22};
  wire [63:0]      dataInMem_hi_lo_hi_8 = {dataInMem_hi_lo_hi_hi_8, dataInMem_hi_lo_hi_lo_8};
  wire [127:0]     dataInMem_hi_lo_136 = {dataInMem_hi_lo_hi_8, dataInMem_hi_lo_lo_8};
  wire [31:0]      dataInMem_hi_hi_lo_lo_8 = {dataRegroupBySew_0_1_25, dataRegroupBySew_0_1_24};
  wire [31:0]      dataInMem_hi_hi_lo_hi_8 = {dataRegroupBySew_0_1_27, dataRegroupBySew_0_1_26};
  wire [63:0]      dataInMem_hi_hi_lo_8 = {dataInMem_hi_hi_lo_hi_8, dataInMem_hi_hi_lo_lo_8};
  wire [31:0]      dataInMem_hi_hi_hi_lo_8 = {dataRegroupBySew_0_1_29, dataRegroupBySew_0_1_28};
  wire [31:0]      dataInMem_hi_hi_hi_hi_8 = {dataRegroupBySew_0_1_31, dataRegroupBySew_0_1_30};
  wire [63:0]      dataInMem_hi_hi_hi_8 = {dataInMem_hi_hi_hi_hi_8, dataInMem_hi_hi_hi_lo_8};
  wire [127:0]     dataInMem_hi_hi_264 = {dataInMem_hi_hi_hi_8, dataInMem_hi_hi_lo_8};
  wire [255:0]     dataInMem_hi_392 = {dataInMem_hi_hi_264, dataInMem_hi_lo_136};
  wire [511:0]     dataInMem_8 = {dataInMem_hi_392, dataInMem_lo_328};
  wire [511:0]     regroupCacheLine_8_0 = dataInMem_8;
  wire [511:0]     res_64 = regroupCacheLine_8_0;
  wire [1023:0]    lo_lo_8 = {512'h0, res_64};
  wire [2047:0]    lo_8 = {1024'h0, lo_lo_8};
  wire [4095:0]    regroupLoadData_1_0 = {2048'h0, lo_8};
  wire [63:0]      dataInMem_lo_lo_lo_lo_9 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1, dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [63:0]      dataInMem_lo_lo_lo_hi_9 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3, dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [127:0]     dataInMem_lo_lo_lo_9 = {dataInMem_lo_lo_lo_hi_9, dataInMem_lo_lo_lo_lo_9};
  wire [63:0]      dataInMem_lo_lo_hi_lo_9 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5, dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [63:0]      dataInMem_lo_lo_hi_hi_9 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7, dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [127:0]     dataInMem_lo_lo_hi_9 = {dataInMem_lo_lo_hi_hi_9, dataInMem_lo_lo_hi_lo_9};
  wire [255:0]     dataInMem_lo_lo_73 = {dataInMem_lo_lo_hi_9, dataInMem_lo_lo_lo_9};
  wire [63:0]      dataInMem_lo_hi_lo_lo_9 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9, dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [63:0]      dataInMem_lo_hi_lo_hi_9 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11, dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [127:0]     dataInMem_lo_hi_lo_9 = {dataInMem_lo_hi_lo_hi_9, dataInMem_lo_hi_lo_lo_9};
  wire [63:0]      dataInMem_lo_hi_hi_lo_9 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13, dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [63:0]      dataInMem_lo_hi_hi_hi_9 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15, dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [127:0]     dataInMem_lo_hi_hi_9 = {dataInMem_lo_hi_hi_hi_9, dataInMem_lo_hi_hi_lo_9};
  wire [255:0]     dataInMem_lo_hi_201 = {dataInMem_lo_hi_hi_9, dataInMem_lo_hi_lo_9};
  wire [511:0]     dataInMem_lo_329 = {dataInMem_lo_hi_201, dataInMem_lo_lo_73};
  wire [63:0]      dataInMem_hi_lo_lo_lo_9 = {dataRegroupBySew_1_1_17, dataRegroupBySew_0_1_17, dataRegroupBySew_1_1_16, dataRegroupBySew_0_1_16};
  wire [63:0]      dataInMem_hi_lo_lo_hi_9 = {dataRegroupBySew_1_1_19, dataRegroupBySew_0_1_19, dataRegroupBySew_1_1_18, dataRegroupBySew_0_1_18};
  wire [127:0]     dataInMem_hi_lo_lo_9 = {dataInMem_hi_lo_lo_hi_9, dataInMem_hi_lo_lo_lo_9};
  wire [63:0]      dataInMem_hi_lo_hi_lo_9 = {dataRegroupBySew_1_1_21, dataRegroupBySew_0_1_21, dataRegroupBySew_1_1_20, dataRegroupBySew_0_1_20};
  wire [63:0]      dataInMem_hi_lo_hi_hi_9 = {dataRegroupBySew_1_1_23, dataRegroupBySew_0_1_23, dataRegroupBySew_1_1_22, dataRegroupBySew_0_1_22};
  wire [127:0]     dataInMem_hi_lo_hi_9 = {dataInMem_hi_lo_hi_hi_9, dataInMem_hi_lo_hi_lo_9};
  wire [255:0]     dataInMem_hi_lo_137 = {dataInMem_hi_lo_hi_9, dataInMem_hi_lo_lo_9};
  wire [63:0]      dataInMem_hi_hi_lo_lo_9 = {dataRegroupBySew_1_1_25, dataRegroupBySew_0_1_25, dataRegroupBySew_1_1_24, dataRegroupBySew_0_1_24};
  wire [63:0]      dataInMem_hi_hi_lo_hi_9 = {dataRegroupBySew_1_1_27, dataRegroupBySew_0_1_27, dataRegroupBySew_1_1_26, dataRegroupBySew_0_1_26};
  wire [127:0]     dataInMem_hi_hi_lo_9 = {dataInMem_hi_hi_lo_hi_9, dataInMem_hi_hi_lo_lo_9};
  wire [63:0]      dataInMem_hi_hi_hi_lo_9 = {dataRegroupBySew_1_1_29, dataRegroupBySew_0_1_29, dataRegroupBySew_1_1_28, dataRegroupBySew_0_1_28};
  wire [63:0]      dataInMem_hi_hi_hi_hi_9 = {dataRegroupBySew_1_1_31, dataRegroupBySew_0_1_31, dataRegroupBySew_1_1_30, dataRegroupBySew_0_1_30};
  wire [127:0]     dataInMem_hi_hi_hi_9 = {dataInMem_hi_hi_hi_hi_9, dataInMem_hi_hi_hi_lo_9};
  wire [255:0]     dataInMem_hi_hi_265 = {dataInMem_hi_hi_hi_9, dataInMem_hi_hi_lo_9};
  wire [511:0]     dataInMem_hi_393 = {dataInMem_hi_hi_265, dataInMem_hi_lo_137};
  wire [1023:0]    dataInMem_9 = {dataInMem_hi_393, dataInMem_lo_329};
  wire [511:0]     regroupCacheLine_9_0 = dataInMem_9[511:0];
  wire [511:0]     regroupCacheLine_9_1 = dataInMem_9[1023:512];
  wire [511:0]     res_72 = regroupCacheLine_9_0;
  wire [511:0]     res_73 = regroupCacheLine_9_1;
  wire [1023:0]    lo_lo_9 = {res_73, res_72};
  wire [2047:0]    lo_9 = {1024'h0, lo_lo_9};
  wire [4095:0]    regroupLoadData_1_1 = {2048'h0, lo_9};
  wire [31:0]      _GEN_325 = {dataRegroupBySew_2_1_0, dataRegroupBySew_1_1_0};
  wire [31:0]      dataInMem_hi_394;
  assign dataInMem_hi_394 = _GEN_325;
  wire [31:0]      dataInMem_lo_hi_205;
  assign dataInMem_lo_hi_205 = _GEN_325;
  wire [31:0]      dataInMem_lo_hi_238;
  assign dataInMem_lo_hi_238 = _GEN_325;
  wire [31:0]      _GEN_326 = {dataRegroupBySew_2_1_1, dataRegroupBySew_1_1_1};
  wire [31:0]      dataInMem_hi_395;
  assign dataInMem_hi_395 = _GEN_326;
  wire [31:0]      dataInMem_lo_hi_206;
  assign dataInMem_lo_hi_206 = _GEN_326;
  wire [31:0]      dataInMem_lo_hi_239;
  assign dataInMem_lo_hi_239 = _GEN_326;
  wire [31:0]      _GEN_327 = {dataRegroupBySew_2_1_2, dataRegroupBySew_1_1_2};
  wire [31:0]      dataInMem_hi_396;
  assign dataInMem_hi_396 = _GEN_327;
  wire [31:0]      dataInMem_lo_hi_207;
  assign dataInMem_lo_hi_207 = _GEN_327;
  wire [31:0]      dataInMem_lo_hi_240;
  assign dataInMem_lo_hi_240 = _GEN_327;
  wire [31:0]      _GEN_328 = {dataRegroupBySew_2_1_3, dataRegroupBySew_1_1_3};
  wire [31:0]      dataInMem_hi_397;
  assign dataInMem_hi_397 = _GEN_328;
  wire [31:0]      dataInMem_lo_hi_208;
  assign dataInMem_lo_hi_208 = _GEN_328;
  wire [31:0]      dataInMem_lo_hi_241;
  assign dataInMem_lo_hi_241 = _GEN_328;
  wire [31:0]      _GEN_329 = {dataRegroupBySew_2_1_4, dataRegroupBySew_1_1_4};
  wire [31:0]      dataInMem_hi_398;
  assign dataInMem_hi_398 = _GEN_329;
  wire [31:0]      dataInMem_lo_hi_209;
  assign dataInMem_lo_hi_209 = _GEN_329;
  wire [31:0]      dataInMem_lo_hi_242;
  assign dataInMem_lo_hi_242 = _GEN_329;
  wire [31:0]      _GEN_330 = {dataRegroupBySew_2_1_5, dataRegroupBySew_1_1_5};
  wire [31:0]      dataInMem_hi_399;
  assign dataInMem_hi_399 = _GEN_330;
  wire [31:0]      dataInMem_lo_hi_210;
  assign dataInMem_lo_hi_210 = _GEN_330;
  wire [31:0]      dataInMem_lo_hi_243;
  assign dataInMem_lo_hi_243 = _GEN_330;
  wire [31:0]      _GEN_331 = {dataRegroupBySew_2_1_6, dataRegroupBySew_1_1_6};
  wire [31:0]      dataInMem_hi_400;
  assign dataInMem_hi_400 = _GEN_331;
  wire [31:0]      dataInMem_lo_hi_211;
  assign dataInMem_lo_hi_211 = _GEN_331;
  wire [31:0]      dataInMem_lo_hi_244;
  assign dataInMem_lo_hi_244 = _GEN_331;
  wire [31:0]      _GEN_332 = {dataRegroupBySew_2_1_7, dataRegroupBySew_1_1_7};
  wire [31:0]      dataInMem_hi_401;
  assign dataInMem_hi_401 = _GEN_332;
  wire [31:0]      dataInMem_lo_hi_212;
  assign dataInMem_lo_hi_212 = _GEN_332;
  wire [31:0]      dataInMem_lo_hi_245;
  assign dataInMem_lo_hi_245 = _GEN_332;
  wire [31:0]      _GEN_333 = {dataRegroupBySew_2_1_8, dataRegroupBySew_1_1_8};
  wire [31:0]      dataInMem_hi_402;
  assign dataInMem_hi_402 = _GEN_333;
  wire [31:0]      dataInMem_lo_hi_213;
  assign dataInMem_lo_hi_213 = _GEN_333;
  wire [31:0]      dataInMem_lo_hi_246;
  assign dataInMem_lo_hi_246 = _GEN_333;
  wire [31:0]      _GEN_334 = {dataRegroupBySew_2_1_9, dataRegroupBySew_1_1_9};
  wire [31:0]      dataInMem_hi_403;
  assign dataInMem_hi_403 = _GEN_334;
  wire [31:0]      dataInMem_lo_hi_214;
  assign dataInMem_lo_hi_214 = _GEN_334;
  wire [31:0]      dataInMem_lo_hi_247;
  assign dataInMem_lo_hi_247 = _GEN_334;
  wire [31:0]      _GEN_335 = {dataRegroupBySew_2_1_10, dataRegroupBySew_1_1_10};
  wire [31:0]      dataInMem_hi_404;
  assign dataInMem_hi_404 = _GEN_335;
  wire [31:0]      dataInMem_lo_hi_215;
  assign dataInMem_lo_hi_215 = _GEN_335;
  wire [31:0]      dataInMem_lo_hi_248;
  assign dataInMem_lo_hi_248 = _GEN_335;
  wire [31:0]      _GEN_336 = {dataRegroupBySew_2_1_11, dataRegroupBySew_1_1_11};
  wire [31:0]      dataInMem_hi_405;
  assign dataInMem_hi_405 = _GEN_336;
  wire [31:0]      dataInMem_lo_hi_216;
  assign dataInMem_lo_hi_216 = _GEN_336;
  wire [31:0]      dataInMem_lo_hi_249;
  assign dataInMem_lo_hi_249 = _GEN_336;
  wire [31:0]      _GEN_337 = {dataRegroupBySew_2_1_12, dataRegroupBySew_1_1_12};
  wire [31:0]      dataInMem_hi_406;
  assign dataInMem_hi_406 = _GEN_337;
  wire [31:0]      dataInMem_lo_hi_217;
  assign dataInMem_lo_hi_217 = _GEN_337;
  wire [31:0]      dataInMem_lo_hi_250;
  assign dataInMem_lo_hi_250 = _GEN_337;
  wire [31:0]      _GEN_338 = {dataRegroupBySew_2_1_13, dataRegroupBySew_1_1_13};
  wire [31:0]      dataInMem_hi_407;
  assign dataInMem_hi_407 = _GEN_338;
  wire [31:0]      dataInMem_lo_hi_218;
  assign dataInMem_lo_hi_218 = _GEN_338;
  wire [31:0]      dataInMem_lo_hi_251;
  assign dataInMem_lo_hi_251 = _GEN_338;
  wire [31:0]      _GEN_339 = {dataRegroupBySew_2_1_14, dataRegroupBySew_1_1_14};
  wire [31:0]      dataInMem_hi_408;
  assign dataInMem_hi_408 = _GEN_339;
  wire [31:0]      dataInMem_lo_hi_219;
  assign dataInMem_lo_hi_219 = _GEN_339;
  wire [31:0]      dataInMem_lo_hi_252;
  assign dataInMem_lo_hi_252 = _GEN_339;
  wire [31:0]      _GEN_340 = {dataRegroupBySew_2_1_15, dataRegroupBySew_1_1_15};
  wire [31:0]      dataInMem_hi_409;
  assign dataInMem_hi_409 = _GEN_340;
  wire [31:0]      dataInMem_lo_hi_220;
  assign dataInMem_lo_hi_220 = _GEN_340;
  wire [31:0]      dataInMem_lo_hi_253;
  assign dataInMem_lo_hi_253 = _GEN_340;
  wire [31:0]      _GEN_341 = {dataRegroupBySew_2_1_16, dataRegroupBySew_1_1_16};
  wire [31:0]      dataInMem_hi_410;
  assign dataInMem_hi_410 = _GEN_341;
  wire [31:0]      dataInMem_lo_hi_221;
  assign dataInMem_lo_hi_221 = _GEN_341;
  wire [31:0]      dataInMem_lo_hi_254;
  assign dataInMem_lo_hi_254 = _GEN_341;
  wire [31:0]      _GEN_342 = {dataRegroupBySew_2_1_17, dataRegroupBySew_1_1_17};
  wire [31:0]      dataInMem_hi_411;
  assign dataInMem_hi_411 = _GEN_342;
  wire [31:0]      dataInMem_lo_hi_222;
  assign dataInMem_lo_hi_222 = _GEN_342;
  wire [31:0]      dataInMem_lo_hi_255;
  assign dataInMem_lo_hi_255 = _GEN_342;
  wire [31:0]      _GEN_343 = {dataRegroupBySew_2_1_18, dataRegroupBySew_1_1_18};
  wire [31:0]      dataInMem_hi_412;
  assign dataInMem_hi_412 = _GEN_343;
  wire [31:0]      dataInMem_lo_hi_223;
  assign dataInMem_lo_hi_223 = _GEN_343;
  wire [31:0]      dataInMem_lo_hi_256;
  assign dataInMem_lo_hi_256 = _GEN_343;
  wire [31:0]      _GEN_344 = {dataRegroupBySew_2_1_19, dataRegroupBySew_1_1_19};
  wire [31:0]      dataInMem_hi_413;
  assign dataInMem_hi_413 = _GEN_344;
  wire [31:0]      dataInMem_lo_hi_224;
  assign dataInMem_lo_hi_224 = _GEN_344;
  wire [31:0]      dataInMem_lo_hi_257;
  assign dataInMem_lo_hi_257 = _GEN_344;
  wire [31:0]      _GEN_345 = {dataRegroupBySew_2_1_20, dataRegroupBySew_1_1_20};
  wire [31:0]      dataInMem_hi_414;
  assign dataInMem_hi_414 = _GEN_345;
  wire [31:0]      dataInMem_lo_hi_225;
  assign dataInMem_lo_hi_225 = _GEN_345;
  wire [31:0]      dataInMem_lo_hi_258;
  assign dataInMem_lo_hi_258 = _GEN_345;
  wire [31:0]      _GEN_346 = {dataRegroupBySew_2_1_21, dataRegroupBySew_1_1_21};
  wire [31:0]      dataInMem_hi_415;
  assign dataInMem_hi_415 = _GEN_346;
  wire [31:0]      dataInMem_lo_hi_226;
  assign dataInMem_lo_hi_226 = _GEN_346;
  wire [31:0]      dataInMem_lo_hi_259;
  assign dataInMem_lo_hi_259 = _GEN_346;
  wire [31:0]      _GEN_347 = {dataRegroupBySew_2_1_22, dataRegroupBySew_1_1_22};
  wire [31:0]      dataInMem_hi_416;
  assign dataInMem_hi_416 = _GEN_347;
  wire [31:0]      dataInMem_lo_hi_227;
  assign dataInMem_lo_hi_227 = _GEN_347;
  wire [31:0]      dataInMem_lo_hi_260;
  assign dataInMem_lo_hi_260 = _GEN_347;
  wire [31:0]      _GEN_348 = {dataRegroupBySew_2_1_23, dataRegroupBySew_1_1_23};
  wire [31:0]      dataInMem_hi_417;
  assign dataInMem_hi_417 = _GEN_348;
  wire [31:0]      dataInMem_lo_hi_228;
  assign dataInMem_lo_hi_228 = _GEN_348;
  wire [31:0]      dataInMem_lo_hi_261;
  assign dataInMem_lo_hi_261 = _GEN_348;
  wire [31:0]      _GEN_349 = {dataRegroupBySew_2_1_24, dataRegroupBySew_1_1_24};
  wire [31:0]      dataInMem_hi_418;
  assign dataInMem_hi_418 = _GEN_349;
  wire [31:0]      dataInMem_lo_hi_229;
  assign dataInMem_lo_hi_229 = _GEN_349;
  wire [31:0]      dataInMem_lo_hi_262;
  assign dataInMem_lo_hi_262 = _GEN_349;
  wire [31:0]      _GEN_350 = {dataRegroupBySew_2_1_25, dataRegroupBySew_1_1_25};
  wire [31:0]      dataInMem_hi_419;
  assign dataInMem_hi_419 = _GEN_350;
  wire [31:0]      dataInMem_lo_hi_230;
  assign dataInMem_lo_hi_230 = _GEN_350;
  wire [31:0]      dataInMem_lo_hi_263;
  assign dataInMem_lo_hi_263 = _GEN_350;
  wire [31:0]      _GEN_351 = {dataRegroupBySew_2_1_26, dataRegroupBySew_1_1_26};
  wire [31:0]      dataInMem_hi_420;
  assign dataInMem_hi_420 = _GEN_351;
  wire [31:0]      dataInMem_lo_hi_231;
  assign dataInMem_lo_hi_231 = _GEN_351;
  wire [31:0]      dataInMem_lo_hi_264;
  assign dataInMem_lo_hi_264 = _GEN_351;
  wire [31:0]      _GEN_352 = {dataRegroupBySew_2_1_27, dataRegroupBySew_1_1_27};
  wire [31:0]      dataInMem_hi_421;
  assign dataInMem_hi_421 = _GEN_352;
  wire [31:0]      dataInMem_lo_hi_232;
  assign dataInMem_lo_hi_232 = _GEN_352;
  wire [31:0]      dataInMem_lo_hi_265;
  assign dataInMem_lo_hi_265 = _GEN_352;
  wire [31:0]      _GEN_353 = {dataRegroupBySew_2_1_28, dataRegroupBySew_1_1_28};
  wire [31:0]      dataInMem_hi_422;
  assign dataInMem_hi_422 = _GEN_353;
  wire [31:0]      dataInMem_lo_hi_233;
  assign dataInMem_lo_hi_233 = _GEN_353;
  wire [31:0]      dataInMem_lo_hi_266;
  assign dataInMem_lo_hi_266 = _GEN_353;
  wire [31:0]      _GEN_354 = {dataRegroupBySew_2_1_29, dataRegroupBySew_1_1_29};
  wire [31:0]      dataInMem_hi_423;
  assign dataInMem_hi_423 = _GEN_354;
  wire [31:0]      dataInMem_lo_hi_234;
  assign dataInMem_lo_hi_234 = _GEN_354;
  wire [31:0]      dataInMem_lo_hi_267;
  assign dataInMem_lo_hi_267 = _GEN_354;
  wire [31:0]      _GEN_355 = {dataRegroupBySew_2_1_30, dataRegroupBySew_1_1_30};
  wire [31:0]      dataInMem_hi_424;
  assign dataInMem_hi_424 = _GEN_355;
  wire [31:0]      dataInMem_lo_hi_235;
  assign dataInMem_lo_hi_235 = _GEN_355;
  wire [31:0]      dataInMem_lo_hi_268;
  assign dataInMem_lo_hi_268 = _GEN_355;
  wire [31:0]      _GEN_356 = {dataRegroupBySew_2_1_31, dataRegroupBySew_1_1_31};
  wire [31:0]      dataInMem_hi_425;
  assign dataInMem_hi_425 = _GEN_356;
  wire [31:0]      dataInMem_lo_hi_236;
  assign dataInMem_lo_hi_236 = _GEN_356;
  wire [31:0]      dataInMem_lo_hi_269;
  assign dataInMem_lo_hi_269 = _GEN_356;
  wire [95:0]      dataInMem_lo_lo_lo_lo_10 = {dataInMem_hi_395, dataRegroupBySew_0_1_1, dataInMem_hi_394, dataRegroupBySew_0_1_0};
  wire [95:0]      dataInMem_lo_lo_lo_hi_10 = {dataInMem_hi_397, dataRegroupBySew_0_1_3, dataInMem_hi_396, dataRegroupBySew_0_1_2};
  wire [191:0]     dataInMem_lo_lo_lo_10 = {dataInMem_lo_lo_lo_hi_10, dataInMem_lo_lo_lo_lo_10};
  wire [95:0]      dataInMem_lo_lo_hi_lo_10 = {dataInMem_hi_399, dataRegroupBySew_0_1_5, dataInMem_hi_398, dataRegroupBySew_0_1_4};
  wire [95:0]      dataInMem_lo_lo_hi_hi_10 = {dataInMem_hi_401, dataRegroupBySew_0_1_7, dataInMem_hi_400, dataRegroupBySew_0_1_6};
  wire [191:0]     dataInMem_lo_lo_hi_10 = {dataInMem_lo_lo_hi_hi_10, dataInMem_lo_lo_hi_lo_10};
  wire [383:0]     dataInMem_lo_lo_74 = {dataInMem_lo_lo_hi_10, dataInMem_lo_lo_lo_10};
  wire [95:0]      dataInMem_lo_hi_lo_lo_10 = {dataInMem_hi_403, dataRegroupBySew_0_1_9, dataInMem_hi_402, dataRegroupBySew_0_1_8};
  wire [95:0]      dataInMem_lo_hi_lo_hi_10 = {dataInMem_hi_405, dataRegroupBySew_0_1_11, dataInMem_hi_404, dataRegroupBySew_0_1_10};
  wire [191:0]     dataInMem_lo_hi_lo_10 = {dataInMem_lo_hi_lo_hi_10, dataInMem_lo_hi_lo_lo_10};
  wire [95:0]      dataInMem_lo_hi_hi_lo_10 = {dataInMem_hi_407, dataRegroupBySew_0_1_13, dataInMem_hi_406, dataRegroupBySew_0_1_12};
  wire [95:0]      dataInMem_lo_hi_hi_hi_10 = {dataInMem_hi_409, dataRegroupBySew_0_1_15, dataInMem_hi_408, dataRegroupBySew_0_1_14};
  wire [191:0]     dataInMem_lo_hi_hi_10 = {dataInMem_lo_hi_hi_hi_10, dataInMem_lo_hi_hi_lo_10};
  wire [383:0]     dataInMem_lo_hi_202 = {dataInMem_lo_hi_hi_10, dataInMem_lo_hi_lo_10};
  wire [767:0]     dataInMem_lo_330 = {dataInMem_lo_hi_202, dataInMem_lo_lo_74};
  wire [95:0]      dataInMem_hi_lo_lo_lo_10 = {dataInMem_hi_411, dataRegroupBySew_0_1_17, dataInMem_hi_410, dataRegroupBySew_0_1_16};
  wire [95:0]      dataInMem_hi_lo_lo_hi_10 = {dataInMem_hi_413, dataRegroupBySew_0_1_19, dataInMem_hi_412, dataRegroupBySew_0_1_18};
  wire [191:0]     dataInMem_hi_lo_lo_10 = {dataInMem_hi_lo_lo_hi_10, dataInMem_hi_lo_lo_lo_10};
  wire [95:0]      dataInMem_hi_lo_hi_lo_10 = {dataInMem_hi_415, dataRegroupBySew_0_1_21, dataInMem_hi_414, dataRegroupBySew_0_1_20};
  wire [95:0]      dataInMem_hi_lo_hi_hi_10 = {dataInMem_hi_417, dataRegroupBySew_0_1_23, dataInMem_hi_416, dataRegroupBySew_0_1_22};
  wire [191:0]     dataInMem_hi_lo_hi_10 = {dataInMem_hi_lo_hi_hi_10, dataInMem_hi_lo_hi_lo_10};
  wire [383:0]     dataInMem_hi_lo_138 = {dataInMem_hi_lo_hi_10, dataInMem_hi_lo_lo_10};
  wire [95:0]      dataInMem_hi_hi_lo_lo_10 = {dataInMem_hi_419, dataRegroupBySew_0_1_25, dataInMem_hi_418, dataRegroupBySew_0_1_24};
  wire [95:0]      dataInMem_hi_hi_lo_hi_10 = {dataInMem_hi_421, dataRegroupBySew_0_1_27, dataInMem_hi_420, dataRegroupBySew_0_1_26};
  wire [191:0]     dataInMem_hi_hi_lo_10 = {dataInMem_hi_hi_lo_hi_10, dataInMem_hi_hi_lo_lo_10};
  wire [95:0]      dataInMem_hi_hi_hi_lo_10 = {dataInMem_hi_423, dataRegroupBySew_0_1_29, dataInMem_hi_422, dataRegroupBySew_0_1_28};
  wire [95:0]      dataInMem_hi_hi_hi_hi_10 = {dataInMem_hi_425, dataRegroupBySew_0_1_31, dataInMem_hi_424, dataRegroupBySew_0_1_30};
  wire [191:0]     dataInMem_hi_hi_hi_10 = {dataInMem_hi_hi_hi_hi_10, dataInMem_hi_hi_hi_lo_10};
  wire [383:0]     dataInMem_hi_hi_266 = {dataInMem_hi_hi_hi_10, dataInMem_hi_hi_lo_10};
  wire [767:0]     dataInMem_hi_426 = {dataInMem_hi_hi_266, dataInMem_hi_lo_138};
  wire [1535:0]    dataInMem_10 = {dataInMem_hi_426, dataInMem_lo_330};
  wire [511:0]     regroupCacheLine_10_0 = dataInMem_10[511:0];
  wire [511:0]     regroupCacheLine_10_1 = dataInMem_10[1023:512];
  wire [511:0]     regroupCacheLine_10_2 = dataInMem_10[1535:1024];
  wire [511:0]     res_80 = regroupCacheLine_10_0;
  wire [511:0]     res_81 = regroupCacheLine_10_1;
  wire [511:0]     res_82 = regroupCacheLine_10_2;
  wire [1023:0]    lo_lo_10 = {res_81, res_80};
  wire [1023:0]    lo_hi_10 = {512'h0, res_82};
  wire [2047:0]    lo_10 = {lo_hi_10, lo_lo_10};
  wire [4095:0]    regroupLoadData_1_2 = {2048'h0, lo_10};
  wire [31:0]      _GEN_357 = {dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_331;
  assign dataInMem_lo_331 = _GEN_357;
  wire [31:0]      dataInMem_lo_364;
  assign dataInMem_lo_364 = _GEN_357;
  wire [31:0]      dataInMem_lo_lo_79;
  assign dataInMem_lo_lo_79 = _GEN_357;
  wire [31:0]      _GEN_358 = {dataRegroupBySew_3_1_0, dataRegroupBySew_2_1_0};
  wire [31:0]      dataInMem_hi_427;
  assign dataInMem_hi_427 = _GEN_358;
  wire [31:0]      dataInMem_lo_hi_271;
  assign dataInMem_lo_hi_271 = _GEN_358;
  wire [31:0]      _GEN_359 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_lo_332;
  assign dataInMem_lo_332 = _GEN_359;
  wire [31:0]      dataInMem_lo_365;
  assign dataInMem_lo_365 = _GEN_359;
  wire [31:0]      dataInMem_lo_lo_80;
  assign dataInMem_lo_lo_80 = _GEN_359;
  wire [31:0]      _GEN_360 = {dataRegroupBySew_3_1_1, dataRegroupBySew_2_1_1};
  wire [31:0]      dataInMem_hi_428;
  assign dataInMem_hi_428 = _GEN_360;
  wire [31:0]      dataInMem_lo_hi_272;
  assign dataInMem_lo_hi_272 = _GEN_360;
  wire [31:0]      _GEN_361 = {dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_lo_333;
  assign dataInMem_lo_333 = _GEN_361;
  wire [31:0]      dataInMem_lo_366;
  assign dataInMem_lo_366 = _GEN_361;
  wire [31:0]      dataInMem_lo_lo_81;
  assign dataInMem_lo_lo_81 = _GEN_361;
  wire [31:0]      _GEN_362 = {dataRegroupBySew_3_1_2, dataRegroupBySew_2_1_2};
  wire [31:0]      dataInMem_hi_429;
  assign dataInMem_hi_429 = _GEN_362;
  wire [31:0]      dataInMem_lo_hi_273;
  assign dataInMem_lo_hi_273 = _GEN_362;
  wire [31:0]      _GEN_363 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_lo_334;
  assign dataInMem_lo_334 = _GEN_363;
  wire [31:0]      dataInMem_lo_367;
  assign dataInMem_lo_367 = _GEN_363;
  wire [31:0]      dataInMem_lo_lo_82;
  assign dataInMem_lo_lo_82 = _GEN_363;
  wire [31:0]      _GEN_364 = {dataRegroupBySew_3_1_3, dataRegroupBySew_2_1_3};
  wire [31:0]      dataInMem_hi_430;
  assign dataInMem_hi_430 = _GEN_364;
  wire [31:0]      dataInMem_lo_hi_274;
  assign dataInMem_lo_hi_274 = _GEN_364;
  wire [31:0]      _GEN_365 = {dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_lo_335;
  assign dataInMem_lo_335 = _GEN_365;
  wire [31:0]      dataInMem_lo_368;
  assign dataInMem_lo_368 = _GEN_365;
  wire [31:0]      dataInMem_lo_lo_83;
  assign dataInMem_lo_lo_83 = _GEN_365;
  wire [31:0]      _GEN_366 = {dataRegroupBySew_3_1_4, dataRegroupBySew_2_1_4};
  wire [31:0]      dataInMem_hi_431;
  assign dataInMem_hi_431 = _GEN_366;
  wire [31:0]      dataInMem_lo_hi_275;
  assign dataInMem_lo_hi_275 = _GEN_366;
  wire [31:0]      _GEN_367 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_lo_336;
  assign dataInMem_lo_336 = _GEN_367;
  wire [31:0]      dataInMem_lo_369;
  assign dataInMem_lo_369 = _GEN_367;
  wire [31:0]      dataInMem_lo_lo_84;
  assign dataInMem_lo_lo_84 = _GEN_367;
  wire [31:0]      _GEN_368 = {dataRegroupBySew_3_1_5, dataRegroupBySew_2_1_5};
  wire [31:0]      dataInMem_hi_432;
  assign dataInMem_hi_432 = _GEN_368;
  wire [31:0]      dataInMem_lo_hi_276;
  assign dataInMem_lo_hi_276 = _GEN_368;
  wire [31:0]      _GEN_369 = {dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_lo_337;
  assign dataInMem_lo_337 = _GEN_369;
  wire [31:0]      dataInMem_lo_370;
  assign dataInMem_lo_370 = _GEN_369;
  wire [31:0]      dataInMem_lo_lo_85;
  assign dataInMem_lo_lo_85 = _GEN_369;
  wire [31:0]      _GEN_370 = {dataRegroupBySew_3_1_6, dataRegroupBySew_2_1_6};
  wire [31:0]      dataInMem_hi_433;
  assign dataInMem_hi_433 = _GEN_370;
  wire [31:0]      dataInMem_lo_hi_277;
  assign dataInMem_lo_hi_277 = _GEN_370;
  wire [31:0]      _GEN_371 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_lo_338;
  assign dataInMem_lo_338 = _GEN_371;
  wire [31:0]      dataInMem_lo_371;
  assign dataInMem_lo_371 = _GEN_371;
  wire [31:0]      dataInMem_lo_lo_86;
  assign dataInMem_lo_lo_86 = _GEN_371;
  wire [31:0]      _GEN_372 = {dataRegroupBySew_3_1_7, dataRegroupBySew_2_1_7};
  wire [31:0]      dataInMem_hi_434;
  assign dataInMem_hi_434 = _GEN_372;
  wire [31:0]      dataInMem_lo_hi_278;
  assign dataInMem_lo_hi_278 = _GEN_372;
  wire [31:0]      _GEN_373 = {dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_lo_339;
  assign dataInMem_lo_339 = _GEN_373;
  wire [31:0]      dataInMem_lo_372;
  assign dataInMem_lo_372 = _GEN_373;
  wire [31:0]      dataInMem_lo_lo_87;
  assign dataInMem_lo_lo_87 = _GEN_373;
  wire [31:0]      _GEN_374 = {dataRegroupBySew_3_1_8, dataRegroupBySew_2_1_8};
  wire [31:0]      dataInMem_hi_435;
  assign dataInMem_hi_435 = _GEN_374;
  wire [31:0]      dataInMem_lo_hi_279;
  assign dataInMem_lo_hi_279 = _GEN_374;
  wire [31:0]      _GEN_375 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9};
  wire [31:0]      dataInMem_lo_340;
  assign dataInMem_lo_340 = _GEN_375;
  wire [31:0]      dataInMem_lo_373;
  assign dataInMem_lo_373 = _GEN_375;
  wire [31:0]      dataInMem_lo_lo_88;
  assign dataInMem_lo_lo_88 = _GEN_375;
  wire [31:0]      _GEN_376 = {dataRegroupBySew_3_1_9, dataRegroupBySew_2_1_9};
  wire [31:0]      dataInMem_hi_436;
  assign dataInMem_hi_436 = _GEN_376;
  wire [31:0]      dataInMem_lo_hi_280;
  assign dataInMem_lo_hi_280 = _GEN_376;
  wire [31:0]      _GEN_377 = {dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [31:0]      dataInMem_lo_341;
  assign dataInMem_lo_341 = _GEN_377;
  wire [31:0]      dataInMem_lo_374;
  assign dataInMem_lo_374 = _GEN_377;
  wire [31:0]      dataInMem_lo_lo_89;
  assign dataInMem_lo_lo_89 = _GEN_377;
  wire [31:0]      _GEN_378 = {dataRegroupBySew_3_1_10, dataRegroupBySew_2_1_10};
  wire [31:0]      dataInMem_hi_437;
  assign dataInMem_hi_437 = _GEN_378;
  wire [31:0]      dataInMem_lo_hi_281;
  assign dataInMem_lo_hi_281 = _GEN_378;
  wire [31:0]      _GEN_379 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11};
  wire [31:0]      dataInMem_lo_342;
  assign dataInMem_lo_342 = _GEN_379;
  wire [31:0]      dataInMem_lo_375;
  assign dataInMem_lo_375 = _GEN_379;
  wire [31:0]      dataInMem_lo_lo_90;
  assign dataInMem_lo_lo_90 = _GEN_379;
  wire [31:0]      _GEN_380 = {dataRegroupBySew_3_1_11, dataRegroupBySew_2_1_11};
  wire [31:0]      dataInMem_hi_438;
  assign dataInMem_hi_438 = _GEN_380;
  wire [31:0]      dataInMem_lo_hi_282;
  assign dataInMem_lo_hi_282 = _GEN_380;
  wire [31:0]      _GEN_381 = {dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_lo_343;
  assign dataInMem_lo_343 = _GEN_381;
  wire [31:0]      dataInMem_lo_376;
  assign dataInMem_lo_376 = _GEN_381;
  wire [31:0]      dataInMem_lo_lo_91;
  assign dataInMem_lo_lo_91 = _GEN_381;
  wire [31:0]      _GEN_382 = {dataRegroupBySew_3_1_12, dataRegroupBySew_2_1_12};
  wire [31:0]      dataInMem_hi_439;
  assign dataInMem_hi_439 = _GEN_382;
  wire [31:0]      dataInMem_lo_hi_283;
  assign dataInMem_lo_hi_283 = _GEN_382;
  wire [31:0]      _GEN_383 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13};
  wire [31:0]      dataInMem_lo_344;
  assign dataInMem_lo_344 = _GEN_383;
  wire [31:0]      dataInMem_lo_377;
  assign dataInMem_lo_377 = _GEN_383;
  wire [31:0]      dataInMem_lo_lo_92;
  assign dataInMem_lo_lo_92 = _GEN_383;
  wire [31:0]      _GEN_384 = {dataRegroupBySew_3_1_13, dataRegroupBySew_2_1_13};
  wire [31:0]      dataInMem_hi_440;
  assign dataInMem_hi_440 = _GEN_384;
  wire [31:0]      dataInMem_lo_hi_284;
  assign dataInMem_lo_hi_284 = _GEN_384;
  wire [31:0]      _GEN_385 = {dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [31:0]      dataInMem_lo_345;
  assign dataInMem_lo_345 = _GEN_385;
  wire [31:0]      dataInMem_lo_378;
  assign dataInMem_lo_378 = _GEN_385;
  wire [31:0]      dataInMem_lo_lo_93;
  assign dataInMem_lo_lo_93 = _GEN_385;
  wire [31:0]      _GEN_386 = {dataRegroupBySew_3_1_14, dataRegroupBySew_2_1_14};
  wire [31:0]      dataInMem_hi_441;
  assign dataInMem_hi_441 = _GEN_386;
  wire [31:0]      dataInMem_lo_hi_285;
  assign dataInMem_lo_hi_285 = _GEN_386;
  wire [31:0]      _GEN_387 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15};
  wire [31:0]      dataInMem_lo_346;
  assign dataInMem_lo_346 = _GEN_387;
  wire [31:0]      dataInMem_lo_379;
  assign dataInMem_lo_379 = _GEN_387;
  wire [31:0]      dataInMem_lo_lo_94;
  assign dataInMem_lo_lo_94 = _GEN_387;
  wire [31:0]      _GEN_388 = {dataRegroupBySew_3_1_15, dataRegroupBySew_2_1_15};
  wire [31:0]      dataInMem_hi_442;
  assign dataInMem_hi_442 = _GEN_388;
  wire [31:0]      dataInMem_lo_hi_286;
  assign dataInMem_lo_hi_286 = _GEN_388;
  wire [31:0]      _GEN_389 = {dataRegroupBySew_1_1_16, dataRegroupBySew_0_1_16};
  wire [31:0]      dataInMem_lo_347;
  assign dataInMem_lo_347 = _GEN_389;
  wire [31:0]      dataInMem_lo_380;
  assign dataInMem_lo_380 = _GEN_389;
  wire [31:0]      dataInMem_lo_lo_95;
  assign dataInMem_lo_lo_95 = _GEN_389;
  wire [31:0]      _GEN_390 = {dataRegroupBySew_3_1_16, dataRegroupBySew_2_1_16};
  wire [31:0]      dataInMem_hi_443;
  assign dataInMem_hi_443 = _GEN_390;
  wire [31:0]      dataInMem_lo_hi_287;
  assign dataInMem_lo_hi_287 = _GEN_390;
  wire [31:0]      _GEN_391 = {dataRegroupBySew_1_1_17, dataRegroupBySew_0_1_17};
  wire [31:0]      dataInMem_lo_348;
  assign dataInMem_lo_348 = _GEN_391;
  wire [31:0]      dataInMem_lo_381;
  assign dataInMem_lo_381 = _GEN_391;
  wire [31:0]      dataInMem_lo_lo_96;
  assign dataInMem_lo_lo_96 = _GEN_391;
  wire [31:0]      _GEN_392 = {dataRegroupBySew_3_1_17, dataRegroupBySew_2_1_17};
  wire [31:0]      dataInMem_hi_444;
  assign dataInMem_hi_444 = _GEN_392;
  wire [31:0]      dataInMem_lo_hi_288;
  assign dataInMem_lo_hi_288 = _GEN_392;
  wire [31:0]      _GEN_393 = {dataRegroupBySew_1_1_18, dataRegroupBySew_0_1_18};
  wire [31:0]      dataInMem_lo_349;
  assign dataInMem_lo_349 = _GEN_393;
  wire [31:0]      dataInMem_lo_382;
  assign dataInMem_lo_382 = _GEN_393;
  wire [31:0]      dataInMem_lo_lo_97;
  assign dataInMem_lo_lo_97 = _GEN_393;
  wire [31:0]      _GEN_394 = {dataRegroupBySew_3_1_18, dataRegroupBySew_2_1_18};
  wire [31:0]      dataInMem_hi_445;
  assign dataInMem_hi_445 = _GEN_394;
  wire [31:0]      dataInMem_lo_hi_289;
  assign dataInMem_lo_hi_289 = _GEN_394;
  wire [31:0]      _GEN_395 = {dataRegroupBySew_1_1_19, dataRegroupBySew_0_1_19};
  wire [31:0]      dataInMem_lo_350;
  assign dataInMem_lo_350 = _GEN_395;
  wire [31:0]      dataInMem_lo_383;
  assign dataInMem_lo_383 = _GEN_395;
  wire [31:0]      dataInMem_lo_lo_98;
  assign dataInMem_lo_lo_98 = _GEN_395;
  wire [31:0]      _GEN_396 = {dataRegroupBySew_3_1_19, dataRegroupBySew_2_1_19};
  wire [31:0]      dataInMem_hi_446;
  assign dataInMem_hi_446 = _GEN_396;
  wire [31:0]      dataInMem_lo_hi_290;
  assign dataInMem_lo_hi_290 = _GEN_396;
  wire [31:0]      _GEN_397 = {dataRegroupBySew_1_1_20, dataRegroupBySew_0_1_20};
  wire [31:0]      dataInMem_lo_351;
  assign dataInMem_lo_351 = _GEN_397;
  wire [31:0]      dataInMem_lo_384;
  assign dataInMem_lo_384 = _GEN_397;
  wire [31:0]      dataInMem_lo_lo_99;
  assign dataInMem_lo_lo_99 = _GEN_397;
  wire [31:0]      _GEN_398 = {dataRegroupBySew_3_1_20, dataRegroupBySew_2_1_20};
  wire [31:0]      dataInMem_hi_447;
  assign dataInMem_hi_447 = _GEN_398;
  wire [31:0]      dataInMem_lo_hi_291;
  assign dataInMem_lo_hi_291 = _GEN_398;
  wire [31:0]      _GEN_399 = {dataRegroupBySew_1_1_21, dataRegroupBySew_0_1_21};
  wire [31:0]      dataInMem_lo_352;
  assign dataInMem_lo_352 = _GEN_399;
  wire [31:0]      dataInMem_lo_385;
  assign dataInMem_lo_385 = _GEN_399;
  wire [31:0]      dataInMem_lo_lo_100;
  assign dataInMem_lo_lo_100 = _GEN_399;
  wire [31:0]      _GEN_400 = {dataRegroupBySew_3_1_21, dataRegroupBySew_2_1_21};
  wire [31:0]      dataInMem_hi_448;
  assign dataInMem_hi_448 = _GEN_400;
  wire [31:0]      dataInMem_lo_hi_292;
  assign dataInMem_lo_hi_292 = _GEN_400;
  wire [31:0]      _GEN_401 = {dataRegroupBySew_1_1_22, dataRegroupBySew_0_1_22};
  wire [31:0]      dataInMem_lo_353;
  assign dataInMem_lo_353 = _GEN_401;
  wire [31:0]      dataInMem_lo_386;
  assign dataInMem_lo_386 = _GEN_401;
  wire [31:0]      dataInMem_lo_lo_101;
  assign dataInMem_lo_lo_101 = _GEN_401;
  wire [31:0]      _GEN_402 = {dataRegroupBySew_3_1_22, dataRegroupBySew_2_1_22};
  wire [31:0]      dataInMem_hi_449;
  assign dataInMem_hi_449 = _GEN_402;
  wire [31:0]      dataInMem_lo_hi_293;
  assign dataInMem_lo_hi_293 = _GEN_402;
  wire [31:0]      _GEN_403 = {dataRegroupBySew_1_1_23, dataRegroupBySew_0_1_23};
  wire [31:0]      dataInMem_lo_354;
  assign dataInMem_lo_354 = _GEN_403;
  wire [31:0]      dataInMem_lo_387;
  assign dataInMem_lo_387 = _GEN_403;
  wire [31:0]      dataInMem_lo_lo_102;
  assign dataInMem_lo_lo_102 = _GEN_403;
  wire [31:0]      _GEN_404 = {dataRegroupBySew_3_1_23, dataRegroupBySew_2_1_23};
  wire [31:0]      dataInMem_hi_450;
  assign dataInMem_hi_450 = _GEN_404;
  wire [31:0]      dataInMem_lo_hi_294;
  assign dataInMem_lo_hi_294 = _GEN_404;
  wire [31:0]      _GEN_405 = {dataRegroupBySew_1_1_24, dataRegroupBySew_0_1_24};
  wire [31:0]      dataInMem_lo_355;
  assign dataInMem_lo_355 = _GEN_405;
  wire [31:0]      dataInMem_lo_388;
  assign dataInMem_lo_388 = _GEN_405;
  wire [31:0]      dataInMem_lo_lo_103;
  assign dataInMem_lo_lo_103 = _GEN_405;
  wire [31:0]      _GEN_406 = {dataRegroupBySew_3_1_24, dataRegroupBySew_2_1_24};
  wire [31:0]      dataInMem_hi_451;
  assign dataInMem_hi_451 = _GEN_406;
  wire [31:0]      dataInMem_lo_hi_295;
  assign dataInMem_lo_hi_295 = _GEN_406;
  wire [31:0]      _GEN_407 = {dataRegroupBySew_1_1_25, dataRegroupBySew_0_1_25};
  wire [31:0]      dataInMem_lo_356;
  assign dataInMem_lo_356 = _GEN_407;
  wire [31:0]      dataInMem_lo_389;
  assign dataInMem_lo_389 = _GEN_407;
  wire [31:0]      dataInMem_lo_lo_104;
  assign dataInMem_lo_lo_104 = _GEN_407;
  wire [31:0]      _GEN_408 = {dataRegroupBySew_3_1_25, dataRegroupBySew_2_1_25};
  wire [31:0]      dataInMem_hi_452;
  assign dataInMem_hi_452 = _GEN_408;
  wire [31:0]      dataInMem_lo_hi_296;
  assign dataInMem_lo_hi_296 = _GEN_408;
  wire [31:0]      _GEN_409 = {dataRegroupBySew_1_1_26, dataRegroupBySew_0_1_26};
  wire [31:0]      dataInMem_lo_357;
  assign dataInMem_lo_357 = _GEN_409;
  wire [31:0]      dataInMem_lo_390;
  assign dataInMem_lo_390 = _GEN_409;
  wire [31:0]      dataInMem_lo_lo_105;
  assign dataInMem_lo_lo_105 = _GEN_409;
  wire [31:0]      _GEN_410 = {dataRegroupBySew_3_1_26, dataRegroupBySew_2_1_26};
  wire [31:0]      dataInMem_hi_453;
  assign dataInMem_hi_453 = _GEN_410;
  wire [31:0]      dataInMem_lo_hi_297;
  assign dataInMem_lo_hi_297 = _GEN_410;
  wire [31:0]      _GEN_411 = {dataRegroupBySew_1_1_27, dataRegroupBySew_0_1_27};
  wire [31:0]      dataInMem_lo_358;
  assign dataInMem_lo_358 = _GEN_411;
  wire [31:0]      dataInMem_lo_391;
  assign dataInMem_lo_391 = _GEN_411;
  wire [31:0]      dataInMem_lo_lo_106;
  assign dataInMem_lo_lo_106 = _GEN_411;
  wire [31:0]      _GEN_412 = {dataRegroupBySew_3_1_27, dataRegroupBySew_2_1_27};
  wire [31:0]      dataInMem_hi_454;
  assign dataInMem_hi_454 = _GEN_412;
  wire [31:0]      dataInMem_lo_hi_298;
  assign dataInMem_lo_hi_298 = _GEN_412;
  wire [31:0]      _GEN_413 = {dataRegroupBySew_1_1_28, dataRegroupBySew_0_1_28};
  wire [31:0]      dataInMem_lo_359;
  assign dataInMem_lo_359 = _GEN_413;
  wire [31:0]      dataInMem_lo_392;
  assign dataInMem_lo_392 = _GEN_413;
  wire [31:0]      dataInMem_lo_lo_107;
  assign dataInMem_lo_lo_107 = _GEN_413;
  wire [31:0]      _GEN_414 = {dataRegroupBySew_3_1_28, dataRegroupBySew_2_1_28};
  wire [31:0]      dataInMem_hi_455;
  assign dataInMem_hi_455 = _GEN_414;
  wire [31:0]      dataInMem_lo_hi_299;
  assign dataInMem_lo_hi_299 = _GEN_414;
  wire [31:0]      _GEN_415 = {dataRegroupBySew_1_1_29, dataRegroupBySew_0_1_29};
  wire [31:0]      dataInMem_lo_360;
  assign dataInMem_lo_360 = _GEN_415;
  wire [31:0]      dataInMem_lo_393;
  assign dataInMem_lo_393 = _GEN_415;
  wire [31:0]      dataInMem_lo_lo_108;
  assign dataInMem_lo_lo_108 = _GEN_415;
  wire [31:0]      _GEN_416 = {dataRegroupBySew_3_1_29, dataRegroupBySew_2_1_29};
  wire [31:0]      dataInMem_hi_456;
  assign dataInMem_hi_456 = _GEN_416;
  wire [31:0]      dataInMem_lo_hi_300;
  assign dataInMem_lo_hi_300 = _GEN_416;
  wire [31:0]      _GEN_417 = {dataRegroupBySew_1_1_30, dataRegroupBySew_0_1_30};
  wire [31:0]      dataInMem_lo_361;
  assign dataInMem_lo_361 = _GEN_417;
  wire [31:0]      dataInMem_lo_394;
  assign dataInMem_lo_394 = _GEN_417;
  wire [31:0]      dataInMem_lo_lo_109;
  assign dataInMem_lo_lo_109 = _GEN_417;
  wire [31:0]      _GEN_418 = {dataRegroupBySew_3_1_30, dataRegroupBySew_2_1_30};
  wire [31:0]      dataInMem_hi_457;
  assign dataInMem_hi_457 = _GEN_418;
  wire [31:0]      dataInMem_lo_hi_301;
  assign dataInMem_lo_hi_301 = _GEN_418;
  wire [31:0]      _GEN_419 = {dataRegroupBySew_1_1_31, dataRegroupBySew_0_1_31};
  wire [31:0]      dataInMem_lo_362;
  assign dataInMem_lo_362 = _GEN_419;
  wire [31:0]      dataInMem_lo_395;
  assign dataInMem_lo_395 = _GEN_419;
  wire [31:0]      dataInMem_lo_lo_110;
  assign dataInMem_lo_lo_110 = _GEN_419;
  wire [31:0]      _GEN_420 = {dataRegroupBySew_3_1_31, dataRegroupBySew_2_1_31};
  wire [31:0]      dataInMem_hi_458;
  assign dataInMem_hi_458 = _GEN_420;
  wire [31:0]      dataInMem_lo_hi_302;
  assign dataInMem_lo_hi_302 = _GEN_420;
  wire [127:0]     dataInMem_lo_lo_lo_lo_11 = {dataInMem_hi_428, dataInMem_lo_332, dataInMem_hi_427, dataInMem_lo_331};
  wire [127:0]     dataInMem_lo_lo_lo_hi_11 = {dataInMem_hi_430, dataInMem_lo_334, dataInMem_hi_429, dataInMem_lo_333};
  wire [255:0]     dataInMem_lo_lo_lo_11 = {dataInMem_lo_lo_lo_hi_11, dataInMem_lo_lo_lo_lo_11};
  wire [127:0]     dataInMem_lo_lo_hi_lo_11 = {dataInMem_hi_432, dataInMem_lo_336, dataInMem_hi_431, dataInMem_lo_335};
  wire [127:0]     dataInMem_lo_lo_hi_hi_11 = {dataInMem_hi_434, dataInMem_lo_338, dataInMem_hi_433, dataInMem_lo_337};
  wire [255:0]     dataInMem_lo_lo_hi_11 = {dataInMem_lo_lo_hi_hi_11, dataInMem_lo_lo_hi_lo_11};
  wire [511:0]     dataInMem_lo_lo_75 = {dataInMem_lo_lo_hi_11, dataInMem_lo_lo_lo_11};
  wire [127:0]     dataInMem_lo_hi_lo_lo_11 = {dataInMem_hi_436, dataInMem_lo_340, dataInMem_hi_435, dataInMem_lo_339};
  wire [127:0]     dataInMem_lo_hi_lo_hi_11 = {dataInMem_hi_438, dataInMem_lo_342, dataInMem_hi_437, dataInMem_lo_341};
  wire [255:0]     dataInMem_lo_hi_lo_11 = {dataInMem_lo_hi_lo_hi_11, dataInMem_lo_hi_lo_lo_11};
  wire [127:0]     dataInMem_lo_hi_hi_lo_11 = {dataInMem_hi_440, dataInMem_lo_344, dataInMem_hi_439, dataInMem_lo_343};
  wire [127:0]     dataInMem_lo_hi_hi_hi_11 = {dataInMem_hi_442, dataInMem_lo_346, dataInMem_hi_441, dataInMem_lo_345};
  wire [255:0]     dataInMem_lo_hi_hi_11 = {dataInMem_lo_hi_hi_hi_11, dataInMem_lo_hi_hi_lo_11};
  wire [511:0]     dataInMem_lo_hi_203 = {dataInMem_lo_hi_hi_11, dataInMem_lo_hi_lo_11};
  wire [1023:0]    dataInMem_lo_363 = {dataInMem_lo_hi_203, dataInMem_lo_lo_75};
  wire [127:0]     dataInMem_hi_lo_lo_lo_11 = {dataInMem_hi_444, dataInMem_lo_348, dataInMem_hi_443, dataInMem_lo_347};
  wire [127:0]     dataInMem_hi_lo_lo_hi_11 = {dataInMem_hi_446, dataInMem_lo_350, dataInMem_hi_445, dataInMem_lo_349};
  wire [255:0]     dataInMem_hi_lo_lo_11 = {dataInMem_hi_lo_lo_hi_11, dataInMem_hi_lo_lo_lo_11};
  wire [127:0]     dataInMem_hi_lo_hi_lo_11 = {dataInMem_hi_448, dataInMem_lo_352, dataInMem_hi_447, dataInMem_lo_351};
  wire [127:0]     dataInMem_hi_lo_hi_hi_11 = {dataInMem_hi_450, dataInMem_lo_354, dataInMem_hi_449, dataInMem_lo_353};
  wire [255:0]     dataInMem_hi_lo_hi_11 = {dataInMem_hi_lo_hi_hi_11, dataInMem_hi_lo_hi_lo_11};
  wire [511:0]     dataInMem_hi_lo_139 = {dataInMem_hi_lo_hi_11, dataInMem_hi_lo_lo_11};
  wire [127:0]     dataInMem_hi_hi_lo_lo_11 = {dataInMem_hi_452, dataInMem_lo_356, dataInMem_hi_451, dataInMem_lo_355};
  wire [127:0]     dataInMem_hi_hi_lo_hi_11 = {dataInMem_hi_454, dataInMem_lo_358, dataInMem_hi_453, dataInMem_lo_357};
  wire [255:0]     dataInMem_hi_hi_lo_11 = {dataInMem_hi_hi_lo_hi_11, dataInMem_hi_hi_lo_lo_11};
  wire [127:0]     dataInMem_hi_hi_hi_lo_11 = {dataInMem_hi_456, dataInMem_lo_360, dataInMem_hi_455, dataInMem_lo_359};
  wire [127:0]     dataInMem_hi_hi_hi_hi_11 = {dataInMem_hi_458, dataInMem_lo_362, dataInMem_hi_457, dataInMem_lo_361};
  wire [255:0]     dataInMem_hi_hi_hi_11 = {dataInMem_hi_hi_hi_hi_11, dataInMem_hi_hi_hi_lo_11};
  wire [511:0]     dataInMem_hi_hi_267 = {dataInMem_hi_hi_hi_11, dataInMem_hi_hi_lo_11};
  wire [1023:0]    dataInMem_hi_459 = {dataInMem_hi_hi_267, dataInMem_hi_lo_139};
  wire [2047:0]    dataInMem_11 = {dataInMem_hi_459, dataInMem_lo_363};
  wire [511:0]     regroupCacheLine_11_0 = dataInMem_11[511:0];
  wire [511:0]     regroupCacheLine_11_1 = dataInMem_11[1023:512];
  wire [511:0]     regroupCacheLine_11_2 = dataInMem_11[1535:1024];
  wire [511:0]     regroupCacheLine_11_3 = dataInMem_11[2047:1536];
  wire [511:0]     res_88 = regroupCacheLine_11_0;
  wire [511:0]     res_89 = regroupCacheLine_11_1;
  wire [511:0]     res_90 = regroupCacheLine_11_2;
  wire [511:0]     res_91 = regroupCacheLine_11_3;
  wire [1023:0]    lo_lo_11 = {res_89, res_88};
  wire [1023:0]    lo_hi_11 = {res_91, res_90};
  wire [2047:0]    lo_11 = {lo_hi_11, lo_lo_11};
  wire [4095:0]    regroupLoadData_1_3 = {2048'h0, lo_11};
  wire [31:0]      _GEN_421 = {dataRegroupBySew_4_1_0, dataRegroupBySew_3_1_0};
  wire [31:0]      dataInMem_hi_hi_268;
  assign dataInMem_hi_hi_268 = _GEN_421;
  wire [31:0]      dataInMem_hi_lo_142;
  assign dataInMem_hi_lo_142 = _GEN_421;
  wire [47:0]      dataInMem_hi_460 = {dataInMem_hi_hi_268, dataRegroupBySew_2_1_0};
  wire [31:0]      _GEN_422 = {dataRegroupBySew_4_1_1, dataRegroupBySew_3_1_1};
  wire [31:0]      dataInMem_hi_hi_269;
  assign dataInMem_hi_hi_269 = _GEN_422;
  wire [31:0]      dataInMem_hi_lo_143;
  assign dataInMem_hi_lo_143 = _GEN_422;
  wire [47:0]      dataInMem_hi_461 = {dataInMem_hi_hi_269, dataRegroupBySew_2_1_1};
  wire [31:0]      _GEN_423 = {dataRegroupBySew_4_1_2, dataRegroupBySew_3_1_2};
  wire [31:0]      dataInMem_hi_hi_270;
  assign dataInMem_hi_hi_270 = _GEN_423;
  wire [31:0]      dataInMem_hi_lo_144;
  assign dataInMem_hi_lo_144 = _GEN_423;
  wire [47:0]      dataInMem_hi_462 = {dataInMem_hi_hi_270, dataRegroupBySew_2_1_2};
  wire [31:0]      _GEN_424 = {dataRegroupBySew_4_1_3, dataRegroupBySew_3_1_3};
  wire [31:0]      dataInMem_hi_hi_271;
  assign dataInMem_hi_hi_271 = _GEN_424;
  wire [31:0]      dataInMem_hi_lo_145;
  assign dataInMem_hi_lo_145 = _GEN_424;
  wire [47:0]      dataInMem_hi_463 = {dataInMem_hi_hi_271, dataRegroupBySew_2_1_3};
  wire [31:0]      _GEN_425 = {dataRegroupBySew_4_1_4, dataRegroupBySew_3_1_4};
  wire [31:0]      dataInMem_hi_hi_272;
  assign dataInMem_hi_hi_272 = _GEN_425;
  wire [31:0]      dataInMem_hi_lo_146;
  assign dataInMem_hi_lo_146 = _GEN_425;
  wire [47:0]      dataInMem_hi_464 = {dataInMem_hi_hi_272, dataRegroupBySew_2_1_4};
  wire [31:0]      _GEN_426 = {dataRegroupBySew_4_1_5, dataRegroupBySew_3_1_5};
  wire [31:0]      dataInMem_hi_hi_273;
  assign dataInMem_hi_hi_273 = _GEN_426;
  wire [31:0]      dataInMem_hi_lo_147;
  assign dataInMem_hi_lo_147 = _GEN_426;
  wire [47:0]      dataInMem_hi_465 = {dataInMem_hi_hi_273, dataRegroupBySew_2_1_5};
  wire [31:0]      _GEN_427 = {dataRegroupBySew_4_1_6, dataRegroupBySew_3_1_6};
  wire [31:0]      dataInMem_hi_hi_274;
  assign dataInMem_hi_hi_274 = _GEN_427;
  wire [31:0]      dataInMem_hi_lo_148;
  assign dataInMem_hi_lo_148 = _GEN_427;
  wire [47:0]      dataInMem_hi_466 = {dataInMem_hi_hi_274, dataRegroupBySew_2_1_6};
  wire [31:0]      _GEN_428 = {dataRegroupBySew_4_1_7, dataRegroupBySew_3_1_7};
  wire [31:0]      dataInMem_hi_hi_275;
  assign dataInMem_hi_hi_275 = _GEN_428;
  wire [31:0]      dataInMem_hi_lo_149;
  assign dataInMem_hi_lo_149 = _GEN_428;
  wire [47:0]      dataInMem_hi_467 = {dataInMem_hi_hi_275, dataRegroupBySew_2_1_7};
  wire [31:0]      _GEN_429 = {dataRegroupBySew_4_1_8, dataRegroupBySew_3_1_8};
  wire [31:0]      dataInMem_hi_hi_276;
  assign dataInMem_hi_hi_276 = _GEN_429;
  wire [31:0]      dataInMem_hi_lo_150;
  assign dataInMem_hi_lo_150 = _GEN_429;
  wire [47:0]      dataInMem_hi_468 = {dataInMem_hi_hi_276, dataRegroupBySew_2_1_8};
  wire [31:0]      _GEN_430 = {dataRegroupBySew_4_1_9, dataRegroupBySew_3_1_9};
  wire [31:0]      dataInMem_hi_hi_277;
  assign dataInMem_hi_hi_277 = _GEN_430;
  wire [31:0]      dataInMem_hi_lo_151;
  assign dataInMem_hi_lo_151 = _GEN_430;
  wire [47:0]      dataInMem_hi_469 = {dataInMem_hi_hi_277, dataRegroupBySew_2_1_9};
  wire [31:0]      _GEN_431 = {dataRegroupBySew_4_1_10, dataRegroupBySew_3_1_10};
  wire [31:0]      dataInMem_hi_hi_278;
  assign dataInMem_hi_hi_278 = _GEN_431;
  wire [31:0]      dataInMem_hi_lo_152;
  assign dataInMem_hi_lo_152 = _GEN_431;
  wire [47:0]      dataInMem_hi_470 = {dataInMem_hi_hi_278, dataRegroupBySew_2_1_10};
  wire [31:0]      _GEN_432 = {dataRegroupBySew_4_1_11, dataRegroupBySew_3_1_11};
  wire [31:0]      dataInMem_hi_hi_279;
  assign dataInMem_hi_hi_279 = _GEN_432;
  wire [31:0]      dataInMem_hi_lo_153;
  assign dataInMem_hi_lo_153 = _GEN_432;
  wire [47:0]      dataInMem_hi_471 = {dataInMem_hi_hi_279, dataRegroupBySew_2_1_11};
  wire [31:0]      _GEN_433 = {dataRegroupBySew_4_1_12, dataRegroupBySew_3_1_12};
  wire [31:0]      dataInMem_hi_hi_280;
  assign dataInMem_hi_hi_280 = _GEN_433;
  wire [31:0]      dataInMem_hi_lo_154;
  assign dataInMem_hi_lo_154 = _GEN_433;
  wire [47:0]      dataInMem_hi_472 = {dataInMem_hi_hi_280, dataRegroupBySew_2_1_12};
  wire [31:0]      _GEN_434 = {dataRegroupBySew_4_1_13, dataRegroupBySew_3_1_13};
  wire [31:0]      dataInMem_hi_hi_281;
  assign dataInMem_hi_hi_281 = _GEN_434;
  wire [31:0]      dataInMem_hi_lo_155;
  assign dataInMem_hi_lo_155 = _GEN_434;
  wire [47:0]      dataInMem_hi_473 = {dataInMem_hi_hi_281, dataRegroupBySew_2_1_13};
  wire [31:0]      _GEN_435 = {dataRegroupBySew_4_1_14, dataRegroupBySew_3_1_14};
  wire [31:0]      dataInMem_hi_hi_282;
  assign dataInMem_hi_hi_282 = _GEN_435;
  wire [31:0]      dataInMem_hi_lo_156;
  assign dataInMem_hi_lo_156 = _GEN_435;
  wire [47:0]      dataInMem_hi_474 = {dataInMem_hi_hi_282, dataRegroupBySew_2_1_14};
  wire [31:0]      _GEN_436 = {dataRegroupBySew_4_1_15, dataRegroupBySew_3_1_15};
  wire [31:0]      dataInMem_hi_hi_283;
  assign dataInMem_hi_hi_283 = _GEN_436;
  wire [31:0]      dataInMem_hi_lo_157;
  assign dataInMem_hi_lo_157 = _GEN_436;
  wire [47:0]      dataInMem_hi_475 = {dataInMem_hi_hi_283, dataRegroupBySew_2_1_15};
  wire [31:0]      _GEN_437 = {dataRegroupBySew_4_1_16, dataRegroupBySew_3_1_16};
  wire [31:0]      dataInMem_hi_hi_284;
  assign dataInMem_hi_hi_284 = _GEN_437;
  wire [31:0]      dataInMem_hi_lo_158;
  assign dataInMem_hi_lo_158 = _GEN_437;
  wire [47:0]      dataInMem_hi_476 = {dataInMem_hi_hi_284, dataRegroupBySew_2_1_16};
  wire [31:0]      _GEN_438 = {dataRegroupBySew_4_1_17, dataRegroupBySew_3_1_17};
  wire [31:0]      dataInMem_hi_hi_285;
  assign dataInMem_hi_hi_285 = _GEN_438;
  wire [31:0]      dataInMem_hi_lo_159;
  assign dataInMem_hi_lo_159 = _GEN_438;
  wire [47:0]      dataInMem_hi_477 = {dataInMem_hi_hi_285, dataRegroupBySew_2_1_17};
  wire [31:0]      _GEN_439 = {dataRegroupBySew_4_1_18, dataRegroupBySew_3_1_18};
  wire [31:0]      dataInMem_hi_hi_286;
  assign dataInMem_hi_hi_286 = _GEN_439;
  wire [31:0]      dataInMem_hi_lo_160;
  assign dataInMem_hi_lo_160 = _GEN_439;
  wire [47:0]      dataInMem_hi_478 = {dataInMem_hi_hi_286, dataRegroupBySew_2_1_18};
  wire [31:0]      _GEN_440 = {dataRegroupBySew_4_1_19, dataRegroupBySew_3_1_19};
  wire [31:0]      dataInMem_hi_hi_287;
  assign dataInMem_hi_hi_287 = _GEN_440;
  wire [31:0]      dataInMem_hi_lo_161;
  assign dataInMem_hi_lo_161 = _GEN_440;
  wire [47:0]      dataInMem_hi_479 = {dataInMem_hi_hi_287, dataRegroupBySew_2_1_19};
  wire [31:0]      _GEN_441 = {dataRegroupBySew_4_1_20, dataRegroupBySew_3_1_20};
  wire [31:0]      dataInMem_hi_hi_288;
  assign dataInMem_hi_hi_288 = _GEN_441;
  wire [31:0]      dataInMem_hi_lo_162;
  assign dataInMem_hi_lo_162 = _GEN_441;
  wire [47:0]      dataInMem_hi_480 = {dataInMem_hi_hi_288, dataRegroupBySew_2_1_20};
  wire [31:0]      _GEN_442 = {dataRegroupBySew_4_1_21, dataRegroupBySew_3_1_21};
  wire [31:0]      dataInMem_hi_hi_289;
  assign dataInMem_hi_hi_289 = _GEN_442;
  wire [31:0]      dataInMem_hi_lo_163;
  assign dataInMem_hi_lo_163 = _GEN_442;
  wire [47:0]      dataInMem_hi_481 = {dataInMem_hi_hi_289, dataRegroupBySew_2_1_21};
  wire [31:0]      _GEN_443 = {dataRegroupBySew_4_1_22, dataRegroupBySew_3_1_22};
  wire [31:0]      dataInMem_hi_hi_290;
  assign dataInMem_hi_hi_290 = _GEN_443;
  wire [31:0]      dataInMem_hi_lo_164;
  assign dataInMem_hi_lo_164 = _GEN_443;
  wire [47:0]      dataInMem_hi_482 = {dataInMem_hi_hi_290, dataRegroupBySew_2_1_22};
  wire [31:0]      _GEN_444 = {dataRegroupBySew_4_1_23, dataRegroupBySew_3_1_23};
  wire [31:0]      dataInMem_hi_hi_291;
  assign dataInMem_hi_hi_291 = _GEN_444;
  wire [31:0]      dataInMem_hi_lo_165;
  assign dataInMem_hi_lo_165 = _GEN_444;
  wire [47:0]      dataInMem_hi_483 = {dataInMem_hi_hi_291, dataRegroupBySew_2_1_23};
  wire [31:0]      _GEN_445 = {dataRegroupBySew_4_1_24, dataRegroupBySew_3_1_24};
  wire [31:0]      dataInMem_hi_hi_292;
  assign dataInMem_hi_hi_292 = _GEN_445;
  wire [31:0]      dataInMem_hi_lo_166;
  assign dataInMem_hi_lo_166 = _GEN_445;
  wire [47:0]      dataInMem_hi_484 = {dataInMem_hi_hi_292, dataRegroupBySew_2_1_24};
  wire [31:0]      _GEN_446 = {dataRegroupBySew_4_1_25, dataRegroupBySew_3_1_25};
  wire [31:0]      dataInMem_hi_hi_293;
  assign dataInMem_hi_hi_293 = _GEN_446;
  wire [31:0]      dataInMem_hi_lo_167;
  assign dataInMem_hi_lo_167 = _GEN_446;
  wire [47:0]      dataInMem_hi_485 = {dataInMem_hi_hi_293, dataRegroupBySew_2_1_25};
  wire [31:0]      _GEN_447 = {dataRegroupBySew_4_1_26, dataRegroupBySew_3_1_26};
  wire [31:0]      dataInMem_hi_hi_294;
  assign dataInMem_hi_hi_294 = _GEN_447;
  wire [31:0]      dataInMem_hi_lo_168;
  assign dataInMem_hi_lo_168 = _GEN_447;
  wire [47:0]      dataInMem_hi_486 = {dataInMem_hi_hi_294, dataRegroupBySew_2_1_26};
  wire [31:0]      _GEN_448 = {dataRegroupBySew_4_1_27, dataRegroupBySew_3_1_27};
  wire [31:0]      dataInMem_hi_hi_295;
  assign dataInMem_hi_hi_295 = _GEN_448;
  wire [31:0]      dataInMem_hi_lo_169;
  assign dataInMem_hi_lo_169 = _GEN_448;
  wire [47:0]      dataInMem_hi_487 = {dataInMem_hi_hi_295, dataRegroupBySew_2_1_27};
  wire [31:0]      _GEN_449 = {dataRegroupBySew_4_1_28, dataRegroupBySew_3_1_28};
  wire [31:0]      dataInMem_hi_hi_296;
  assign dataInMem_hi_hi_296 = _GEN_449;
  wire [31:0]      dataInMem_hi_lo_170;
  assign dataInMem_hi_lo_170 = _GEN_449;
  wire [47:0]      dataInMem_hi_488 = {dataInMem_hi_hi_296, dataRegroupBySew_2_1_28};
  wire [31:0]      _GEN_450 = {dataRegroupBySew_4_1_29, dataRegroupBySew_3_1_29};
  wire [31:0]      dataInMem_hi_hi_297;
  assign dataInMem_hi_hi_297 = _GEN_450;
  wire [31:0]      dataInMem_hi_lo_171;
  assign dataInMem_hi_lo_171 = _GEN_450;
  wire [47:0]      dataInMem_hi_489 = {dataInMem_hi_hi_297, dataRegroupBySew_2_1_29};
  wire [31:0]      _GEN_451 = {dataRegroupBySew_4_1_30, dataRegroupBySew_3_1_30};
  wire [31:0]      dataInMem_hi_hi_298;
  assign dataInMem_hi_hi_298 = _GEN_451;
  wire [31:0]      dataInMem_hi_lo_172;
  assign dataInMem_hi_lo_172 = _GEN_451;
  wire [47:0]      dataInMem_hi_490 = {dataInMem_hi_hi_298, dataRegroupBySew_2_1_30};
  wire [31:0]      _GEN_452 = {dataRegroupBySew_4_1_31, dataRegroupBySew_3_1_31};
  wire [31:0]      dataInMem_hi_hi_299;
  assign dataInMem_hi_hi_299 = _GEN_452;
  wire [31:0]      dataInMem_hi_lo_173;
  assign dataInMem_hi_lo_173 = _GEN_452;
  wire [47:0]      dataInMem_hi_491 = {dataInMem_hi_hi_299, dataRegroupBySew_2_1_31};
  wire [159:0]     dataInMem_lo_lo_lo_lo_12 = {dataInMem_hi_461, dataInMem_lo_365, dataInMem_hi_460, dataInMem_lo_364};
  wire [159:0]     dataInMem_lo_lo_lo_hi_12 = {dataInMem_hi_463, dataInMem_lo_367, dataInMem_hi_462, dataInMem_lo_366};
  wire [319:0]     dataInMem_lo_lo_lo_12 = {dataInMem_lo_lo_lo_hi_12, dataInMem_lo_lo_lo_lo_12};
  wire [159:0]     dataInMem_lo_lo_hi_lo_12 = {dataInMem_hi_465, dataInMem_lo_369, dataInMem_hi_464, dataInMem_lo_368};
  wire [159:0]     dataInMem_lo_lo_hi_hi_12 = {dataInMem_hi_467, dataInMem_lo_371, dataInMem_hi_466, dataInMem_lo_370};
  wire [319:0]     dataInMem_lo_lo_hi_12 = {dataInMem_lo_lo_hi_hi_12, dataInMem_lo_lo_hi_lo_12};
  wire [639:0]     dataInMem_lo_lo_76 = {dataInMem_lo_lo_hi_12, dataInMem_lo_lo_lo_12};
  wire [159:0]     dataInMem_lo_hi_lo_lo_12 = {dataInMem_hi_469, dataInMem_lo_373, dataInMem_hi_468, dataInMem_lo_372};
  wire [159:0]     dataInMem_lo_hi_lo_hi_12 = {dataInMem_hi_471, dataInMem_lo_375, dataInMem_hi_470, dataInMem_lo_374};
  wire [319:0]     dataInMem_lo_hi_lo_12 = {dataInMem_lo_hi_lo_hi_12, dataInMem_lo_hi_lo_lo_12};
  wire [159:0]     dataInMem_lo_hi_hi_lo_12 = {dataInMem_hi_473, dataInMem_lo_377, dataInMem_hi_472, dataInMem_lo_376};
  wire [159:0]     dataInMem_lo_hi_hi_hi_12 = {dataInMem_hi_475, dataInMem_lo_379, dataInMem_hi_474, dataInMem_lo_378};
  wire [319:0]     dataInMem_lo_hi_hi_12 = {dataInMem_lo_hi_hi_hi_12, dataInMem_lo_hi_hi_lo_12};
  wire [639:0]     dataInMem_lo_hi_204 = {dataInMem_lo_hi_hi_12, dataInMem_lo_hi_lo_12};
  wire [1279:0]    dataInMem_lo_396 = {dataInMem_lo_hi_204, dataInMem_lo_lo_76};
  wire [159:0]     dataInMem_hi_lo_lo_lo_12 = {dataInMem_hi_477, dataInMem_lo_381, dataInMem_hi_476, dataInMem_lo_380};
  wire [159:0]     dataInMem_hi_lo_lo_hi_12 = {dataInMem_hi_479, dataInMem_lo_383, dataInMem_hi_478, dataInMem_lo_382};
  wire [319:0]     dataInMem_hi_lo_lo_12 = {dataInMem_hi_lo_lo_hi_12, dataInMem_hi_lo_lo_lo_12};
  wire [159:0]     dataInMem_hi_lo_hi_lo_12 = {dataInMem_hi_481, dataInMem_lo_385, dataInMem_hi_480, dataInMem_lo_384};
  wire [159:0]     dataInMem_hi_lo_hi_hi_12 = {dataInMem_hi_483, dataInMem_lo_387, dataInMem_hi_482, dataInMem_lo_386};
  wire [319:0]     dataInMem_hi_lo_hi_12 = {dataInMem_hi_lo_hi_hi_12, dataInMem_hi_lo_hi_lo_12};
  wire [639:0]     dataInMem_hi_lo_140 = {dataInMem_hi_lo_hi_12, dataInMem_hi_lo_lo_12};
  wire [159:0]     dataInMem_hi_hi_lo_lo_12 = {dataInMem_hi_485, dataInMem_lo_389, dataInMem_hi_484, dataInMem_lo_388};
  wire [159:0]     dataInMem_hi_hi_lo_hi_12 = {dataInMem_hi_487, dataInMem_lo_391, dataInMem_hi_486, dataInMem_lo_390};
  wire [319:0]     dataInMem_hi_hi_lo_12 = {dataInMem_hi_hi_lo_hi_12, dataInMem_hi_hi_lo_lo_12};
  wire [159:0]     dataInMem_hi_hi_hi_lo_12 = {dataInMem_hi_489, dataInMem_lo_393, dataInMem_hi_488, dataInMem_lo_392};
  wire [159:0]     dataInMem_hi_hi_hi_hi_12 = {dataInMem_hi_491, dataInMem_lo_395, dataInMem_hi_490, dataInMem_lo_394};
  wire [319:0]     dataInMem_hi_hi_hi_12 = {dataInMem_hi_hi_hi_hi_12, dataInMem_hi_hi_hi_lo_12};
  wire [639:0]     dataInMem_hi_hi_300 = {dataInMem_hi_hi_hi_12, dataInMem_hi_hi_lo_12};
  wire [1279:0]    dataInMem_hi_492 = {dataInMem_hi_hi_300, dataInMem_hi_lo_140};
  wire [2559:0]    dataInMem_12 = {dataInMem_hi_492, dataInMem_lo_396};
  wire [511:0]     regroupCacheLine_12_0 = dataInMem_12[511:0];
  wire [511:0]     regroupCacheLine_12_1 = dataInMem_12[1023:512];
  wire [511:0]     regroupCacheLine_12_2 = dataInMem_12[1535:1024];
  wire [511:0]     regroupCacheLine_12_3 = dataInMem_12[2047:1536];
  wire [511:0]     regroupCacheLine_12_4 = dataInMem_12[2559:2048];
  wire [511:0]     res_96 = regroupCacheLine_12_0;
  wire [511:0]     res_97 = regroupCacheLine_12_1;
  wire [511:0]     res_98 = regroupCacheLine_12_2;
  wire [511:0]     res_99 = regroupCacheLine_12_3;
  wire [511:0]     res_100 = regroupCacheLine_12_4;
  wire [1023:0]    lo_lo_12 = {res_97, res_96};
  wire [1023:0]    lo_hi_12 = {res_99, res_98};
  wire [2047:0]    lo_12 = {lo_hi_12, lo_lo_12};
  wire [1023:0]    hi_lo_12 = {512'h0, res_100};
  wire [2047:0]    hi_12 = {1024'h0, hi_lo_12};
  wire [4095:0]    regroupLoadData_1_4 = {hi_12, lo_12};
  wire [47:0]      dataInMem_lo_397 = {dataInMem_lo_hi_205, dataRegroupBySew_0_1_0};
  wire [31:0]      _GEN_453 = {dataRegroupBySew_5_1_0, dataRegroupBySew_4_1_0};
  wire [31:0]      dataInMem_hi_hi_301;
  assign dataInMem_hi_hi_301 = _GEN_453;
  wire [31:0]      dataInMem_hi_lo_175;
  assign dataInMem_hi_lo_175 = _GEN_453;
  wire [47:0]      dataInMem_hi_493 = {dataInMem_hi_hi_301, dataRegroupBySew_3_1_0};
  wire [47:0]      dataInMem_lo_398 = {dataInMem_lo_hi_206, dataRegroupBySew_0_1_1};
  wire [31:0]      _GEN_454 = {dataRegroupBySew_5_1_1, dataRegroupBySew_4_1_1};
  wire [31:0]      dataInMem_hi_hi_302;
  assign dataInMem_hi_hi_302 = _GEN_454;
  wire [31:0]      dataInMem_hi_lo_176;
  assign dataInMem_hi_lo_176 = _GEN_454;
  wire [47:0]      dataInMem_hi_494 = {dataInMem_hi_hi_302, dataRegroupBySew_3_1_1};
  wire [47:0]      dataInMem_lo_399 = {dataInMem_lo_hi_207, dataRegroupBySew_0_1_2};
  wire [31:0]      _GEN_455 = {dataRegroupBySew_5_1_2, dataRegroupBySew_4_1_2};
  wire [31:0]      dataInMem_hi_hi_303;
  assign dataInMem_hi_hi_303 = _GEN_455;
  wire [31:0]      dataInMem_hi_lo_177;
  assign dataInMem_hi_lo_177 = _GEN_455;
  wire [47:0]      dataInMem_hi_495 = {dataInMem_hi_hi_303, dataRegroupBySew_3_1_2};
  wire [47:0]      dataInMem_lo_400 = {dataInMem_lo_hi_208, dataRegroupBySew_0_1_3};
  wire [31:0]      _GEN_456 = {dataRegroupBySew_5_1_3, dataRegroupBySew_4_1_3};
  wire [31:0]      dataInMem_hi_hi_304;
  assign dataInMem_hi_hi_304 = _GEN_456;
  wire [31:0]      dataInMem_hi_lo_178;
  assign dataInMem_hi_lo_178 = _GEN_456;
  wire [47:0]      dataInMem_hi_496 = {dataInMem_hi_hi_304, dataRegroupBySew_3_1_3};
  wire [47:0]      dataInMem_lo_401 = {dataInMem_lo_hi_209, dataRegroupBySew_0_1_4};
  wire [31:0]      _GEN_457 = {dataRegroupBySew_5_1_4, dataRegroupBySew_4_1_4};
  wire [31:0]      dataInMem_hi_hi_305;
  assign dataInMem_hi_hi_305 = _GEN_457;
  wire [31:0]      dataInMem_hi_lo_179;
  assign dataInMem_hi_lo_179 = _GEN_457;
  wire [47:0]      dataInMem_hi_497 = {dataInMem_hi_hi_305, dataRegroupBySew_3_1_4};
  wire [47:0]      dataInMem_lo_402 = {dataInMem_lo_hi_210, dataRegroupBySew_0_1_5};
  wire [31:0]      _GEN_458 = {dataRegroupBySew_5_1_5, dataRegroupBySew_4_1_5};
  wire [31:0]      dataInMem_hi_hi_306;
  assign dataInMem_hi_hi_306 = _GEN_458;
  wire [31:0]      dataInMem_hi_lo_180;
  assign dataInMem_hi_lo_180 = _GEN_458;
  wire [47:0]      dataInMem_hi_498 = {dataInMem_hi_hi_306, dataRegroupBySew_3_1_5};
  wire [47:0]      dataInMem_lo_403 = {dataInMem_lo_hi_211, dataRegroupBySew_0_1_6};
  wire [31:0]      _GEN_459 = {dataRegroupBySew_5_1_6, dataRegroupBySew_4_1_6};
  wire [31:0]      dataInMem_hi_hi_307;
  assign dataInMem_hi_hi_307 = _GEN_459;
  wire [31:0]      dataInMem_hi_lo_181;
  assign dataInMem_hi_lo_181 = _GEN_459;
  wire [47:0]      dataInMem_hi_499 = {dataInMem_hi_hi_307, dataRegroupBySew_3_1_6};
  wire [47:0]      dataInMem_lo_404 = {dataInMem_lo_hi_212, dataRegroupBySew_0_1_7};
  wire [31:0]      _GEN_460 = {dataRegroupBySew_5_1_7, dataRegroupBySew_4_1_7};
  wire [31:0]      dataInMem_hi_hi_308;
  assign dataInMem_hi_hi_308 = _GEN_460;
  wire [31:0]      dataInMem_hi_lo_182;
  assign dataInMem_hi_lo_182 = _GEN_460;
  wire [47:0]      dataInMem_hi_500 = {dataInMem_hi_hi_308, dataRegroupBySew_3_1_7};
  wire [47:0]      dataInMem_lo_405 = {dataInMem_lo_hi_213, dataRegroupBySew_0_1_8};
  wire [31:0]      _GEN_461 = {dataRegroupBySew_5_1_8, dataRegroupBySew_4_1_8};
  wire [31:0]      dataInMem_hi_hi_309;
  assign dataInMem_hi_hi_309 = _GEN_461;
  wire [31:0]      dataInMem_hi_lo_183;
  assign dataInMem_hi_lo_183 = _GEN_461;
  wire [47:0]      dataInMem_hi_501 = {dataInMem_hi_hi_309, dataRegroupBySew_3_1_8};
  wire [47:0]      dataInMem_lo_406 = {dataInMem_lo_hi_214, dataRegroupBySew_0_1_9};
  wire [31:0]      _GEN_462 = {dataRegroupBySew_5_1_9, dataRegroupBySew_4_1_9};
  wire [31:0]      dataInMem_hi_hi_310;
  assign dataInMem_hi_hi_310 = _GEN_462;
  wire [31:0]      dataInMem_hi_lo_184;
  assign dataInMem_hi_lo_184 = _GEN_462;
  wire [47:0]      dataInMem_hi_502 = {dataInMem_hi_hi_310, dataRegroupBySew_3_1_9};
  wire [47:0]      dataInMem_lo_407 = {dataInMem_lo_hi_215, dataRegroupBySew_0_1_10};
  wire [31:0]      _GEN_463 = {dataRegroupBySew_5_1_10, dataRegroupBySew_4_1_10};
  wire [31:0]      dataInMem_hi_hi_311;
  assign dataInMem_hi_hi_311 = _GEN_463;
  wire [31:0]      dataInMem_hi_lo_185;
  assign dataInMem_hi_lo_185 = _GEN_463;
  wire [47:0]      dataInMem_hi_503 = {dataInMem_hi_hi_311, dataRegroupBySew_3_1_10};
  wire [47:0]      dataInMem_lo_408 = {dataInMem_lo_hi_216, dataRegroupBySew_0_1_11};
  wire [31:0]      _GEN_464 = {dataRegroupBySew_5_1_11, dataRegroupBySew_4_1_11};
  wire [31:0]      dataInMem_hi_hi_312;
  assign dataInMem_hi_hi_312 = _GEN_464;
  wire [31:0]      dataInMem_hi_lo_186;
  assign dataInMem_hi_lo_186 = _GEN_464;
  wire [47:0]      dataInMem_hi_504 = {dataInMem_hi_hi_312, dataRegroupBySew_3_1_11};
  wire [47:0]      dataInMem_lo_409 = {dataInMem_lo_hi_217, dataRegroupBySew_0_1_12};
  wire [31:0]      _GEN_465 = {dataRegroupBySew_5_1_12, dataRegroupBySew_4_1_12};
  wire [31:0]      dataInMem_hi_hi_313;
  assign dataInMem_hi_hi_313 = _GEN_465;
  wire [31:0]      dataInMem_hi_lo_187;
  assign dataInMem_hi_lo_187 = _GEN_465;
  wire [47:0]      dataInMem_hi_505 = {dataInMem_hi_hi_313, dataRegroupBySew_3_1_12};
  wire [47:0]      dataInMem_lo_410 = {dataInMem_lo_hi_218, dataRegroupBySew_0_1_13};
  wire [31:0]      _GEN_466 = {dataRegroupBySew_5_1_13, dataRegroupBySew_4_1_13};
  wire [31:0]      dataInMem_hi_hi_314;
  assign dataInMem_hi_hi_314 = _GEN_466;
  wire [31:0]      dataInMem_hi_lo_188;
  assign dataInMem_hi_lo_188 = _GEN_466;
  wire [47:0]      dataInMem_hi_506 = {dataInMem_hi_hi_314, dataRegroupBySew_3_1_13};
  wire [47:0]      dataInMem_lo_411 = {dataInMem_lo_hi_219, dataRegroupBySew_0_1_14};
  wire [31:0]      _GEN_467 = {dataRegroupBySew_5_1_14, dataRegroupBySew_4_1_14};
  wire [31:0]      dataInMem_hi_hi_315;
  assign dataInMem_hi_hi_315 = _GEN_467;
  wire [31:0]      dataInMem_hi_lo_189;
  assign dataInMem_hi_lo_189 = _GEN_467;
  wire [47:0]      dataInMem_hi_507 = {dataInMem_hi_hi_315, dataRegroupBySew_3_1_14};
  wire [47:0]      dataInMem_lo_412 = {dataInMem_lo_hi_220, dataRegroupBySew_0_1_15};
  wire [31:0]      _GEN_468 = {dataRegroupBySew_5_1_15, dataRegroupBySew_4_1_15};
  wire [31:0]      dataInMem_hi_hi_316;
  assign dataInMem_hi_hi_316 = _GEN_468;
  wire [31:0]      dataInMem_hi_lo_190;
  assign dataInMem_hi_lo_190 = _GEN_468;
  wire [47:0]      dataInMem_hi_508 = {dataInMem_hi_hi_316, dataRegroupBySew_3_1_15};
  wire [47:0]      dataInMem_lo_413 = {dataInMem_lo_hi_221, dataRegroupBySew_0_1_16};
  wire [31:0]      _GEN_469 = {dataRegroupBySew_5_1_16, dataRegroupBySew_4_1_16};
  wire [31:0]      dataInMem_hi_hi_317;
  assign dataInMem_hi_hi_317 = _GEN_469;
  wire [31:0]      dataInMem_hi_lo_191;
  assign dataInMem_hi_lo_191 = _GEN_469;
  wire [47:0]      dataInMem_hi_509 = {dataInMem_hi_hi_317, dataRegroupBySew_3_1_16};
  wire [47:0]      dataInMem_lo_414 = {dataInMem_lo_hi_222, dataRegroupBySew_0_1_17};
  wire [31:0]      _GEN_470 = {dataRegroupBySew_5_1_17, dataRegroupBySew_4_1_17};
  wire [31:0]      dataInMem_hi_hi_318;
  assign dataInMem_hi_hi_318 = _GEN_470;
  wire [31:0]      dataInMem_hi_lo_192;
  assign dataInMem_hi_lo_192 = _GEN_470;
  wire [47:0]      dataInMem_hi_510 = {dataInMem_hi_hi_318, dataRegroupBySew_3_1_17};
  wire [47:0]      dataInMem_lo_415 = {dataInMem_lo_hi_223, dataRegroupBySew_0_1_18};
  wire [31:0]      _GEN_471 = {dataRegroupBySew_5_1_18, dataRegroupBySew_4_1_18};
  wire [31:0]      dataInMem_hi_hi_319;
  assign dataInMem_hi_hi_319 = _GEN_471;
  wire [31:0]      dataInMem_hi_lo_193;
  assign dataInMem_hi_lo_193 = _GEN_471;
  wire [47:0]      dataInMem_hi_511 = {dataInMem_hi_hi_319, dataRegroupBySew_3_1_18};
  wire [47:0]      dataInMem_lo_416 = {dataInMem_lo_hi_224, dataRegroupBySew_0_1_19};
  wire [31:0]      _GEN_472 = {dataRegroupBySew_5_1_19, dataRegroupBySew_4_1_19};
  wire [31:0]      dataInMem_hi_hi_320;
  assign dataInMem_hi_hi_320 = _GEN_472;
  wire [31:0]      dataInMem_hi_lo_194;
  assign dataInMem_hi_lo_194 = _GEN_472;
  wire [47:0]      dataInMem_hi_512 = {dataInMem_hi_hi_320, dataRegroupBySew_3_1_19};
  wire [47:0]      dataInMem_lo_417 = {dataInMem_lo_hi_225, dataRegroupBySew_0_1_20};
  wire [31:0]      _GEN_473 = {dataRegroupBySew_5_1_20, dataRegroupBySew_4_1_20};
  wire [31:0]      dataInMem_hi_hi_321;
  assign dataInMem_hi_hi_321 = _GEN_473;
  wire [31:0]      dataInMem_hi_lo_195;
  assign dataInMem_hi_lo_195 = _GEN_473;
  wire [47:0]      dataInMem_hi_513 = {dataInMem_hi_hi_321, dataRegroupBySew_3_1_20};
  wire [47:0]      dataInMem_lo_418 = {dataInMem_lo_hi_226, dataRegroupBySew_0_1_21};
  wire [31:0]      _GEN_474 = {dataRegroupBySew_5_1_21, dataRegroupBySew_4_1_21};
  wire [31:0]      dataInMem_hi_hi_322;
  assign dataInMem_hi_hi_322 = _GEN_474;
  wire [31:0]      dataInMem_hi_lo_196;
  assign dataInMem_hi_lo_196 = _GEN_474;
  wire [47:0]      dataInMem_hi_514 = {dataInMem_hi_hi_322, dataRegroupBySew_3_1_21};
  wire [47:0]      dataInMem_lo_419 = {dataInMem_lo_hi_227, dataRegroupBySew_0_1_22};
  wire [31:0]      _GEN_475 = {dataRegroupBySew_5_1_22, dataRegroupBySew_4_1_22};
  wire [31:0]      dataInMem_hi_hi_323;
  assign dataInMem_hi_hi_323 = _GEN_475;
  wire [31:0]      dataInMem_hi_lo_197;
  assign dataInMem_hi_lo_197 = _GEN_475;
  wire [47:0]      dataInMem_hi_515 = {dataInMem_hi_hi_323, dataRegroupBySew_3_1_22};
  wire [47:0]      dataInMem_lo_420 = {dataInMem_lo_hi_228, dataRegroupBySew_0_1_23};
  wire [31:0]      _GEN_476 = {dataRegroupBySew_5_1_23, dataRegroupBySew_4_1_23};
  wire [31:0]      dataInMem_hi_hi_324;
  assign dataInMem_hi_hi_324 = _GEN_476;
  wire [31:0]      dataInMem_hi_lo_198;
  assign dataInMem_hi_lo_198 = _GEN_476;
  wire [47:0]      dataInMem_hi_516 = {dataInMem_hi_hi_324, dataRegroupBySew_3_1_23};
  wire [47:0]      dataInMem_lo_421 = {dataInMem_lo_hi_229, dataRegroupBySew_0_1_24};
  wire [31:0]      _GEN_477 = {dataRegroupBySew_5_1_24, dataRegroupBySew_4_1_24};
  wire [31:0]      dataInMem_hi_hi_325;
  assign dataInMem_hi_hi_325 = _GEN_477;
  wire [31:0]      dataInMem_hi_lo_199;
  assign dataInMem_hi_lo_199 = _GEN_477;
  wire [47:0]      dataInMem_hi_517 = {dataInMem_hi_hi_325, dataRegroupBySew_3_1_24};
  wire [47:0]      dataInMem_lo_422 = {dataInMem_lo_hi_230, dataRegroupBySew_0_1_25};
  wire [31:0]      _GEN_478 = {dataRegroupBySew_5_1_25, dataRegroupBySew_4_1_25};
  wire [31:0]      dataInMem_hi_hi_326;
  assign dataInMem_hi_hi_326 = _GEN_478;
  wire [31:0]      dataInMem_hi_lo_200;
  assign dataInMem_hi_lo_200 = _GEN_478;
  wire [47:0]      dataInMem_hi_518 = {dataInMem_hi_hi_326, dataRegroupBySew_3_1_25};
  wire [47:0]      dataInMem_lo_423 = {dataInMem_lo_hi_231, dataRegroupBySew_0_1_26};
  wire [31:0]      _GEN_479 = {dataRegroupBySew_5_1_26, dataRegroupBySew_4_1_26};
  wire [31:0]      dataInMem_hi_hi_327;
  assign dataInMem_hi_hi_327 = _GEN_479;
  wire [31:0]      dataInMem_hi_lo_201;
  assign dataInMem_hi_lo_201 = _GEN_479;
  wire [47:0]      dataInMem_hi_519 = {dataInMem_hi_hi_327, dataRegroupBySew_3_1_26};
  wire [47:0]      dataInMem_lo_424 = {dataInMem_lo_hi_232, dataRegroupBySew_0_1_27};
  wire [31:0]      _GEN_480 = {dataRegroupBySew_5_1_27, dataRegroupBySew_4_1_27};
  wire [31:0]      dataInMem_hi_hi_328;
  assign dataInMem_hi_hi_328 = _GEN_480;
  wire [31:0]      dataInMem_hi_lo_202;
  assign dataInMem_hi_lo_202 = _GEN_480;
  wire [47:0]      dataInMem_hi_520 = {dataInMem_hi_hi_328, dataRegroupBySew_3_1_27};
  wire [47:0]      dataInMem_lo_425 = {dataInMem_lo_hi_233, dataRegroupBySew_0_1_28};
  wire [31:0]      _GEN_481 = {dataRegroupBySew_5_1_28, dataRegroupBySew_4_1_28};
  wire [31:0]      dataInMem_hi_hi_329;
  assign dataInMem_hi_hi_329 = _GEN_481;
  wire [31:0]      dataInMem_hi_lo_203;
  assign dataInMem_hi_lo_203 = _GEN_481;
  wire [47:0]      dataInMem_hi_521 = {dataInMem_hi_hi_329, dataRegroupBySew_3_1_28};
  wire [47:0]      dataInMem_lo_426 = {dataInMem_lo_hi_234, dataRegroupBySew_0_1_29};
  wire [31:0]      _GEN_482 = {dataRegroupBySew_5_1_29, dataRegroupBySew_4_1_29};
  wire [31:0]      dataInMem_hi_hi_330;
  assign dataInMem_hi_hi_330 = _GEN_482;
  wire [31:0]      dataInMem_hi_lo_204;
  assign dataInMem_hi_lo_204 = _GEN_482;
  wire [47:0]      dataInMem_hi_522 = {dataInMem_hi_hi_330, dataRegroupBySew_3_1_29};
  wire [47:0]      dataInMem_lo_427 = {dataInMem_lo_hi_235, dataRegroupBySew_0_1_30};
  wire [31:0]      _GEN_483 = {dataRegroupBySew_5_1_30, dataRegroupBySew_4_1_30};
  wire [31:0]      dataInMem_hi_hi_331;
  assign dataInMem_hi_hi_331 = _GEN_483;
  wire [31:0]      dataInMem_hi_lo_205;
  assign dataInMem_hi_lo_205 = _GEN_483;
  wire [47:0]      dataInMem_hi_523 = {dataInMem_hi_hi_331, dataRegroupBySew_3_1_30};
  wire [47:0]      dataInMem_lo_428 = {dataInMem_lo_hi_236, dataRegroupBySew_0_1_31};
  wire [31:0]      _GEN_484 = {dataRegroupBySew_5_1_31, dataRegroupBySew_4_1_31};
  wire [31:0]      dataInMem_hi_hi_332;
  assign dataInMem_hi_hi_332 = _GEN_484;
  wire [31:0]      dataInMem_hi_lo_206;
  assign dataInMem_hi_lo_206 = _GEN_484;
  wire [47:0]      dataInMem_hi_524 = {dataInMem_hi_hi_332, dataRegroupBySew_3_1_31};
  wire [191:0]     dataInMem_lo_lo_lo_lo_13 = {dataInMem_hi_494, dataInMem_lo_398, dataInMem_hi_493, dataInMem_lo_397};
  wire [191:0]     dataInMem_lo_lo_lo_hi_13 = {dataInMem_hi_496, dataInMem_lo_400, dataInMem_hi_495, dataInMem_lo_399};
  wire [383:0]     dataInMem_lo_lo_lo_13 = {dataInMem_lo_lo_lo_hi_13, dataInMem_lo_lo_lo_lo_13};
  wire [191:0]     dataInMem_lo_lo_hi_lo_13 = {dataInMem_hi_498, dataInMem_lo_402, dataInMem_hi_497, dataInMem_lo_401};
  wire [191:0]     dataInMem_lo_lo_hi_hi_13 = {dataInMem_hi_500, dataInMem_lo_404, dataInMem_hi_499, dataInMem_lo_403};
  wire [383:0]     dataInMem_lo_lo_hi_13 = {dataInMem_lo_lo_hi_hi_13, dataInMem_lo_lo_hi_lo_13};
  wire [767:0]     dataInMem_lo_lo_77 = {dataInMem_lo_lo_hi_13, dataInMem_lo_lo_lo_13};
  wire [191:0]     dataInMem_lo_hi_lo_lo_13 = {dataInMem_hi_502, dataInMem_lo_406, dataInMem_hi_501, dataInMem_lo_405};
  wire [191:0]     dataInMem_lo_hi_lo_hi_13 = {dataInMem_hi_504, dataInMem_lo_408, dataInMem_hi_503, dataInMem_lo_407};
  wire [383:0]     dataInMem_lo_hi_lo_13 = {dataInMem_lo_hi_lo_hi_13, dataInMem_lo_hi_lo_lo_13};
  wire [191:0]     dataInMem_lo_hi_hi_lo_13 = {dataInMem_hi_506, dataInMem_lo_410, dataInMem_hi_505, dataInMem_lo_409};
  wire [191:0]     dataInMem_lo_hi_hi_hi_13 = {dataInMem_hi_508, dataInMem_lo_412, dataInMem_hi_507, dataInMem_lo_411};
  wire [383:0]     dataInMem_lo_hi_hi_13 = {dataInMem_lo_hi_hi_hi_13, dataInMem_lo_hi_hi_lo_13};
  wire [767:0]     dataInMem_lo_hi_237 = {dataInMem_lo_hi_hi_13, dataInMem_lo_hi_lo_13};
  wire [1535:0]    dataInMem_lo_429 = {dataInMem_lo_hi_237, dataInMem_lo_lo_77};
  wire [191:0]     dataInMem_hi_lo_lo_lo_13 = {dataInMem_hi_510, dataInMem_lo_414, dataInMem_hi_509, dataInMem_lo_413};
  wire [191:0]     dataInMem_hi_lo_lo_hi_13 = {dataInMem_hi_512, dataInMem_lo_416, dataInMem_hi_511, dataInMem_lo_415};
  wire [383:0]     dataInMem_hi_lo_lo_13 = {dataInMem_hi_lo_lo_hi_13, dataInMem_hi_lo_lo_lo_13};
  wire [191:0]     dataInMem_hi_lo_hi_lo_13 = {dataInMem_hi_514, dataInMem_lo_418, dataInMem_hi_513, dataInMem_lo_417};
  wire [191:0]     dataInMem_hi_lo_hi_hi_13 = {dataInMem_hi_516, dataInMem_lo_420, dataInMem_hi_515, dataInMem_lo_419};
  wire [383:0]     dataInMem_hi_lo_hi_13 = {dataInMem_hi_lo_hi_hi_13, dataInMem_hi_lo_hi_lo_13};
  wire [767:0]     dataInMem_hi_lo_141 = {dataInMem_hi_lo_hi_13, dataInMem_hi_lo_lo_13};
  wire [191:0]     dataInMem_hi_hi_lo_lo_13 = {dataInMem_hi_518, dataInMem_lo_422, dataInMem_hi_517, dataInMem_lo_421};
  wire [191:0]     dataInMem_hi_hi_lo_hi_13 = {dataInMem_hi_520, dataInMem_lo_424, dataInMem_hi_519, dataInMem_lo_423};
  wire [383:0]     dataInMem_hi_hi_lo_13 = {dataInMem_hi_hi_lo_hi_13, dataInMem_hi_hi_lo_lo_13};
  wire [191:0]     dataInMem_hi_hi_hi_lo_13 = {dataInMem_hi_522, dataInMem_lo_426, dataInMem_hi_521, dataInMem_lo_425};
  wire [191:0]     dataInMem_hi_hi_hi_hi_13 = {dataInMem_hi_524, dataInMem_lo_428, dataInMem_hi_523, dataInMem_lo_427};
  wire [383:0]     dataInMem_hi_hi_hi_13 = {dataInMem_hi_hi_hi_hi_13, dataInMem_hi_hi_hi_lo_13};
  wire [767:0]     dataInMem_hi_hi_333 = {dataInMem_hi_hi_hi_13, dataInMem_hi_hi_lo_13};
  wire [1535:0]    dataInMem_hi_525 = {dataInMem_hi_hi_333, dataInMem_hi_lo_141};
  wire [3071:0]    dataInMem_13 = {dataInMem_hi_525, dataInMem_lo_429};
  wire [511:0]     regroupCacheLine_13_0 = dataInMem_13[511:0];
  wire [511:0]     regroupCacheLine_13_1 = dataInMem_13[1023:512];
  wire [511:0]     regroupCacheLine_13_2 = dataInMem_13[1535:1024];
  wire [511:0]     regroupCacheLine_13_3 = dataInMem_13[2047:1536];
  wire [511:0]     regroupCacheLine_13_4 = dataInMem_13[2559:2048];
  wire [511:0]     regroupCacheLine_13_5 = dataInMem_13[3071:2560];
  wire [511:0]     res_104 = regroupCacheLine_13_0;
  wire [511:0]     res_105 = regroupCacheLine_13_1;
  wire [511:0]     res_106 = regroupCacheLine_13_2;
  wire [511:0]     res_107 = regroupCacheLine_13_3;
  wire [511:0]     res_108 = regroupCacheLine_13_4;
  wire [511:0]     res_109 = regroupCacheLine_13_5;
  wire [1023:0]    lo_lo_13 = {res_105, res_104};
  wire [1023:0]    lo_hi_13 = {res_107, res_106};
  wire [2047:0]    lo_13 = {lo_hi_13, lo_lo_13};
  wire [1023:0]    hi_lo_13 = {res_109, res_108};
  wire [2047:0]    hi_13 = {1024'h0, hi_lo_13};
  wire [4095:0]    regroupLoadData_1_5 = {hi_13, lo_13};
  wire [47:0]      dataInMem_lo_430 = {dataInMem_lo_hi_238, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_hi_hi_334 = {dataRegroupBySew_6_1_0, dataRegroupBySew_5_1_0};
  wire [63:0]      dataInMem_hi_526 = {dataInMem_hi_hi_334, dataInMem_hi_lo_142};
  wire [47:0]      dataInMem_lo_431 = {dataInMem_lo_hi_239, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_hi_hi_335 = {dataRegroupBySew_6_1_1, dataRegroupBySew_5_1_1};
  wire [63:0]      dataInMem_hi_527 = {dataInMem_hi_hi_335, dataInMem_hi_lo_143};
  wire [47:0]      dataInMem_lo_432 = {dataInMem_lo_hi_240, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_hi_hi_336 = {dataRegroupBySew_6_1_2, dataRegroupBySew_5_1_2};
  wire [63:0]      dataInMem_hi_528 = {dataInMem_hi_hi_336, dataInMem_hi_lo_144};
  wire [47:0]      dataInMem_lo_433 = {dataInMem_lo_hi_241, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_hi_hi_337 = {dataRegroupBySew_6_1_3, dataRegroupBySew_5_1_3};
  wire [63:0]      dataInMem_hi_529 = {dataInMem_hi_hi_337, dataInMem_hi_lo_145};
  wire [47:0]      dataInMem_lo_434 = {dataInMem_lo_hi_242, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_hi_hi_338 = {dataRegroupBySew_6_1_4, dataRegroupBySew_5_1_4};
  wire [63:0]      dataInMem_hi_530 = {dataInMem_hi_hi_338, dataInMem_hi_lo_146};
  wire [47:0]      dataInMem_lo_435 = {dataInMem_lo_hi_243, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_hi_hi_339 = {dataRegroupBySew_6_1_5, dataRegroupBySew_5_1_5};
  wire [63:0]      dataInMem_hi_531 = {dataInMem_hi_hi_339, dataInMem_hi_lo_147};
  wire [47:0]      dataInMem_lo_436 = {dataInMem_lo_hi_244, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_hi_hi_340 = {dataRegroupBySew_6_1_6, dataRegroupBySew_5_1_6};
  wire [63:0]      dataInMem_hi_532 = {dataInMem_hi_hi_340, dataInMem_hi_lo_148};
  wire [47:0]      dataInMem_lo_437 = {dataInMem_lo_hi_245, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_hi_hi_341 = {dataRegroupBySew_6_1_7, dataRegroupBySew_5_1_7};
  wire [63:0]      dataInMem_hi_533 = {dataInMem_hi_hi_341, dataInMem_hi_lo_149};
  wire [47:0]      dataInMem_lo_438 = {dataInMem_lo_hi_246, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_hi_hi_342 = {dataRegroupBySew_6_1_8, dataRegroupBySew_5_1_8};
  wire [63:0]      dataInMem_hi_534 = {dataInMem_hi_hi_342, dataInMem_hi_lo_150};
  wire [47:0]      dataInMem_lo_439 = {dataInMem_lo_hi_247, dataRegroupBySew_0_1_9};
  wire [31:0]      dataInMem_hi_hi_343 = {dataRegroupBySew_6_1_9, dataRegroupBySew_5_1_9};
  wire [63:0]      dataInMem_hi_535 = {dataInMem_hi_hi_343, dataInMem_hi_lo_151};
  wire [47:0]      dataInMem_lo_440 = {dataInMem_lo_hi_248, dataRegroupBySew_0_1_10};
  wire [31:0]      dataInMem_hi_hi_344 = {dataRegroupBySew_6_1_10, dataRegroupBySew_5_1_10};
  wire [63:0]      dataInMem_hi_536 = {dataInMem_hi_hi_344, dataInMem_hi_lo_152};
  wire [47:0]      dataInMem_lo_441 = {dataInMem_lo_hi_249, dataRegroupBySew_0_1_11};
  wire [31:0]      dataInMem_hi_hi_345 = {dataRegroupBySew_6_1_11, dataRegroupBySew_5_1_11};
  wire [63:0]      dataInMem_hi_537 = {dataInMem_hi_hi_345, dataInMem_hi_lo_153};
  wire [47:0]      dataInMem_lo_442 = {dataInMem_lo_hi_250, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_hi_hi_346 = {dataRegroupBySew_6_1_12, dataRegroupBySew_5_1_12};
  wire [63:0]      dataInMem_hi_538 = {dataInMem_hi_hi_346, dataInMem_hi_lo_154};
  wire [47:0]      dataInMem_lo_443 = {dataInMem_lo_hi_251, dataRegroupBySew_0_1_13};
  wire [31:0]      dataInMem_hi_hi_347 = {dataRegroupBySew_6_1_13, dataRegroupBySew_5_1_13};
  wire [63:0]      dataInMem_hi_539 = {dataInMem_hi_hi_347, dataInMem_hi_lo_155};
  wire [47:0]      dataInMem_lo_444 = {dataInMem_lo_hi_252, dataRegroupBySew_0_1_14};
  wire [31:0]      dataInMem_hi_hi_348 = {dataRegroupBySew_6_1_14, dataRegroupBySew_5_1_14};
  wire [63:0]      dataInMem_hi_540 = {dataInMem_hi_hi_348, dataInMem_hi_lo_156};
  wire [47:0]      dataInMem_lo_445 = {dataInMem_lo_hi_253, dataRegroupBySew_0_1_15};
  wire [31:0]      dataInMem_hi_hi_349 = {dataRegroupBySew_6_1_15, dataRegroupBySew_5_1_15};
  wire [63:0]      dataInMem_hi_541 = {dataInMem_hi_hi_349, dataInMem_hi_lo_157};
  wire [47:0]      dataInMem_lo_446 = {dataInMem_lo_hi_254, dataRegroupBySew_0_1_16};
  wire [31:0]      dataInMem_hi_hi_350 = {dataRegroupBySew_6_1_16, dataRegroupBySew_5_1_16};
  wire [63:0]      dataInMem_hi_542 = {dataInMem_hi_hi_350, dataInMem_hi_lo_158};
  wire [47:0]      dataInMem_lo_447 = {dataInMem_lo_hi_255, dataRegroupBySew_0_1_17};
  wire [31:0]      dataInMem_hi_hi_351 = {dataRegroupBySew_6_1_17, dataRegroupBySew_5_1_17};
  wire [63:0]      dataInMem_hi_543 = {dataInMem_hi_hi_351, dataInMem_hi_lo_159};
  wire [47:0]      dataInMem_lo_448 = {dataInMem_lo_hi_256, dataRegroupBySew_0_1_18};
  wire [31:0]      dataInMem_hi_hi_352 = {dataRegroupBySew_6_1_18, dataRegroupBySew_5_1_18};
  wire [63:0]      dataInMem_hi_544 = {dataInMem_hi_hi_352, dataInMem_hi_lo_160};
  wire [47:0]      dataInMem_lo_449 = {dataInMem_lo_hi_257, dataRegroupBySew_0_1_19};
  wire [31:0]      dataInMem_hi_hi_353 = {dataRegroupBySew_6_1_19, dataRegroupBySew_5_1_19};
  wire [63:0]      dataInMem_hi_545 = {dataInMem_hi_hi_353, dataInMem_hi_lo_161};
  wire [47:0]      dataInMem_lo_450 = {dataInMem_lo_hi_258, dataRegroupBySew_0_1_20};
  wire [31:0]      dataInMem_hi_hi_354 = {dataRegroupBySew_6_1_20, dataRegroupBySew_5_1_20};
  wire [63:0]      dataInMem_hi_546 = {dataInMem_hi_hi_354, dataInMem_hi_lo_162};
  wire [47:0]      dataInMem_lo_451 = {dataInMem_lo_hi_259, dataRegroupBySew_0_1_21};
  wire [31:0]      dataInMem_hi_hi_355 = {dataRegroupBySew_6_1_21, dataRegroupBySew_5_1_21};
  wire [63:0]      dataInMem_hi_547 = {dataInMem_hi_hi_355, dataInMem_hi_lo_163};
  wire [47:0]      dataInMem_lo_452 = {dataInMem_lo_hi_260, dataRegroupBySew_0_1_22};
  wire [31:0]      dataInMem_hi_hi_356 = {dataRegroupBySew_6_1_22, dataRegroupBySew_5_1_22};
  wire [63:0]      dataInMem_hi_548 = {dataInMem_hi_hi_356, dataInMem_hi_lo_164};
  wire [47:0]      dataInMem_lo_453 = {dataInMem_lo_hi_261, dataRegroupBySew_0_1_23};
  wire [31:0]      dataInMem_hi_hi_357 = {dataRegroupBySew_6_1_23, dataRegroupBySew_5_1_23};
  wire [63:0]      dataInMem_hi_549 = {dataInMem_hi_hi_357, dataInMem_hi_lo_165};
  wire [47:0]      dataInMem_lo_454 = {dataInMem_lo_hi_262, dataRegroupBySew_0_1_24};
  wire [31:0]      dataInMem_hi_hi_358 = {dataRegroupBySew_6_1_24, dataRegroupBySew_5_1_24};
  wire [63:0]      dataInMem_hi_550 = {dataInMem_hi_hi_358, dataInMem_hi_lo_166};
  wire [47:0]      dataInMem_lo_455 = {dataInMem_lo_hi_263, dataRegroupBySew_0_1_25};
  wire [31:0]      dataInMem_hi_hi_359 = {dataRegroupBySew_6_1_25, dataRegroupBySew_5_1_25};
  wire [63:0]      dataInMem_hi_551 = {dataInMem_hi_hi_359, dataInMem_hi_lo_167};
  wire [47:0]      dataInMem_lo_456 = {dataInMem_lo_hi_264, dataRegroupBySew_0_1_26};
  wire [31:0]      dataInMem_hi_hi_360 = {dataRegroupBySew_6_1_26, dataRegroupBySew_5_1_26};
  wire [63:0]      dataInMem_hi_552 = {dataInMem_hi_hi_360, dataInMem_hi_lo_168};
  wire [47:0]      dataInMem_lo_457 = {dataInMem_lo_hi_265, dataRegroupBySew_0_1_27};
  wire [31:0]      dataInMem_hi_hi_361 = {dataRegroupBySew_6_1_27, dataRegroupBySew_5_1_27};
  wire [63:0]      dataInMem_hi_553 = {dataInMem_hi_hi_361, dataInMem_hi_lo_169};
  wire [47:0]      dataInMem_lo_458 = {dataInMem_lo_hi_266, dataRegroupBySew_0_1_28};
  wire [31:0]      dataInMem_hi_hi_362 = {dataRegroupBySew_6_1_28, dataRegroupBySew_5_1_28};
  wire [63:0]      dataInMem_hi_554 = {dataInMem_hi_hi_362, dataInMem_hi_lo_170};
  wire [47:0]      dataInMem_lo_459 = {dataInMem_lo_hi_267, dataRegroupBySew_0_1_29};
  wire [31:0]      dataInMem_hi_hi_363 = {dataRegroupBySew_6_1_29, dataRegroupBySew_5_1_29};
  wire [63:0]      dataInMem_hi_555 = {dataInMem_hi_hi_363, dataInMem_hi_lo_171};
  wire [47:0]      dataInMem_lo_460 = {dataInMem_lo_hi_268, dataRegroupBySew_0_1_30};
  wire [31:0]      dataInMem_hi_hi_364 = {dataRegroupBySew_6_1_30, dataRegroupBySew_5_1_30};
  wire [63:0]      dataInMem_hi_556 = {dataInMem_hi_hi_364, dataInMem_hi_lo_172};
  wire [47:0]      dataInMem_lo_461 = {dataInMem_lo_hi_269, dataRegroupBySew_0_1_31};
  wire [31:0]      dataInMem_hi_hi_365 = {dataRegroupBySew_6_1_31, dataRegroupBySew_5_1_31};
  wire [63:0]      dataInMem_hi_557 = {dataInMem_hi_hi_365, dataInMem_hi_lo_173};
  wire [223:0]     dataInMem_lo_lo_lo_lo_14 = {dataInMem_hi_527, dataInMem_lo_431, dataInMem_hi_526, dataInMem_lo_430};
  wire [223:0]     dataInMem_lo_lo_lo_hi_14 = {dataInMem_hi_529, dataInMem_lo_433, dataInMem_hi_528, dataInMem_lo_432};
  wire [447:0]     dataInMem_lo_lo_lo_14 = {dataInMem_lo_lo_lo_hi_14, dataInMem_lo_lo_lo_lo_14};
  wire [223:0]     dataInMem_lo_lo_hi_lo_14 = {dataInMem_hi_531, dataInMem_lo_435, dataInMem_hi_530, dataInMem_lo_434};
  wire [223:0]     dataInMem_lo_lo_hi_hi_14 = {dataInMem_hi_533, dataInMem_lo_437, dataInMem_hi_532, dataInMem_lo_436};
  wire [447:0]     dataInMem_lo_lo_hi_14 = {dataInMem_lo_lo_hi_hi_14, dataInMem_lo_lo_hi_lo_14};
  wire [895:0]     dataInMem_lo_lo_78 = {dataInMem_lo_lo_hi_14, dataInMem_lo_lo_lo_14};
  wire [223:0]     dataInMem_lo_hi_lo_lo_14 = {dataInMem_hi_535, dataInMem_lo_439, dataInMem_hi_534, dataInMem_lo_438};
  wire [223:0]     dataInMem_lo_hi_lo_hi_14 = {dataInMem_hi_537, dataInMem_lo_441, dataInMem_hi_536, dataInMem_lo_440};
  wire [447:0]     dataInMem_lo_hi_lo_14 = {dataInMem_lo_hi_lo_hi_14, dataInMem_lo_hi_lo_lo_14};
  wire [223:0]     dataInMem_lo_hi_hi_lo_14 = {dataInMem_hi_539, dataInMem_lo_443, dataInMem_hi_538, dataInMem_lo_442};
  wire [223:0]     dataInMem_lo_hi_hi_hi_14 = {dataInMem_hi_541, dataInMem_lo_445, dataInMem_hi_540, dataInMem_lo_444};
  wire [447:0]     dataInMem_lo_hi_hi_14 = {dataInMem_lo_hi_hi_hi_14, dataInMem_lo_hi_hi_lo_14};
  wire [895:0]     dataInMem_lo_hi_270 = {dataInMem_lo_hi_hi_14, dataInMem_lo_hi_lo_14};
  wire [1791:0]    dataInMem_lo_462 = {dataInMem_lo_hi_270, dataInMem_lo_lo_78};
  wire [223:0]     dataInMem_hi_lo_lo_lo_14 = {dataInMem_hi_543, dataInMem_lo_447, dataInMem_hi_542, dataInMem_lo_446};
  wire [223:0]     dataInMem_hi_lo_lo_hi_14 = {dataInMem_hi_545, dataInMem_lo_449, dataInMem_hi_544, dataInMem_lo_448};
  wire [447:0]     dataInMem_hi_lo_lo_14 = {dataInMem_hi_lo_lo_hi_14, dataInMem_hi_lo_lo_lo_14};
  wire [223:0]     dataInMem_hi_lo_hi_lo_14 = {dataInMem_hi_547, dataInMem_lo_451, dataInMem_hi_546, dataInMem_lo_450};
  wire [223:0]     dataInMem_hi_lo_hi_hi_14 = {dataInMem_hi_549, dataInMem_lo_453, dataInMem_hi_548, dataInMem_lo_452};
  wire [447:0]     dataInMem_hi_lo_hi_14 = {dataInMem_hi_lo_hi_hi_14, dataInMem_hi_lo_hi_lo_14};
  wire [895:0]     dataInMem_hi_lo_174 = {dataInMem_hi_lo_hi_14, dataInMem_hi_lo_lo_14};
  wire [223:0]     dataInMem_hi_hi_lo_lo_14 = {dataInMem_hi_551, dataInMem_lo_455, dataInMem_hi_550, dataInMem_lo_454};
  wire [223:0]     dataInMem_hi_hi_lo_hi_14 = {dataInMem_hi_553, dataInMem_lo_457, dataInMem_hi_552, dataInMem_lo_456};
  wire [447:0]     dataInMem_hi_hi_lo_14 = {dataInMem_hi_hi_lo_hi_14, dataInMem_hi_hi_lo_lo_14};
  wire [223:0]     dataInMem_hi_hi_hi_lo_14 = {dataInMem_hi_555, dataInMem_lo_459, dataInMem_hi_554, dataInMem_lo_458};
  wire [223:0]     dataInMem_hi_hi_hi_hi_14 = {dataInMem_hi_557, dataInMem_lo_461, dataInMem_hi_556, dataInMem_lo_460};
  wire [447:0]     dataInMem_hi_hi_hi_14 = {dataInMem_hi_hi_hi_hi_14, dataInMem_hi_hi_hi_lo_14};
  wire [895:0]     dataInMem_hi_hi_366 = {dataInMem_hi_hi_hi_14, dataInMem_hi_hi_lo_14};
  wire [1791:0]    dataInMem_hi_558 = {dataInMem_hi_hi_366, dataInMem_hi_lo_174};
  wire [3583:0]    dataInMem_14 = {dataInMem_hi_558, dataInMem_lo_462};
  wire [511:0]     regroupCacheLine_14_0 = dataInMem_14[511:0];
  wire [511:0]     regroupCacheLine_14_1 = dataInMem_14[1023:512];
  wire [511:0]     regroupCacheLine_14_2 = dataInMem_14[1535:1024];
  wire [511:0]     regroupCacheLine_14_3 = dataInMem_14[2047:1536];
  wire [511:0]     regroupCacheLine_14_4 = dataInMem_14[2559:2048];
  wire [511:0]     regroupCacheLine_14_5 = dataInMem_14[3071:2560];
  wire [511:0]     regroupCacheLine_14_6 = dataInMem_14[3583:3072];
  wire [511:0]     res_112 = regroupCacheLine_14_0;
  wire [511:0]     res_113 = regroupCacheLine_14_1;
  wire [511:0]     res_114 = regroupCacheLine_14_2;
  wire [511:0]     res_115 = regroupCacheLine_14_3;
  wire [511:0]     res_116 = regroupCacheLine_14_4;
  wire [511:0]     res_117 = regroupCacheLine_14_5;
  wire [511:0]     res_118 = regroupCacheLine_14_6;
  wire [1023:0]    lo_lo_14 = {res_113, res_112};
  wire [1023:0]    lo_hi_14 = {res_115, res_114};
  wire [2047:0]    lo_14 = {lo_hi_14, lo_lo_14};
  wire [1023:0]    hi_lo_14 = {res_117, res_116};
  wire [1023:0]    hi_hi_14 = {512'h0, res_118};
  wire [2047:0]    hi_14 = {hi_hi_14, hi_lo_14};
  wire [4095:0]    regroupLoadData_1_6 = {hi_14, lo_14};
  wire [63:0]      dataInMem_lo_463 = {dataInMem_lo_hi_271, dataInMem_lo_lo_79};
  wire [31:0]      dataInMem_hi_hi_367 = {dataRegroupBySew_7_1_0, dataRegroupBySew_6_1_0};
  wire [63:0]      dataInMem_hi_559 = {dataInMem_hi_hi_367, dataInMem_hi_lo_175};
  wire [63:0]      dataInMem_lo_464 = {dataInMem_lo_hi_272, dataInMem_lo_lo_80};
  wire [31:0]      dataInMem_hi_hi_368 = {dataRegroupBySew_7_1_1, dataRegroupBySew_6_1_1};
  wire [63:0]      dataInMem_hi_560 = {dataInMem_hi_hi_368, dataInMem_hi_lo_176};
  wire [63:0]      dataInMem_lo_465 = {dataInMem_lo_hi_273, dataInMem_lo_lo_81};
  wire [31:0]      dataInMem_hi_hi_369 = {dataRegroupBySew_7_1_2, dataRegroupBySew_6_1_2};
  wire [63:0]      dataInMem_hi_561 = {dataInMem_hi_hi_369, dataInMem_hi_lo_177};
  wire [63:0]      dataInMem_lo_466 = {dataInMem_lo_hi_274, dataInMem_lo_lo_82};
  wire [31:0]      dataInMem_hi_hi_370 = {dataRegroupBySew_7_1_3, dataRegroupBySew_6_1_3};
  wire [63:0]      dataInMem_hi_562 = {dataInMem_hi_hi_370, dataInMem_hi_lo_178};
  wire [63:0]      dataInMem_lo_467 = {dataInMem_lo_hi_275, dataInMem_lo_lo_83};
  wire [31:0]      dataInMem_hi_hi_371 = {dataRegroupBySew_7_1_4, dataRegroupBySew_6_1_4};
  wire [63:0]      dataInMem_hi_563 = {dataInMem_hi_hi_371, dataInMem_hi_lo_179};
  wire [63:0]      dataInMem_lo_468 = {dataInMem_lo_hi_276, dataInMem_lo_lo_84};
  wire [31:0]      dataInMem_hi_hi_372 = {dataRegroupBySew_7_1_5, dataRegroupBySew_6_1_5};
  wire [63:0]      dataInMem_hi_564 = {dataInMem_hi_hi_372, dataInMem_hi_lo_180};
  wire [63:0]      dataInMem_lo_469 = {dataInMem_lo_hi_277, dataInMem_lo_lo_85};
  wire [31:0]      dataInMem_hi_hi_373 = {dataRegroupBySew_7_1_6, dataRegroupBySew_6_1_6};
  wire [63:0]      dataInMem_hi_565 = {dataInMem_hi_hi_373, dataInMem_hi_lo_181};
  wire [63:0]      dataInMem_lo_470 = {dataInMem_lo_hi_278, dataInMem_lo_lo_86};
  wire [31:0]      dataInMem_hi_hi_374 = {dataRegroupBySew_7_1_7, dataRegroupBySew_6_1_7};
  wire [63:0]      dataInMem_hi_566 = {dataInMem_hi_hi_374, dataInMem_hi_lo_182};
  wire [63:0]      dataInMem_lo_471 = {dataInMem_lo_hi_279, dataInMem_lo_lo_87};
  wire [31:0]      dataInMem_hi_hi_375 = {dataRegroupBySew_7_1_8, dataRegroupBySew_6_1_8};
  wire [63:0]      dataInMem_hi_567 = {dataInMem_hi_hi_375, dataInMem_hi_lo_183};
  wire [63:0]      dataInMem_lo_472 = {dataInMem_lo_hi_280, dataInMem_lo_lo_88};
  wire [31:0]      dataInMem_hi_hi_376 = {dataRegroupBySew_7_1_9, dataRegroupBySew_6_1_9};
  wire [63:0]      dataInMem_hi_568 = {dataInMem_hi_hi_376, dataInMem_hi_lo_184};
  wire [63:0]      dataInMem_lo_473 = {dataInMem_lo_hi_281, dataInMem_lo_lo_89};
  wire [31:0]      dataInMem_hi_hi_377 = {dataRegroupBySew_7_1_10, dataRegroupBySew_6_1_10};
  wire [63:0]      dataInMem_hi_569 = {dataInMem_hi_hi_377, dataInMem_hi_lo_185};
  wire [63:0]      dataInMem_lo_474 = {dataInMem_lo_hi_282, dataInMem_lo_lo_90};
  wire [31:0]      dataInMem_hi_hi_378 = {dataRegroupBySew_7_1_11, dataRegroupBySew_6_1_11};
  wire [63:0]      dataInMem_hi_570 = {dataInMem_hi_hi_378, dataInMem_hi_lo_186};
  wire [63:0]      dataInMem_lo_475 = {dataInMem_lo_hi_283, dataInMem_lo_lo_91};
  wire [31:0]      dataInMem_hi_hi_379 = {dataRegroupBySew_7_1_12, dataRegroupBySew_6_1_12};
  wire [63:0]      dataInMem_hi_571 = {dataInMem_hi_hi_379, dataInMem_hi_lo_187};
  wire [63:0]      dataInMem_lo_476 = {dataInMem_lo_hi_284, dataInMem_lo_lo_92};
  wire [31:0]      dataInMem_hi_hi_380 = {dataRegroupBySew_7_1_13, dataRegroupBySew_6_1_13};
  wire [63:0]      dataInMem_hi_572 = {dataInMem_hi_hi_380, dataInMem_hi_lo_188};
  wire [63:0]      dataInMem_lo_477 = {dataInMem_lo_hi_285, dataInMem_lo_lo_93};
  wire [31:0]      dataInMem_hi_hi_381 = {dataRegroupBySew_7_1_14, dataRegroupBySew_6_1_14};
  wire [63:0]      dataInMem_hi_573 = {dataInMem_hi_hi_381, dataInMem_hi_lo_189};
  wire [63:0]      dataInMem_lo_478 = {dataInMem_lo_hi_286, dataInMem_lo_lo_94};
  wire [31:0]      dataInMem_hi_hi_382 = {dataRegroupBySew_7_1_15, dataRegroupBySew_6_1_15};
  wire [63:0]      dataInMem_hi_574 = {dataInMem_hi_hi_382, dataInMem_hi_lo_190};
  wire [63:0]      dataInMem_lo_479 = {dataInMem_lo_hi_287, dataInMem_lo_lo_95};
  wire [31:0]      dataInMem_hi_hi_383 = {dataRegroupBySew_7_1_16, dataRegroupBySew_6_1_16};
  wire [63:0]      dataInMem_hi_575 = {dataInMem_hi_hi_383, dataInMem_hi_lo_191};
  wire [63:0]      dataInMem_lo_480 = {dataInMem_lo_hi_288, dataInMem_lo_lo_96};
  wire [31:0]      dataInMem_hi_hi_384 = {dataRegroupBySew_7_1_17, dataRegroupBySew_6_1_17};
  wire [63:0]      dataInMem_hi_576 = {dataInMem_hi_hi_384, dataInMem_hi_lo_192};
  wire [63:0]      dataInMem_lo_481 = {dataInMem_lo_hi_289, dataInMem_lo_lo_97};
  wire [31:0]      dataInMem_hi_hi_385 = {dataRegroupBySew_7_1_18, dataRegroupBySew_6_1_18};
  wire [63:0]      dataInMem_hi_577 = {dataInMem_hi_hi_385, dataInMem_hi_lo_193};
  wire [63:0]      dataInMem_lo_482 = {dataInMem_lo_hi_290, dataInMem_lo_lo_98};
  wire [31:0]      dataInMem_hi_hi_386 = {dataRegroupBySew_7_1_19, dataRegroupBySew_6_1_19};
  wire [63:0]      dataInMem_hi_578 = {dataInMem_hi_hi_386, dataInMem_hi_lo_194};
  wire [63:0]      dataInMem_lo_483 = {dataInMem_lo_hi_291, dataInMem_lo_lo_99};
  wire [31:0]      dataInMem_hi_hi_387 = {dataRegroupBySew_7_1_20, dataRegroupBySew_6_1_20};
  wire [63:0]      dataInMem_hi_579 = {dataInMem_hi_hi_387, dataInMem_hi_lo_195};
  wire [63:0]      dataInMem_lo_484 = {dataInMem_lo_hi_292, dataInMem_lo_lo_100};
  wire [31:0]      dataInMem_hi_hi_388 = {dataRegroupBySew_7_1_21, dataRegroupBySew_6_1_21};
  wire [63:0]      dataInMem_hi_580 = {dataInMem_hi_hi_388, dataInMem_hi_lo_196};
  wire [63:0]      dataInMem_lo_485 = {dataInMem_lo_hi_293, dataInMem_lo_lo_101};
  wire [31:0]      dataInMem_hi_hi_389 = {dataRegroupBySew_7_1_22, dataRegroupBySew_6_1_22};
  wire [63:0]      dataInMem_hi_581 = {dataInMem_hi_hi_389, dataInMem_hi_lo_197};
  wire [63:0]      dataInMem_lo_486 = {dataInMem_lo_hi_294, dataInMem_lo_lo_102};
  wire [31:0]      dataInMem_hi_hi_390 = {dataRegroupBySew_7_1_23, dataRegroupBySew_6_1_23};
  wire [63:0]      dataInMem_hi_582 = {dataInMem_hi_hi_390, dataInMem_hi_lo_198};
  wire [63:0]      dataInMem_lo_487 = {dataInMem_lo_hi_295, dataInMem_lo_lo_103};
  wire [31:0]      dataInMem_hi_hi_391 = {dataRegroupBySew_7_1_24, dataRegroupBySew_6_1_24};
  wire [63:0]      dataInMem_hi_583 = {dataInMem_hi_hi_391, dataInMem_hi_lo_199};
  wire [63:0]      dataInMem_lo_488 = {dataInMem_lo_hi_296, dataInMem_lo_lo_104};
  wire [31:0]      dataInMem_hi_hi_392 = {dataRegroupBySew_7_1_25, dataRegroupBySew_6_1_25};
  wire [63:0]      dataInMem_hi_584 = {dataInMem_hi_hi_392, dataInMem_hi_lo_200};
  wire [63:0]      dataInMem_lo_489 = {dataInMem_lo_hi_297, dataInMem_lo_lo_105};
  wire [31:0]      dataInMem_hi_hi_393 = {dataRegroupBySew_7_1_26, dataRegroupBySew_6_1_26};
  wire [63:0]      dataInMem_hi_585 = {dataInMem_hi_hi_393, dataInMem_hi_lo_201};
  wire [63:0]      dataInMem_lo_490 = {dataInMem_lo_hi_298, dataInMem_lo_lo_106};
  wire [31:0]      dataInMem_hi_hi_394 = {dataRegroupBySew_7_1_27, dataRegroupBySew_6_1_27};
  wire [63:0]      dataInMem_hi_586 = {dataInMem_hi_hi_394, dataInMem_hi_lo_202};
  wire [63:0]      dataInMem_lo_491 = {dataInMem_lo_hi_299, dataInMem_lo_lo_107};
  wire [31:0]      dataInMem_hi_hi_395 = {dataRegroupBySew_7_1_28, dataRegroupBySew_6_1_28};
  wire [63:0]      dataInMem_hi_587 = {dataInMem_hi_hi_395, dataInMem_hi_lo_203};
  wire [63:0]      dataInMem_lo_492 = {dataInMem_lo_hi_300, dataInMem_lo_lo_108};
  wire [31:0]      dataInMem_hi_hi_396 = {dataRegroupBySew_7_1_29, dataRegroupBySew_6_1_29};
  wire [63:0]      dataInMem_hi_588 = {dataInMem_hi_hi_396, dataInMem_hi_lo_204};
  wire [63:0]      dataInMem_lo_493 = {dataInMem_lo_hi_301, dataInMem_lo_lo_109};
  wire [31:0]      dataInMem_hi_hi_397 = {dataRegroupBySew_7_1_30, dataRegroupBySew_6_1_30};
  wire [63:0]      dataInMem_hi_589 = {dataInMem_hi_hi_397, dataInMem_hi_lo_205};
  wire [63:0]      dataInMem_lo_494 = {dataInMem_lo_hi_302, dataInMem_lo_lo_110};
  wire [31:0]      dataInMem_hi_hi_398 = {dataRegroupBySew_7_1_31, dataRegroupBySew_6_1_31};
  wire [63:0]      dataInMem_hi_590 = {dataInMem_hi_hi_398, dataInMem_hi_lo_206};
  wire [255:0]     dataInMem_lo_lo_lo_lo_15 = {dataInMem_hi_560, dataInMem_lo_464, dataInMem_hi_559, dataInMem_lo_463};
  wire [255:0]     dataInMem_lo_lo_lo_hi_15 = {dataInMem_hi_562, dataInMem_lo_466, dataInMem_hi_561, dataInMem_lo_465};
  wire [511:0]     dataInMem_lo_lo_lo_15 = {dataInMem_lo_lo_lo_hi_15, dataInMem_lo_lo_lo_lo_15};
  wire [255:0]     dataInMem_lo_lo_hi_lo_15 = {dataInMem_hi_564, dataInMem_lo_468, dataInMem_hi_563, dataInMem_lo_467};
  wire [255:0]     dataInMem_lo_lo_hi_hi_15 = {dataInMem_hi_566, dataInMem_lo_470, dataInMem_hi_565, dataInMem_lo_469};
  wire [511:0]     dataInMem_lo_lo_hi_15 = {dataInMem_lo_lo_hi_hi_15, dataInMem_lo_lo_hi_lo_15};
  wire [1023:0]    dataInMem_lo_lo_111 = {dataInMem_lo_lo_hi_15, dataInMem_lo_lo_lo_15};
  wire [255:0]     dataInMem_lo_hi_lo_lo_15 = {dataInMem_hi_568, dataInMem_lo_472, dataInMem_hi_567, dataInMem_lo_471};
  wire [255:0]     dataInMem_lo_hi_lo_hi_15 = {dataInMem_hi_570, dataInMem_lo_474, dataInMem_hi_569, dataInMem_lo_473};
  wire [511:0]     dataInMem_lo_hi_lo_15 = {dataInMem_lo_hi_lo_hi_15, dataInMem_lo_hi_lo_lo_15};
  wire [255:0]     dataInMem_lo_hi_hi_lo_15 = {dataInMem_hi_572, dataInMem_lo_476, dataInMem_hi_571, dataInMem_lo_475};
  wire [255:0]     dataInMem_lo_hi_hi_hi_15 = {dataInMem_hi_574, dataInMem_lo_478, dataInMem_hi_573, dataInMem_lo_477};
  wire [511:0]     dataInMem_lo_hi_hi_15 = {dataInMem_lo_hi_hi_hi_15, dataInMem_lo_hi_hi_lo_15};
  wire [1023:0]    dataInMem_lo_hi_303 = {dataInMem_lo_hi_hi_15, dataInMem_lo_hi_lo_15};
  wire [2047:0]    dataInMem_lo_495 = {dataInMem_lo_hi_303, dataInMem_lo_lo_111};
  wire [255:0]     dataInMem_hi_lo_lo_lo_15 = {dataInMem_hi_576, dataInMem_lo_480, dataInMem_hi_575, dataInMem_lo_479};
  wire [255:0]     dataInMem_hi_lo_lo_hi_15 = {dataInMem_hi_578, dataInMem_lo_482, dataInMem_hi_577, dataInMem_lo_481};
  wire [511:0]     dataInMem_hi_lo_lo_15 = {dataInMem_hi_lo_lo_hi_15, dataInMem_hi_lo_lo_lo_15};
  wire [255:0]     dataInMem_hi_lo_hi_lo_15 = {dataInMem_hi_580, dataInMem_lo_484, dataInMem_hi_579, dataInMem_lo_483};
  wire [255:0]     dataInMem_hi_lo_hi_hi_15 = {dataInMem_hi_582, dataInMem_lo_486, dataInMem_hi_581, dataInMem_lo_485};
  wire [511:0]     dataInMem_hi_lo_hi_15 = {dataInMem_hi_lo_hi_hi_15, dataInMem_hi_lo_hi_lo_15};
  wire [1023:0]    dataInMem_hi_lo_207 = {dataInMem_hi_lo_hi_15, dataInMem_hi_lo_lo_15};
  wire [255:0]     dataInMem_hi_hi_lo_lo_15 = {dataInMem_hi_584, dataInMem_lo_488, dataInMem_hi_583, dataInMem_lo_487};
  wire [255:0]     dataInMem_hi_hi_lo_hi_15 = {dataInMem_hi_586, dataInMem_lo_490, dataInMem_hi_585, dataInMem_lo_489};
  wire [511:0]     dataInMem_hi_hi_lo_15 = {dataInMem_hi_hi_lo_hi_15, dataInMem_hi_hi_lo_lo_15};
  wire [255:0]     dataInMem_hi_hi_hi_lo_15 = {dataInMem_hi_588, dataInMem_lo_492, dataInMem_hi_587, dataInMem_lo_491};
  wire [255:0]     dataInMem_hi_hi_hi_hi_15 = {dataInMem_hi_590, dataInMem_lo_494, dataInMem_hi_589, dataInMem_lo_493};
  wire [511:0]     dataInMem_hi_hi_hi_15 = {dataInMem_hi_hi_hi_hi_15, dataInMem_hi_hi_hi_lo_15};
  wire [1023:0]    dataInMem_hi_hi_399 = {dataInMem_hi_hi_hi_15, dataInMem_hi_hi_lo_15};
  wire [2047:0]    dataInMem_hi_591 = {dataInMem_hi_hi_399, dataInMem_hi_lo_207};
  wire [4095:0]    dataInMem_15 = {dataInMem_hi_591, dataInMem_lo_495};
  wire [511:0]     regroupCacheLine_15_0 = dataInMem_15[511:0];
  wire [511:0]     regroupCacheLine_15_1 = dataInMem_15[1023:512];
  wire [511:0]     regroupCacheLine_15_2 = dataInMem_15[1535:1024];
  wire [511:0]     regroupCacheLine_15_3 = dataInMem_15[2047:1536];
  wire [511:0]     regroupCacheLine_15_4 = dataInMem_15[2559:2048];
  wire [511:0]     regroupCacheLine_15_5 = dataInMem_15[3071:2560];
  wire [511:0]     regroupCacheLine_15_6 = dataInMem_15[3583:3072];
  wire [511:0]     regroupCacheLine_15_7 = dataInMem_15[4095:3584];
  wire [511:0]     res_120 = regroupCacheLine_15_0;
  wire [511:0]     res_121 = regroupCacheLine_15_1;
  wire [511:0]     res_122 = regroupCacheLine_15_2;
  wire [511:0]     res_123 = regroupCacheLine_15_3;
  wire [511:0]     res_124 = regroupCacheLine_15_4;
  wire [511:0]     res_125 = regroupCacheLine_15_5;
  wire [511:0]     res_126 = regroupCacheLine_15_6;
  wire [511:0]     res_127 = regroupCacheLine_15_7;
  wire [1023:0]    lo_lo_15 = {res_121, res_120};
  wire [1023:0]    lo_hi_15 = {res_123, res_122};
  wire [2047:0]    lo_15 = {lo_hi_15, lo_lo_15};
  wire [1023:0]    hi_lo_15 = {res_125, res_124};
  wire [1023:0]    hi_hi_15 = {res_127, res_126};
  wire [2047:0]    hi_15 = {hi_hi_15, hi_lo_15};
  wire [4095:0]    regroupLoadData_1_7 = {hi_15, lo_15};
  wire [31:0]      dataRegroupBySew_0_2_0 = bufferStageEnqueueData_0[31:0];
  wire [31:0]      dataRegroupBySew_0_2_1 = bufferStageEnqueueData_0[63:32];
  wire [31:0]      dataRegroupBySew_0_2_2 = bufferStageEnqueueData_0[95:64];
  wire [31:0]      dataRegroupBySew_0_2_3 = bufferStageEnqueueData_0[127:96];
  wire [31:0]      dataRegroupBySew_0_2_4 = bufferStageEnqueueData_0[159:128];
  wire [31:0]      dataRegroupBySew_0_2_5 = bufferStageEnqueueData_0[191:160];
  wire [31:0]      dataRegroupBySew_0_2_6 = bufferStageEnqueueData_0[223:192];
  wire [31:0]      dataRegroupBySew_0_2_7 = bufferStageEnqueueData_0[255:224];
  wire [31:0]      dataRegroupBySew_0_2_8 = bufferStageEnqueueData_0[287:256];
  wire [31:0]      dataRegroupBySew_0_2_9 = bufferStageEnqueueData_0[319:288];
  wire [31:0]      dataRegroupBySew_0_2_10 = bufferStageEnqueueData_0[351:320];
  wire [31:0]      dataRegroupBySew_0_2_11 = bufferStageEnqueueData_0[383:352];
  wire [31:0]      dataRegroupBySew_0_2_12 = bufferStageEnqueueData_0[415:384];
  wire [31:0]      dataRegroupBySew_0_2_13 = bufferStageEnqueueData_0[447:416];
  wire [31:0]      dataRegroupBySew_0_2_14 = bufferStageEnqueueData_0[479:448];
  wire [31:0]      dataRegroupBySew_0_2_15 = bufferStageEnqueueData_0[511:480];
  wire [31:0]      dataRegroupBySew_1_2_0 = bufferStageEnqueueData_1[31:0];
  wire [31:0]      dataRegroupBySew_1_2_1 = bufferStageEnqueueData_1[63:32];
  wire [31:0]      dataRegroupBySew_1_2_2 = bufferStageEnqueueData_1[95:64];
  wire [31:0]      dataRegroupBySew_1_2_3 = bufferStageEnqueueData_1[127:96];
  wire [31:0]      dataRegroupBySew_1_2_4 = bufferStageEnqueueData_1[159:128];
  wire [31:0]      dataRegroupBySew_1_2_5 = bufferStageEnqueueData_1[191:160];
  wire [31:0]      dataRegroupBySew_1_2_6 = bufferStageEnqueueData_1[223:192];
  wire [31:0]      dataRegroupBySew_1_2_7 = bufferStageEnqueueData_1[255:224];
  wire [31:0]      dataRegroupBySew_1_2_8 = bufferStageEnqueueData_1[287:256];
  wire [31:0]      dataRegroupBySew_1_2_9 = bufferStageEnqueueData_1[319:288];
  wire [31:0]      dataRegroupBySew_1_2_10 = bufferStageEnqueueData_1[351:320];
  wire [31:0]      dataRegroupBySew_1_2_11 = bufferStageEnqueueData_1[383:352];
  wire [31:0]      dataRegroupBySew_1_2_12 = bufferStageEnqueueData_1[415:384];
  wire [31:0]      dataRegroupBySew_1_2_13 = bufferStageEnqueueData_1[447:416];
  wire [31:0]      dataRegroupBySew_1_2_14 = bufferStageEnqueueData_1[479:448];
  wire [31:0]      dataRegroupBySew_1_2_15 = bufferStageEnqueueData_1[511:480];
  wire [31:0]      dataRegroupBySew_2_2_0 = bufferStageEnqueueData_2[31:0];
  wire [31:0]      dataRegroupBySew_2_2_1 = bufferStageEnqueueData_2[63:32];
  wire [31:0]      dataRegroupBySew_2_2_2 = bufferStageEnqueueData_2[95:64];
  wire [31:0]      dataRegroupBySew_2_2_3 = bufferStageEnqueueData_2[127:96];
  wire [31:0]      dataRegroupBySew_2_2_4 = bufferStageEnqueueData_2[159:128];
  wire [31:0]      dataRegroupBySew_2_2_5 = bufferStageEnqueueData_2[191:160];
  wire [31:0]      dataRegroupBySew_2_2_6 = bufferStageEnqueueData_2[223:192];
  wire [31:0]      dataRegroupBySew_2_2_7 = bufferStageEnqueueData_2[255:224];
  wire [31:0]      dataRegroupBySew_2_2_8 = bufferStageEnqueueData_2[287:256];
  wire [31:0]      dataRegroupBySew_2_2_9 = bufferStageEnqueueData_2[319:288];
  wire [31:0]      dataRegroupBySew_2_2_10 = bufferStageEnqueueData_2[351:320];
  wire [31:0]      dataRegroupBySew_2_2_11 = bufferStageEnqueueData_2[383:352];
  wire [31:0]      dataRegroupBySew_2_2_12 = bufferStageEnqueueData_2[415:384];
  wire [31:0]      dataRegroupBySew_2_2_13 = bufferStageEnqueueData_2[447:416];
  wire [31:0]      dataRegroupBySew_2_2_14 = bufferStageEnqueueData_2[479:448];
  wire [31:0]      dataRegroupBySew_2_2_15 = bufferStageEnqueueData_2[511:480];
  wire [31:0]      dataRegroupBySew_3_2_0 = bufferStageEnqueueData_3[31:0];
  wire [31:0]      dataRegroupBySew_3_2_1 = bufferStageEnqueueData_3[63:32];
  wire [31:0]      dataRegroupBySew_3_2_2 = bufferStageEnqueueData_3[95:64];
  wire [31:0]      dataRegroupBySew_3_2_3 = bufferStageEnqueueData_3[127:96];
  wire [31:0]      dataRegroupBySew_3_2_4 = bufferStageEnqueueData_3[159:128];
  wire [31:0]      dataRegroupBySew_3_2_5 = bufferStageEnqueueData_3[191:160];
  wire [31:0]      dataRegroupBySew_3_2_6 = bufferStageEnqueueData_3[223:192];
  wire [31:0]      dataRegroupBySew_3_2_7 = bufferStageEnqueueData_3[255:224];
  wire [31:0]      dataRegroupBySew_3_2_8 = bufferStageEnqueueData_3[287:256];
  wire [31:0]      dataRegroupBySew_3_2_9 = bufferStageEnqueueData_3[319:288];
  wire [31:0]      dataRegroupBySew_3_2_10 = bufferStageEnqueueData_3[351:320];
  wire [31:0]      dataRegroupBySew_3_2_11 = bufferStageEnqueueData_3[383:352];
  wire [31:0]      dataRegroupBySew_3_2_12 = bufferStageEnqueueData_3[415:384];
  wire [31:0]      dataRegroupBySew_3_2_13 = bufferStageEnqueueData_3[447:416];
  wire [31:0]      dataRegroupBySew_3_2_14 = bufferStageEnqueueData_3[479:448];
  wire [31:0]      dataRegroupBySew_3_2_15 = bufferStageEnqueueData_3[511:480];
  wire [31:0]      dataRegroupBySew_4_2_0 = bufferStageEnqueueData_4[31:0];
  wire [31:0]      dataRegroupBySew_4_2_1 = bufferStageEnqueueData_4[63:32];
  wire [31:0]      dataRegroupBySew_4_2_2 = bufferStageEnqueueData_4[95:64];
  wire [31:0]      dataRegroupBySew_4_2_3 = bufferStageEnqueueData_4[127:96];
  wire [31:0]      dataRegroupBySew_4_2_4 = bufferStageEnqueueData_4[159:128];
  wire [31:0]      dataRegroupBySew_4_2_5 = bufferStageEnqueueData_4[191:160];
  wire [31:0]      dataRegroupBySew_4_2_6 = bufferStageEnqueueData_4[223:192];
  wire [31:0]      dataRegroupBySew_4_2_7 = bufferStageEnqueueData_4[255:224];
  wire [31:0]      dataRegroupBySew_4_2_8 = bufferStageEnqueueData_4[287:256];
  wire [31:0]      dataRegroupBySew_4_2_9 = bufferStageEnqueueData_4[319:288];
  wire [31:0]      dataRegroupBySew_4_2_10 = bufferStageEnqueueData_4[351:320];
  wire [31:0]      dataRegroupBySew_4_2_11 = bufferStageEnqueueData_4[383:352];
  wire [31:0]      dataRegroupBySew_4_2_12 = bufferStageEnqueueData_4[415:384];
  wire [31:0]      dataRegroupBySew_4_2_13 = bufferStageEnqueueData_4[447:416];
  wire [31:0]      dataRegroupBySew_4_2_14 = bufferStageEnqueueData_4[479:448];
  wire [31:0]      dataRegroupBySew_4_2_15 = bufferStageEnqueueData_4[511:480];
  wire [31:0]      dataRegroupBySew_5_2_0 = bufferStageEnqueueData_5[31:0];
  wire [31:0]      dataRegroupBySew_5_2_1 = bufferStageEnqueueData_5[63:32];
  wire [31:0]      dataRegroupBySew_5_2_2 = bufferStageEnqueueData_5[95:64];
  wire [31:0]      dataRegroupBySew_5_2_3 = bufferStageEnqueueData_5[127:96];
  wire [31:0]      dataRegroupBySew_5_2_4 = bufferStageEnqueueData_5[159:128];
  wire [31:0]      dataRegroupBySew_5_2_5 = bufferStageEnqueueData_5[191:160];
  wire [31:0]      dataRegroupBySew_5_2_6 = bufferStageEnqueueData_5[223:192];
  wire [31:0]      dataRegroupBySew_5_2_7 = bufferStageEnqueueData_5[255:224];
  wire [31:0]      dataRegroupBySew_5_2_8 = bufferStageEnqueueData_5[287:256];
  wire [31:0]      dataRegroupBySew_5_2_9 = bufferStageEnqueueData_5[319:288];
  wire [31:0]      dataRegroupBySew_5_2_10 = bufferStageEnqueueData_5[351:320];
  wire [31:0]      dataRegroupBySew_5_2_11 = bufferStageEnqueueData_5[383:352];
  wire [31:0]      dataRegroupBySew_5_2_12 = bufferStageEnqueueData_5[415:384];
  wire [31:0]      dataRegroupBySew_5_2_13 = bufferStageEnqueueData_5[447:416];
  wire [31:0]      dataRegroupBySew_5_2_14 = bufferStageEnqueueData_5[479:448];
  wire [31:0]      dataRegroupBySew_5_2_15 = bufferStageEnqueueData_5[511:480];
  wire [31:0]      dataRegroupBySew_6_2_0 = bufferStageEnqueueData_6[31:0];
  wire [31:0]      dataRegroupBySew_6_2_1 = bufferStageEnqueueData_6[63:32];
  wire [31:0]      dataRegroupBySew_6_2_2 = bufferStageEnqueueData_6[95:64];
  wire [31:0]      dataRegroupBySew_6_2_3 = bufferStageEnqueueData_6[127:96];
  wire [31:0]      dataRegroupBySew_6_2_4 = bufferStageEnqueueData_6[159:128];
  wire [31:0]      dataRegroupBySew_6_2_5 = bufferStageEnqueueData_6[191:160];
  wire [31:0]      dataRegroupBySew_6_2_6 = bufferStageEnqueueData_6[223:192];
  wire [31:0]      dataRegroupBySew_6_2_7 = bufferStageEnqueueData_6[255:224];
  wire [31:0]      dataRegroupBySew_6_2_8 = bufferStageEnqueueData_6[287:256];
  wire [31:0]      dataRegroupBySew_6_2_9 = bufferStageEnqueueData_6[319:288];
  wire [31:0]      dataRegroupBySew_6_2_10 = bufferStageEnqueueData_6[351:320];
  wire [31:0]      dataRegroupBySew_6_2_11 = bufferStageEnqueueData_6[383:352];
  wire [31:0]      dataRegroupBySew_6_2_12 = bufferStageEnqueueData_6[415:384];
  wire [31:0]      dataRegroupBySew_6_2_13 = bufferStageEnqueueData_6[447:416];
  wire [31:0]      dataRegroupBySew_6_2_14 = bufferStageEnqueueData_6[479:448];
  wire [31:0]      dataRegroupBySew_6_2_15 = bufferStageEnqueueData_6[511:480];
  wire [31:0]      dataRegroupBySew_7_2_0 = bufferStageEnqueueData_7[31:0];
  wire [31:0]      dataRegroupBySew_7_2_1 = bufferStageEnqueueData_7[63:32];
  wire [31:0]      dataRegroupBySew_7_2_2 = bufferStageEnqueueData_7[95:64];
  wire [31:0]      dataRegroupBySew_7_2_3 = bufferStageEnqueueData_7[127:96];
  wire [31:0]      dataRegroupBySew_7_2_4 = bufferStageEnqueueData_7[159:128];
  wire [31:0]      dataRegroupBySew_7_2_5 = bufferStageEnqueueData_7[191:160];
  wire [31:0]      dataRegroupBySew_7_2_6 = bufferStageEnqueueData_7[223:192];
  wire [31:0]      dataRegroupBySew_7_2_7 = bufferStageEnqueueData_7[255:224];
  wire [31:0]      dataRegroupBySew_7_2_8 = bufferStageEnqueueData_7[287:256];
  wire [31:0]      dataRegroupBySew_7_2_9 = bufferStageEnqueueData_7[319:288];
  wire [31:0]      dataRegroupBySew_7_2_10 = bufferStageEnqueueData_7[351:320];
  wire [31:0]      dataRegroupBySew_7_2_11 = bufferStageEnqueueData_7[383:352];
  wire [31:0]      dataRegroupBySew_7_2_12 = bufferStageEnqueueData_7[415:384];
  wire [31:0]      dataRegroupBySew_7_2_13 = bufferStageEnqueueData_7[447:416];
  wire [31:0]      dataRegroupBySew_7_2_14 = bufferStageEnqueueData_7[479:448];
  wire [31:0]      dataRegroupBySew_7_2_15 = bufferStageEnqueueData_7[511:480];
  wire [63:0]      dataInMem_lo_lo_lo_16 = {dataRegroupBySew_0_2_1, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_lo_lo_hi_16 = {dataRegroupBySew_0_2_3, dataRegroupBySew_0_2_2};
  wire [127:0]     dataInMem_lo_lo_112 = {dataInMem_lo_lo_hi_16, dataInMem_lo_lo_lo_16};
  wire [63:0]      dataInMem_lo_hi_lo_16 = {dataRegroupBySew_0_2_5, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_lo_hi_hi_16 = {dataRegroupBySew_0_2_7, dataRegroupBySew_0_2_6};
  wire [127:0]     dataInMem_lo_hi_304 = {dataInMem_lo_hi_hi_16, dataInMem_lo_hi_lo_16};
  wire [255:0]     dataInMem_lo_496 = {dataInMem_lo_hi_304, dataInMem_lo_lo_112};
  wire [63:0]      dataInMem_hi_lo_lo_16 = {dataRegroupBySew_0_2_9, dataRegroupBySew_0_2_8};
  wire [63:0]      dataInMem_hi_lo_hi_16 = {dataRegroupBySew_0_2_11, dataRegroupBySew_0_2_10};
  wire [127:0]     dataInMem_hi_lo_208 = {dataInMem_hi_lo_hi_16, dataInMem_hi_lo_lo_16};
  wire [63:0]      dataInMem_hi_hi_lo_16 = {dataRegroupBySew_0_2_13, dataRegroupBySew_0_2_12};
  wire [63:0]      dataInMem_hi_hi_hi_16 = {dataRegroupBySew_0_2_15, dataRegroupBySew_0_2_14};
  wire [127:0]     dataInMem_hi_hi_400 = {dataInMem_hi_hi_hi_16, dataInMem_hi_hi_lo_16};
  wire [255:0]     dataInMem_hi_592 = {dataInMem_hi_hi_400, dataInMem_hi_lo_208};
  wire [511:0]     dataInMem_16 = {dataInMem_hi_592, dataInMem_lo_496};
  wire [511:0]     regroupCacheLine_16_0 = dataInMem_16;
  wire [511:0]     res_128 = regroupCacheLine_16_0;
  wire [1023:0]    lo_lo_16 = {512'h0, res_128};
  wire [2047:0]    lo_16 = {1024'h0, lo_lo_16};
  wire [4095:0]    regroupLoadData_2_0 = {2048'h0, lo_16};
  wire [127:0]     dataInMem_lo_lo_lo_17 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1, dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [127:0]     dataInMem_lo_lo_hi_17 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3, dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [255:0]     dataInMem_lo_lo_113 = {dataInMem_lo_lo_hi_17, dataInMem_lo_lo_lo_17};
  wire [127:0]     dataInMem_lo_hi_lo_17 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5, dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [127:0]     dataInMem_lo_hi_hi_17 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7, dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [255:0]     dataInMem_lo_hi_305 = {dataInMem_lo_hi_hi_17, dataInMem_lo_hi_lo_17};
  wire [511:0]     dataInMem_lo_497 = {dataInMem_lo_hi_305, dataInMem_lo_lo_113};
  wire [127:0]     dataInMem_hi_lo_lo_17 = {dataRegroupBySew_1_2_9, dataRegroupBySew_0_2_9, dataRegroupBySew_1_2_8, dataRegroupBySew_0_2_8};
  wire [127:0]     dataInMem_hi_lo_hi_17 = {dataRegroupBySew_1_2_11, dataRegroupBySew_0_2_11, dataRegroupBySew_1_2_10, dataRegroupBySew_0_2_10};
  wire [255:0]     dataInMem_hi_lo_209 = {dataInMem_hi_lo_hi_17, dataInMem_hi_lo_lo_17};
  wire [127:0]     dataInMem_hi_hi_lo_17 = {dataRegroupBySew_1_2_13, dataRegroupBySew_0_2_13, dataRegroupBySew_1_2_12, dataRegroupBySew_0_2_12};
  wire [127:0]     dataInMem_hi_hi_hi_17 = {dataRegroupBySew_1_2_15, dataRegroupBySew_0_2_15, dataRegroupBySew_1_2_14, dataRegroupBySew_0_2_14};
  wire [255:0]     dataInMem_hi_hi_401 = {dataInMem_hi_hi_hi_17, dataInMem_hi_hi_lo_17};
  wire [511:0]     dataInMem_hi_593 = {dataInMem_hi_hi_401, dataInMem_hi_lo_209};
  wire [1023:0]    dataInMem_17 = {dataInMem_hi_593, dataInMem_lo_497};
  wire [511:0]     regroupCacheLine_17_0 = dataInMem_17[511:0];
  wire [511:0]     regroupCacheLine_17_1 = dataInMem_17[1023:512];
  wire [511:0]     res_136 = regroupCacheLine_17_0;
  wire [511:0]     res_137 = regroupCacheLine_17_1;
  wire [1023:0]    lo_lo_17 = {res_137, res_136};
  wire [2047:0]    lo_17 = {1024'h0, lo_lo_17};
  wire [4095:0]    regroupLoadData_2_1 = {2048'h0, lo_17};
  wire [63:0]      _GEN_485 = {dataRegroupBySew_2_2_0, dataRegroupBySew_1_2_0};
  wire [63:0]      dataInMem_hi_594;
  assign dataInMem_hi_594 = _GEN_485;
  wire [63:0]      dataInMem_lo_hi_309;
  assign dataInMem_lo_hi_309 = _GEN_485;
  wire [63:0]      dataInMem_lo_hi_326;
  assign dataInMem_lo_hi_326 = _GEN_485;
  wire [63:0]      _GEN_486 = {dataRegroupBySew_2_2_1, dataRegroupBySew_1_2_1};
  wire [63:0]      dataInMem_hi_595;
  assign dataInMem_hi_595 = _GEN_486;
  wire [63:0]      dataInMem_lo_hi_310;
  assign dataInMem_lo_hi_310 = _GEN_486;
  wire [63:0]      dataInMem_lo_hi_327;
  assign dataInMem_lo_hi_327 = _GEN_486;
  wire [63:0]      _GEN_487 = {dataRegroupBySew_2_2_2, dataRegroupBySew_1_2_2};
  wire [63:0]      dataInMem_hi_596;
  assign dataInMem_hi_596 = _GEN_487;
  wire [63:0]      dataInMem_lo_hi_311;
  assign dataInMem_lo_hi_311 = _GEN_487;
  wire [63:0]      dataInMem_lo_hi_328;
  assign dataInMem_lo_hi_328 = _GEN_487;
  wire [63:0]      _GEN_488 = {dataRegroupBySew_2_2_3, dataRegroupBySew_1_2_3};
  wire [63:0]      dataInMem_hi_597;
  assign dataInMem_hi_597 = _GEN_488;
  wire [63:0]      dataInMem_lo_hi_312;
  assign dataInMem_lo_hi_312 = _GEN_488;
  wire [63:0]      dataInMem_lo_hi_329;
  assign dataInMem_lo_hi_329 = _GEN_488;
  wire [63:0]      _GEN_489 = {dataRegroupBySew_2_2_4, dataRegroupBySew_1_2_4};
  wire [63:0]      dataInMem_hi_598;
  assign dataInMem_hi_598 = _GEN_489;
  wire [63:0]      dataInMem_lo_hi_313;
  assign dataInMem_lo_hi_313 = _GEN_489;
  wire [63:0]      dataInMem_lo_hi_330;
  assign dataInMem_lo_hi_330 = _GEN_489;
  wire [63:0]      _GEN_490 = {dataRegroupBySew_2_2_5, dataRegroupBySew_1_2_5};
  wire [63:0]      dataInMem_hi_599;
  assign dataInMem_hi_599 = _GEN_490;
  wire [63:0]      dataInMem_lo_hi_314;
  assign dataInMem_lo_hi_314 = _GEN_490;
  wire [63:0]      dataInMem_lo_hi_331;
  assign dataInMem_lo_hi_331 = _GEN_490;
  wire [63:0]      _GEN_491 = {dataRegroupBySew_2_2_6, dataRegroupBySew_1_2_6};
  wire [63:0]      dataInMem_hi_600;
  assign dataInMem_hi_600 = _GEN_491;
  wire [63:0]      dataInMem_lo_hi_315;
  assign dataInMem_lo_hi_315 = _GEN_491;
  wire [63:0]      dataInMem_lo_hi_332;
  assign dataInMem_lo_hi_332 = _GEN_491;
  wire [63:0]      _GEN_492 = {dataRegroupBySew_2_2_7, dataRegroupBySew_1_2_7};
  wire [63:0]      dataInMem_hi_601;
  assign dataInMem_hi_601 = _GEN_492;
  wire [63:0]      dataInMem_lo_hi_316;
  assign dataInMem_lo_hi_316 = _GEN_492;
  wire [63:0]      dataInMem_lo_hi_333;
  assign dataInMem_lo_hi_333 = _GEN_492;
  wire [63:0]      _GEN_493 = {dataRegroupBySew_2_2_8, dataRegroupBySew_1_2_8};
  wire [63:0]      dataInMem_hi_602;
  assign dataInMem_hi_602 = _GEN_493;
  wire [63:0]      dataInMem_lo_hi_317;
  assign dataInMem_lo_hi_317 = _GEN_493;
  wire [63:0]      dataInMem_lo_hi_334;
  assign dataInMem_lo_hi_334 = _GEN_493;
  wire [63:0]      _GEN_494 = {dataRegroupBySew_2_2_9, dataRegroupBySew_1_2_9};
  wire [63:0]      dataInMem_hi_603;
  assign dataInMem_hi_603 = _GEN_494;
  wire [63:0]      dataInMem_lo_hi_318;
  assign dataInMem_lo_hi_318 = _GEN_494;
  wire [63:0]      dataInMem_lo_hi_335;
  assign dataInMem_lo_hi_335 = _GEN_494;
  wire [63:0]      _GEN_495 = {dataRegroupBySew_2_2_10, dataRegroupBySew_1_2_10};
  wire [63:0]      dataInMem_hi_604;
  assign dataInMem_hi_604 = _GEN_495;
  wire [63:0]      dataInMem_lo_hi_319;
  assign dataInMem_lo_hi_319 = _GEN_495;
  wire [63:0]      dataInMem_lo_hi_336;
  assign dataInMem_lo_hi_336 = _GEN_495;
  wire [63:0]      _GEN_496 = {dataRegroupBySew_2_2_11, dataRegroupBySew_1_2_11};
  wire [63:0]      dataInMem_hi_605;
  assign dataInMem_hi_605 = _GEN_496;
  wire [63:0]      dataInMem_lo_hi_320;
  assign dataInMem_lo_hi_320 = _GEN_496;
  wire [63:0]      dataInMem_lo_hi_337;
  assign dataInMem_lo_hi_337 = _GEN_496;
  wire [63:0]      _GEN_497 = {dataRegroupBySew_2_2_12, dataRegroupBySew_1_2_12};
  wire [63:0]      dataInMem_hi_606;
  assign dataInMem_hi_606 = _GEN_497;
  wire [63:0]      dataInMem_lo_hi_321;
  assign dataInMem_lo_hi_321 = _GEN_497;
  wire [63:0]      dataInMem_lo_hi_338;
  assign dataInMem_lo_hi_338 = _GEN_497;
  wire [63:0]      _GEN_498 = {dataRegroupBySew_2_2_13, dataRegroupBySew_1_2_13};
  wire [63:0]      dataInMem_hi_607;
  assign dataInMem_hi_607 = _GEN_498;
  wire [63:0]      dataInMem_lo_hi_322;
  assign dataInMem_lo_hi_322 = _GEN_498;
  wire [63:0]      dataInMem_lo_hi_339;
  assign dataInMem_lo_hi_339 = _GEN_498;
  wire [63:0]      _GEN_499 = {dataRegroupBySew_2_2_14, dataRegroupBySew_1_2_14};
  wire [63:0]      dataInMem_hi_608;
  assign dataInMem_hi_608 = _GEN_499;
  wire [63:0]      dataInMem_lo_hi_323;
  assign dataInMem_lo_hi_323 = _GEN_499;
  wire [63:0]      dataInMem_lo_hi_340;
  assign dataInMem_lo_hi_340 = _GEN_499;
  wire [63:0]      _GEN_500 = {dataRegroupBySew_2_2_15, dataRegroupBySew_1_2_15};
  wire [63:0]      dataInMem_hi_609;
  assign dataInMem_hi_609 = _GEN_500;
  wire [63:0]      dataInMem_lo_hi_324;
  assign dataInMem_lo_hi_324 = _GEN_500;
  wire [63:0]      dataInMem_lo_hi_341;
  assign dataInMem_lo_hi_341 = _GEN_500;
  wire [191:0]     dataInMem_lo_lo_lo_18 = {dataInMem_hi_595, dataRegroupBySew_0_2_1, dataInMem_hi_594, dataRegroupBySew_0_2_0};
  wire [191:0]     dataInMem_lo_lo_hi_18 = {dataInMem_hi_597, dataRegroupBySew_0_2_3, dataInMem_hi_596, dataRegroupBySew_0_2_2};
  wire [383:0]     dataInMem_lo_lo_114 = {dataInMem_lo_lo_hi_18, dataInMem_lo_lo_lo_18};
  wire [191:0]     dataInMem_lo_hi_lo_18 = {dataInMem_hi_599, dataRegroupBySew_0_2_5, dataInMem_hi_598, dataRegroupBySew_0_2_4};
  wire [191:0]     dataInMem_lo_hi_hi_18 = {dataInMem_hi_601, dataRegroupBySew_0_2_7, dataInMem_hi_600, dataRegroupBySew_0_2_6};
  wire [383:0]     dataInMem_lo_hi_306 = {dataInMem_lo_hi_hi_18, dataInMem_lo_hi_lo_18};
  wire [767:0]     dataInMem_lo_498 = {dataInMem_lo_hi_306, dataInMem_lo_lo_114};
  wire [191:0]     dataInMem_hi_lo_lo_18 = {dataInMem_hi_603, dataRegroupBySew_0_2_9, dataInMem_hi_602, dataRegroupBySew_0_2_8};
  wire [191:0]     dataInMem_hi_lo_hi_18 = {dataInMem_hi_605, dataRegroupBySew_0_2_11, dataInMem_hi_604, dataRegroupBySew_0_2_10};
  wire [383:0]     dataInMem_hi_lo_210 = {dataInMem_hi_lo_hi_18, dataInMem_hi_lo_lo_18};
  wire [191:0]     dataInMem_hi_hi_lo_18 = {dataInMem_hi_607, dataRegroupBySew_0_2_13, dataInMem_hi_606, dataRegroupBySew_0_2_12};
  wire [191:0]     dataInMem_hi_hi_hi_18 = {dataInMem_hi_609, dataRegroupBySew_0_2_15, dataInMem_hi_608, dataRegroupBySew_0_2_14};
  wire [383:0]     dataInMem_hi_hi_402 = {dataInMem_hi_hi_hi_18, dataInMem_hi_hi_lo_18};
  wire [767:0]     dataInMem_hi_610 = {dataInMem_hi_hi_402, dataInMem_hi_lo_210};
  wire [1535:0]    dataInMem_18 = {dataInMem_hi_610, dataInMem_lo_498};
  wire [511:0]     regroupCacheLine_18_0 = dataInMem_18[511:0];
  wire [511:0]     regroupCacheLine_18_1 = dataInMem_18[1023:512];
  wire [511:0]     regroupCacheLine_18_2 = dataInMem_18[1535:1024];
  wire [511:0]     res_144 = regroupCacheLine_18_0;
  wire [511:0]     res_145 = regroupCacheLine_18_1;
  wire [511:0]     res_146 = regroupCacheLine_18_2;
  wire [1023:0]    lo_lo_18 = {res_145, res_144};
  wire [1023:0]    lo_hi_18 = {512'h0, res_146};
  wire [2047:0]    lo_18 = {lo_hi_18, lo_lo_18};
  wire [4095:0]    regroupLoadData_2_2 = {2048'h0, lo_18};
  wire [63:0]      _GEN_501 = {dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_lo_499;
  assign dataInMem_lo_499 = _GEN_501;
  wire [63:0]      dataInMem_lo_516;
  assign dataInMem_lo_516 = _GEN_501;
  wire [63:0]      dataInMem_lo_lo_119;
  assign dataInMem_lo_lo_119 = _GEN_501;
  wire [63:0]      _GEN_502 = {dataRegroupBySew_3_2_0, dataRegroupBySew_2_2_0};
  wire [63:0]      dataInMem_hi_611;
  assign dataInMem_hi_611 = _GEN_502;
  wire [63:0]      dataInMem_lo_hi_343;
  assign dataInMem_lo_hi_343 = _GEN_502;
  wire [63:0]      _GEN_503 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_lo_500;
  assign dataInMem_lo_500 = _GEN_503;
  wire [63:0]      dataInMem_lo_517;
  assign dataInMem_lo_517 = _GEN_503;
  wire [63:0]      dataInMem_lo_lo_120;
  assign dataInMem_lo_lo_120 = _GEN_503;
  wire [63:0]      _GEN_504 = {dataRegroupBySew_3_2_1, dataRegroupBySew_2_2_1};
  wire [63:0]      dataInMem_hi_612;
  assign dataInMem_hi_612 = _GEN_504;
  wire [63:0]      dataInMem_lo_hi_344;
  assign dataInMem_lo_hi_344 = _GEN_504;
  wire [63:0]      _GEN_505 = {dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_lo_501;
  assign dataInMem_lo_501 = _GEN_505;
  wire [63:0]      dataInMem_lo_518;
  assign dataInMem_lo_518 = _GEN_505;
  wire [63:0]      dataInMem_lo_lo_121;
  assign dataInMem_lo_lo_121 = _GEN_505;
  wire [63:0]      _GEN_506 = {dataRegroupBySew_3_2_2, dataRegroupBySew_2_2_2};
  wire [63:0]      dataInMem_hi_613;
  assign dataInMem_hi_613 = _GEN_506;
  wire [63:0]      dataInMem_lo_hi_345;
  assign dataInMem_lo_hi_345 = _GEN_506;
  wire [63:0]      _GEN_507 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_lo_502;
  assign dataInMem_lo_502 = _GEN_507;
  wire [63:0]      dataInMem_lo_519;
  assign dataInMem_lo_519 = _GEN_507;
  wire [63:0]      dataInMem_lo_lo_122;
  assign dataInMem_lo_lo_122 = _GEN_507;
  wire [63:0]      _GEN_508 = {dataRegroupBySew_3_2_3, dataRegroupBySew_2_2_3};
  wire [63:0]      dataInMem_hi_614;
  assign dataInMem_hi_614 = _GEN_508;
  wire [63:0]      dataInMem_lo_hi_346;
  assign dataInMem_lo_hi_346 = _GEN_508;
  wire [63:0]      _GEN_509 = {dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_lo_503;
  assign dataInMem_lo_503 = _GEN_509;
  wire [63:0]      dataInMem_lo_520;
  assign dataInMem_lo_520 = _GEN_509;
  wire [63:0]      dataInMem_lo_lo_123;
  assign dataInMem_lo_lo_123 = _GEN_509;
  wire [63:0]      _GEN_510 = {dataRegroupBySew_3_2_4, dataRegroupBySew_2_2_4};
  wire [63:0]      dataInMem_hi_615;
  assign dataInMem_hi_615 = _GEN_510;
  wire [63:0]      dataInMem_lo_hi_347;
  assign dataInMem_lo_hi_347 = _GEN_510;
  wire [63:0]      _GEN_511 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5};
  wire [63:0]      dataInMem_lo_504;
  assign dataInMem_lo_504 = _GEN_511;
  wire [63:0]      dataInMem_lo_521;
  assign dataInMem_lo_521 = _GEN_511;
  wire [63:0]      dataInMem_lo_lo_124;
  assign dataInMem_lo_lo_124 = _GEN_511;
  wire [63:0]      _GEN_512 = {dataRegroupBySew_3_2_5, dataRegroupBySew_2_2_5};
  wire [63:0]      dataInMem_hi_616;
  assign dataInMem_hi_616 = _GEN_512;
  wire [63:0]      dataInMem_lo_hi_348;
  assign dataInMem_lo_hi_348 = _GEN_512;
  wire [63:0]      _GEN_513 = {dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [63:0]      dataInMem_lo_505;
  assign dataInMem_lo_505 = _GEN_513;
  wire [63:0]      dataInMem_lo_522;
  assign dataInMem_lo_522 = _GEN_513;
  wire [63:0]      dataInMem_lo_lo_125;
  assign dataInMem_lo_lo_125 = _GEN_513;
  wire [63:0]      _GEN_514 = {dataRegroupBySew_3_2_6, dataRegroupBySew_2_2_6};
  wire [63:0]      dataInMem_hi_617;
  assign dataInMem_hi_617 = _GEN_514;
  wire [63:0]      dataInMem_lo_hi_349;
  assign dataInMem_lo_hi_349 = _GEN_514;
  wire [63:0]      _GEN_515 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7};
  wire [63:0]      dataInMem_lo_506;
  assign dataInMem_lo_506 = _GEN_515;
  wire [63:0]      dataInMem_lo_523;
  assign dataInMem_lo_523 = _GEN_515;
  wire [63:0]      dataInMem_lo_lo_126;
  assign dataInMem_lo_lo_126 = _GEN_515;
  wire [63:0]      _GEN_516 = {dataRegroupBySew_3_2_7, dataRegroupBySew_2_2_7};
  wire [63:0]      dataInMem_hi_618;
  assign dataInMem_hi_618 = _GEN_516;
  wire [63:0]      dataInMem_lo_hi_350;
  assign dataInMem_lo_hi_350 = _GEN_516;
  wire [63:0]      _GEN_517 = {dataRegroupBySew_1_2_8, dataRegroupBySew_0_2_8};
  wire [63:0]      dataInMem_lo_507;
  assign dataInMem_lo_507 = _GEN_517;
  wire [63:0]      dataInMem_lo_524;
  assign dataInMem_lo_524 = _GEN_517;
  wire [63:0]      dataInMem_lo_lo_127;
  assign dataInMem_lo_lo_127 = _GEN_517;
  wire [63:0]      _GEN_518 = {dataRegroupBySew_3_2_8, dataRegroupBySew_2_2_8};
  wire [63:0]      dataInMem_hi_619;
  assign dataInMem_hi_619 = _GEN_518;
  wire [63:0]      dataInMem_lo_hi_351;
  assign dataInMem_lo_hi_351 = _GEN_518;
  wire [63:0]      _GEN_519 = {dataRegroupBySew_1_2_9, dataRegroupBySew_0_2_9};
  wire [63:0]      dataInMem_lo_508;
  assign dataInMem_lo_508 = _GEN_519;
  wire [63:0]      dataInMem_lo_525;
  assign dataInMem_lo_525 = _GEN_519;
  wire [63:0]      dataInMem_lo_lo_128;
  assign dataInMem_lo_lo_128 = _GEN_519;
  wire [63:0]      _GEN_520 = {dataRegroupBySew_3_2_9, dataRegroupBySew_2_2_9};
  wire [63:0]      dataInMem_hi_620;
  assign dataInMem_hi_620 = _GEN_520;
  wire [63:0]      dataInMem_lo_hi_352;
  assign dataInMem_lo_hi_352 = _GEN_520;
  wire [63:0]      _GEN_521 = {dataRegroupBySew_1_2_10, dataRegroupBySew_0_2_10};
  wire [63:0]      dataInMem_lo_509;
  assign dataInMem_lo_509 = _GEN_521;
  wire [63:0]      dataInMem_lo_526;
  assign dataInMem_lo_526 = _GEN_521;
  wire [63:0]      dataInMem_lo_lo_129;
  assign dataInMem_lo_lo_129 = _GEN_521;
  wire [63:0]      _GEN_522 = {dataRegroupBySew_3_2_10, dataRegroupBySew_2_2_10};
  wire [63:0]      dataInMem_hi_621;
  assign dataInMem_hi_621 = _GEN_522;
  wire [63:0]      dataInMem_lo_hi_353;
  assign dataInMem_lo_hi_353 = _GEN_522;
  wire [63:0]      _GEN_523 = {dataRegroupBySew_1_2_11, dataRegroupBySew_0_2_11};
  wire [63:0]      dataInMem_lo_510;
  assign dataInMem_lo_510 = _GEN_523;
  wire [63:0]      dataInMem_lo_527;
  assign dataInMem_lo_527 = _GEN_523;
  wire [63:0]      dataInMem_lo_lo_130;
  assign dataInMem_lo_lo_130 = _GEN_523;
  wire [63:0]      _GEN_524 = {dataRegroupBySew_3_2_11, dataRegroupBySew_2_2_11};
  wire [63:0]      dataInMem_hi_622;
  assign dataInMem_hi_622 = _GEN_524;
  wire [63:0]      dataInMem_lo_hi_354;
  assign dataInMem_lo_hi_354 = _GEN_524;
  wire [63:0]      _GEN_525 = {dataRegroupBySew_1_2_12, dataRegroupBySew_0_2_12};
  wire [63:0]      dataInMem_lo_511;
  assign dataInMem_lo_511 = _GEN_525;
  wire [63:0]      dataInMem_lo_528;
  assign dataInMem_lo_528 = _GEN_525;
  wire [63:0]      dataInMem_lo_lo_131;
  assign dataInMem_lo_lo_131 = _GEN_525;
  wire [63:0]      _GEN_526 = {dataRegroupBySew_3_2_12, dataRegroupBySew_2_2_12};
  wire [63:0]      dataInMem_hi_623;
  assign dataInMem_hi_623 = _GEN_526;
  wire [63:0]      dataInMem_lo_hi_355;
  assign dataInMem_lo_hi_355 = _GEN_526;
  wire [63:0]      _GEN_527 = {dataRegroupBySew_1_2_13, dataRegroupBySew_0_2_13};
  wire [63:0]      dataInMem_lo_512;
  assign dataInMem_lo_512 = _GEN_527;
  wire [63:0]      dataInMem_lo_529;
  assign dataInMem_lo_529 = _GEN_527;
  wire [63:0]      dataInMem_lo_lo_132;
  assign dataInMem_lo_lo_132 = _GEN_527;
  wire [63:0]      _GEN_528 = {dataRegroupBySew_3_2_13, dataRegroupBySew_2_2_13};
  wire [63:0]      dataInMem_hi_624;
  assign dataInMem_hi_624 = _GEN_528;
  wire [63:0]      dataInMem_lo_hi_356;
  assign dataInMem_lo_hi_356 = _GEN_528;
  wire [63:0]      _GEN_529 = {dataRegroupBySew_1_2_14, dataRegroupBySew_0_2_14};
  wire [63:0]      dataInMem_lo_513;
  assign dataInMem_lo_513 = _GEN_529;
  wire [63:0]      dataInMem_lo_530;
  assign dataInMem_lo_530 = _GEN_529;
  wire [63:0]      dataInMem_lo_lo_133;
  assign dataInMem_lo_lo_133 = _GEN_529;
  wire [63:0]      _GEN_530 = {dataRegroupBySew_3_2_14, dataRegroupBySew_2_2_14};
  wire [63:0]      dataInMem_hi_625;
  assign dataInMem_hi_625 = _GEN_530;
  wire [63:0]      dataInMem_lo_hi_357;
  assign dataInMem_lo_hi_357 = _GEN_530;
  wire [63:0]      _GEN_531 = {dataRegroupBySew_1_2_15, dataRegroupBySew_0_2_15};
  wire [63:0]      dataInMem_lo_514;
  assign dataInMem_lo_514 = _GEN_531;
  wire [63:0]      dataInMem_lo_531;
  assign dataInMem_lo_531 = _GEN_531;
  wire [63:0]      dataInMem_lo_lo_134;
  assign dataInMem_lo_lo_134 = _GEN_531;
  wire [63:0]      _GEN_532 = {dataRegroupBySew_3_2_15, dataRegroupBySew_2_2_15};
  wire [63:0]      dataInMem_hi_626;
  assign dataInMem_hi_626 = _GEN_532;
  wire [63:0]      dataInMem_lo_hi_358;
  assign dataInMem_lo_hi_358 = _GEN_532;
  wire [255:0]     dataInMem_lo_lo_lo_19 = {dataInMem_hi_612, dataInMem_lo_500, dataInMem_hi_611, dataInMem_lo_499};
  wire [255:0]     dataInMem_lo_lo_hi_19 = {dataInMem_hi_614, dataInMem_lo_502, dataInMem_hi_613, dataInMem_lo_501};
  wire [511:0]     dataInMem_lo_lo_115 = {dataInMem_lo_lo_hi_19, dataInMem_lo_lo_lo_19};
  wire [255:0]     dataInMem_lo_hi_lo_19 = {dataInMem_hi_616, dataInMem_lo_504, dataInMem_hi_615, dataInMem_lo_503};
  wire [255:0]     dataInMem_lo_hi_hi_19 = {dataInMem_hi_618, dataInMem_lo_506, dataInMem_hi_617, dataInMem_lo_505};
  wire [511:0]     dataInMem_lo_hi_307 = {dataInMem_lo_hi_hi_19, dataInMem_lo_hi_lo_19};
  wire [1023:0]    dataInMem_lo_515 = {dataInMem_lo_hi_307, dataInMem_lo_lo_115};
  wire [255:0]     dataInMem_hi_lo_lo_19 = {dataInMem_hi_620, dataInMem_lo_508, dataInMem_hi_619, dataInMem_lo_507};
  wire [255:0]     dataInMem_hi_lo_hi_19 = {dataInMem_hi_622, dataInMem_lo_510, dataInMem_hi_621, dataInMem_lo_509};
  wire [511:0]     dataInMem_hi_lo_211 = {dataInMem_hi_lo_hi_19, dataInMem_hi_lo_lo_19};
  wire [255:0]     dataInMem_hi_hi_lo_19 = {dataInMem_hi_624, dataInMem_lo_512, dataInMem_hi_623, dataInMem_lo_511};
  wire [255:0]     dataInMem_hi_hi_hi_19 = {dataInMem_hi_626, dataInMem_lo_514, dataInMem_hi_625, dataInMem_lo_513};
  wire [511:0]     dataInMem_hi_hi_403 = {dataInMem_hi_hi_hi_19, dataInMem_hi_hi_lo_19};
  wire [1023:0]    dataInMem_hi_627 = {dataInMem_hi_hi_403, dataInMem_hi_lo_211};
  wire [2047:0]    dataInMem_19 = {dataInMem_hi_627, dataInMem_lo_515};
  wire [511:0]     regroupCacheLine_19_0 = dataInMem_19[511:0];
  wire [511:0]     regroupCacheLine_19_1 = dataInMem_19[1023:512];
  wire [511:0]     regroupCacheLine_19_2 = dataInMem_19[1535:1024];
  wire [511:0]     regroupCacheLine_19_3 = dataInMem_19[2047:1536];
  wire [511:0]     res_152 = regroupCacheLine_19_0;
  wire [511:0]     res_153 = regroupCacheLine_19_1;
  wire [511:0]     res_154 = regroupCacheLine_19_2;
  wire [511:0]     res_155 = regroupCacheLine_19_3;
  wire [1023:0]    lo_lo_19 = {res_153, res_152};
  wire [1023:0]    lo_hi_19 = {res_155, res_154};
  wire [2047:0]    lo_19 = {lo_hi_19, lo_lo_19};
  wire [4095:0]    regroupLoadData_2_3 = {2048'h0, lo_19};
  wire [63:0]      _GEN_533 = {dataRegroupBySew_4_2_0, dataRegroupBySew_3_2_0};
  wire [63:0]      dataInMem_hi_hi_404;
  assign dataInMem_hi_hi_404 = _GEN_533;
  wire [63:0]      dataInMem_hi_lo_214;
  assign dataInMem_hi_lo_214 = _GEN_533;
  wire [95:0]      dataInMem_hi_628 = {dataInMem_hi_hi_404, dataRegroupBySew_2_2_0};
  wire [63:0]      _GEN_534 = {dataRegroupBySew_4_2_1, dataRegroupBySew_3_2_1};
  wire [63:0]      dataInMem_hi_hi_405;
  assign dataInMem_hi_hi_405 = _GEN_534;
  wire [63:0]      dataInMem_hi_lo_215;
  assign dataInMem_hi_lo_215 = _GEN_534;
  wire [95:0]      dataInMem_hi_629 = {dataInMem_hi_hi_405, dataRegroupBySew_2_2_1};
  wire [63:0]      _GEN_535 = {dataRegroupBySew_4_2_2, dataRegroupBySew_3_2_2};
  wire [63:0]      dataInMem_hi_hi_406;
  assign dataInMem_hi_hi_406 = _GEN_535;
  wire [63:0]      dataInMem_hi_lo_216;
  assign dataInMem_hi_lo_216 = _GEN_535;
  wire [95:0]      dataInMem_hi_630 = {dataInMem_hi_hi_406, dataRegroupBySew_2_2_2};
  wire [63:0]      _GEN_536 = {dataRegroupBySew_4_2_3, dataRegroupBySew_3_2_3};
  wire [63:0]      dataInMem_hi_hi_407;
  assign dataInMem_hi_hi_407 = _GEN_536;
  wire [63:0]      dataInMem_hi_lo_217;
  assign dataInMem_hi_lo_217 = _GEN_536;
  wire [95:0]      dataInMem_hi_631 = {dataInMem_hi_hi_407, dataRegroupBySew_2_2_3};
  wire [63:0]      _GEN_537 = {dataRegroupBySew_4_2_4, dataRegroupBySew_3_2_4};
  wire [63:0]      dataInMem_hi_hi_408;
  assign dataInMem_hi_hi_408 = _GEN_537;
  wire [63:0]      dataInMem_hi_lo_218;
  assign dataInMem_hi_lo_218 = _GEN_537;
  wire [95:0]      dataInMem_hi_632 = {dataInMem_hi_hi_408, dataRegroupBySew_2_2_4};
  wire [63:0]      _GEN_538 = {dataRegroupBySew_4_2_5, dataRegroupBySew_3_2_5};
  wire [63:0]      dataInMem_hi_hi_409;
  assign dataInMem_hi_hi_409 = _GEN_538;
  wire [63:0]      dataInMem_hi_lo_219;
  assign dataInMem_hi_lo_219 = _GEN_538;
  wire [95:0]      dataInMem_hi_633 = {dataInMem_hi_hi_409, dataRegroupBySew_2_2_5};
  wire [63:0]      _GEN_539 = {dataRegroupBySew_4_2_6, dataRegroupBySew_3_2_6};
  wire [63:0]      dataInMem_hi_hi_410;
  assign dataInMem_hi_hi_410 = _GEN_539;
  wire [63:0]      dataInMem_hi_lo_220;
  assign dataInMem_hi_lo_220 = _GEN_539;
  wire [95:0]      dataInMem_hi_634 = {dataInMem_hi_hi_410, dataRegroupBySew_2_2_6};
  wire [63:0]      _GEN_540 = {dataRegroupBySew_4_2_7, dataRegroupBySew_3_2_7};
  wire [63:0]      dataInMem_hi_hi_411;
  assign dataInMem_hi_hi_411 = _GEN_540;
  wire [63:0]      dataInMem_hi_lo_221;
  assign dataInMem_hi_lo_221 = _GEN_540;
  wire [95:0]      dataInMem_hi_635 = {dataInMem_hi_hi_411, dataRegroupBySew_2_2_7};
  wire [63:0]      _GEN_541 = {dataRegroupBySew_4_2_8, dataRegroupBySew_3_2_8};
  wire [63:0]      dataInMem_hi_hi_412;
  assign dataInMem_hi_hi_412 = _GEN_541;
  wire [63:0]      dataInMem_hi_lo_222;
  assign dataInMem_hi_lo_222 = _GEN_541;
  wire [95:0]      dataInMem_hi_636 = {dataInMem_hi_hi_412, dataRegroupBySew_2_2_8};
  wire [63:0]      _GEN_542 = {dataRegroupBySew_4_2_9, dataRegroupBySew_3_2_9};
  wire [63:0]      dataInMem_hi_hi_413;
  assign dataInMem_hi_hi_413 = _GEN_542;
  wire [63:0]      dataInMem_hi_lo_223;
  assign dataInMem_hi_lo_223 = _GEN_542;
  wire [95:0]      dataInMem_hi_637 = {dataInMem_hi_hi_413, dataRegroupBySew_2_2_9};
  wire [63:0]      _GEN_543 = {dataRegroupBySew_4_2_10, dataRegroupBySew_3_2_10};
  wire [63:0]      dataInMem_hi_hi_414;
  assign dataInMem_hi_hi_414 = _GEN_543;
  wire [63:0]      dataInMem_hi_lo_224;
  assign dataInMem_hi_lo_224 = _GEN_543;
  wire [95:0]      dataInMem_hi_638 = {dataInMem_hi_hi_414, dataRegroupBySew_2_2_10};
  wire [63:0]      _GEN_544 = {dataRegroupBySew_4_2_11, dataRegroupBySew_3_2_11};
  wire [63:0]      dataInMem_hi_hi_415;
  assign dataInMem_hi_hi_415 = _GEN_544;
  wire [63:0]      dataInMem_hi_lo_225;
  assign dataInMem_hi_lo_225 = _GEN_544;
  wire [95:0]      dataInMem_hi_639 = {dataInMem_hi_hi_415, dataRegroupBySew_2_2_11};
  wire [63:0]      _GEN_545 = {dataRegroupBySew_4_2_12, dataRegroupBySew_3_2_12};
  wire [63:0]      dataInMem_hi_hi_416;
  assign dataInMem_hi_hi_416 = _GEN_545;
  wire [63:0]      dataInMem_hi_lo_226;
  assign dataInMem_hi_lo_226 = _GEN_545;
  wire [95:0]      dataInMem_hi_640 = {dataInMem_hi_hi_416, dataRegroupBySew_2_2_12};
  wire [63:0]      _GEN_546 = {dataRegroupBySew_4_2_13, dataRegroupBySew_3_2_13};
  wire [63:0]      dataInMem_hi_hi_417;
  assign dataInMem_hi_hi_417 = _GEN_546;
  wire [63:0]      dataInMem_hi_lo_227;
  assign dataInMem_hi_lo_227 = _GEN_546;
  wire [95:0]      dataInMem_hi_641 = {dataInMem_hi_hi_417, dataRegroupBySew_2_2_13};
  wire [63:0]      _GEN_547 = {dataRegroupBySew_4_2_14, dataRegroupBySew_3_2_14};
  wire [63:0]      dataInMem_hi_hi_418;
  assign dataInMem_hi_hi_418 = _GEN_547;
  wire [63:0]      dataInMem_hi_lo_228;
  assign dataInMem_hi_lo_228 = _GEN_547;
  wire [95:0]      dataInMem_hi_642 = {dataInMem_hi_hi_418, dataRegroupBySew_2_2_14};
  wire [63:0]      _GEN_548 = {dataRegroupBySew_4_2_15, dataRegroupBySew_3_2_15};
  wire [63:0]      dataInMem_hi_hi_419;
  assign dataInMem_hi_hi_419 = _GEN_548;
  wire [63:0]      dataInMem_hi_lo_229;
  assign dataInMem_hi_lo_229 = _GEN_548;
  wire [95:0]      dataInMem_hi_643 = {dataInMem_hi_hi_419, dataRegroupBySew_2_2_15};
  wire [319:0]     dataInMem_lo_lo_lo_20 = {dataInMem_hi_629, dataInMem_lo_517, dataInMem_hi_628, dataInMem_lo_516};
  wire [319:0]     dataInMem_lo_lo_hi_20 = {dataInMem_hi_631, dataInMem_lo_519, dataInMem_hi_630, dataInMem_lo_518};
  wire [639:0]     dataInMem_lo_lo_116 = {dataInMem_lo_lo_hi_20, dataInMem_lo_lo_lo_20};
  wire [319:0]     dataInMem_lo_hi_lo_20 = {dataInMem_hi_633, dataInMem_lo_521, dataInMem_hi_632, dataInMem_lo_520};
  wire [319:0]     dataInMem_lo_hi_hi_20 = {dataInMem_hi_635, dataInMem_lo_523, dataInMem_hi_634, dataInMem_lo_522};
  wire [639:0]     dataInMem_lo_hi_308 = {dataInMem_lo_hi_hi_20, dataInMem_lo_hi_lo_20};
  wire [1279:0]    dataInMem_lo_532 = {dataInMem_lo_hi_308, dataInMem_lo_lo_116};
  wire [319:0]     dataInMem_hi_lo_lo_20 = {dataInMem_hi_637, dataInMem_lo_525, dataInMem_hi_636, dataInMem_lo_524};
  wire [319:0]     dataInMem_hi_lo_hi_20 = {dataInMem_hi_639, dataInMem_lo_527, dataInMem_hi_638, dataInMem_lo_526};
  wire [639:0]     dataInMem_hi_lo_212 = {dataInMem_hi_lo_hi_20, dataInMem_hi_lo_lo_20};
  wire [319:0]     dataInMem_hi_hi_lo_20 = {dataInMem_hi_641, dataInMem_lo_529, dataInMem_hi_640, dataInMem_lo_528};
  wire [319:0]     dataInMem_hi_hi_hi_20 = {dataInMem_hi_643, dataInMem_lo_531, dataInMem_hi_642, dataInMem_lo_530};
  wire [639:0]     dataInMem_hi_hi_420 = {dataInMem_hi_hi_hi_20, dataInMem_hi_hi_lo_20};
  wire [1279:0]    dataInMem_hi_644 = {dataInMem_hi_hi_420, dataInMem_hi_lo_212};
  wire [2559:0]    dataInMem_20 = {dataInMem_hi_644, dataInMem_lo_532};
  wire [511:0]     regroupCacheLine_20_0 = dataInMem_20[511:0];
  wire [511:0]     regroupCacheLine_20_1 = dataInMem_20[1023:512];
  wire [511:0]     regroupCacheLine_20_2 = dataInMem_20[1535:1024];
  wire [511:0]     regroupCacheLine_20_3 = dataInMem_20[2047:1536];
  wire [511:0]     regroupCacheLine_20_4 = dataInMem_20[2559:2048];
  wire [511:0]     res_160 = regroupCacheLine_20_0;
  wire [511:0]     res_161 = regroupCacheLine_20_1;
  wire [511:0]     res_162 = regroupCacheLine_20_2;
  wire [511:0]     res_163 = regroupCacheLine_20_3;
  wire [511:0]     res_164 = regroupCacheLine_20_4;
  wire [1023:0]    lo_lo_20 = {res_161, res_160};
  wire [1023:0]    lo_hi_20 = {res_163, res_162};
  wire [2047:0]    lo_20 = {lo_hi_20, lo_lo_20};
  wire [1023:0]    hi_lo_20 = {512'h0, res_164};
  wire [2047:0]    hi_20 = {1024'h0, hi_lo_20};
  wire [4095:0]    regroupLoadData_2_4 = {hi_20, lo_20};
  wire [95:0]      dataInMem_lo_533 = {dataInMem_lo_hi_309, dataRegroupBySew_0_2_0};
  wire [63:0]      _GEN_549 = {dataRegroupBySew_5_2_0, dataRegroupBySew_4_2_0};
  wire [63:0]      dataInMem_hi_hi_421;
  assign dataInMem_hi_hi_421 = _GEN_549;
  wire [63:0]      dataInMem_hi_lo_231;
  assign dataInMem_hi_lo_231 = _GEN_549;
  wire [95:0]      dataInMem_hi_645 = {dataInMem_hi_hi_421, dataRegroupBySew_3_2_0};
  wire [95:0]      dataInMem_lo_534 = {dataInMem_lo_hi_310, dataRegroupBySew_0_2_1};
  wire [63:0]      _GEN_550 = {dataRegroupBySew_5_2_1, dataRegroupBySew_4_2_1};
  wire [63:0]      dataInMem_hi_hi_422;
  assign dataInMem_hi_hi_422 = _GEN_550;
  wire [63:0]      dataInMem_hi_lo_232;
  assign dataInMem_hi_lo_232 = _GEN_550;
  wire [95:0]      dataInMem_hi_646 = {dataInMem_hi_hi_422, dataRegroupBySew_3_2_1};
  wire [95:0]      dataInMem_lo_535 = {dataInMem_lo_hi_311, dataRegroupBySew_0_2_2};
  wire [63:0]      _GEN_551 = {dataRegroupBySew_5_2_2, dataRegroupBySew_4_2_2};
  wire [63:0]      dataInMem_hi_hi_423;
  assign dataInMem_hi_hi_423 = _GEN_551;
  wire [63:0]      dataInMem_hi_lo_233;
  assign dataInMem_hi_lo_233 = _GEN_551;
  wire [95:0]      dataInMem_hi_647 = {dataInMem_hi_hi_423, dataRegroupBySew_3_2_2};
  wire [95:0]      dataInMem_lo_536 = {dataInMem_lo_hi_312, dataRegroupBySew_0_2_3};
  wire [63:0]      _GEN_552 = {dataRegroupBySew_5_2_3, dataRegroupBySew_4_2_3};
  wire [63:0]      dataInMem_hi_hi_424;
  assign dataInMem_hi_hi_424 = _GEN_552;
  wire [63:0]      dataInMem_hi_lo_234;
  assign dataInMem_hi_lo_234 = _GEN_552;
  wire [95:0]      dataInMem_hi_648 = {dataInMem_hi_hi_424, dataRegroupBySew_3_2_3};
  wire [95:0]      dataInMem_lo_537 = {dataInMem_lo_hi_313, dataRegroupBySew_0_2_4};
  wire [63:0]      _GEN_553 = {dataRegroupBySew_5_2_4, dataRegroupBySew_4_2_4};
  wire [63:0]      dataInMem_hi_hi_425;
  assign dataInMem_hi_hi_425 = _GEN_553;
  wire [63:0]      dataInMem_hi_lo_235;
  assign dataInMem_hi_lo_235 = _GEN_553;
  wire [95:0]      dataInMem_hi_649 = {dataInMem_hi_hi_425, dataRegroupBySew_3_2_4};
  wire [95:0]      dataInMem_lo_538 = {dataInMem_lo_hi_314, dataRegroupBySew_0_2_5};
  wire [63:0]      _GEN_554 = {dataRegroupBySew_5_2_5, dataRegroupBySew_4_2_5};
  wire [63:0]      dataInMem_hi_hi_426;
  assign dataInMem_hi_hi_426 = _GEN_554;
  wire [63:0]      dataInMem_hi_lo_236;
  assign dataInMem_hi_lo_236 = _GEN_554;
  wire [95:0]      dataInMem_hi_650 = {dataInMem_hi_hi_426, dataRegroupBySew_3_2_5};
  wire [95:0]      dataInMem_lo_539 = {dataInMem_lo_hi_315, dataRegroupBySew_0_2_6};
  wire [63:0]      _GEN_555 = {dataRegroupBySew_5_2_6, dataRegroupBySew_4_2_6};
  wire [63:0]      dataInMem_hi_hi_427;
  assign dataInMem_hi_hi_427 = _GEN_555;
  wire [63:0]      dataInMem_hi_lo_237;
  assign dataInMem_hi_lo_237 = _GEN_555;
  wire [95:0]      dataInMem_hi_651 = {dataInMem_hi_hi_427, dataRegroupBySew_3_2_6};
  wire [95:0]      dataInMem_lo_540 = {dataInMem_lo_hi_316, dataRegroupBySew_0_2_7};
  wire [63:0]      _GEN_556 = {dataRegroupBySew_5_2_7, dataRegroupBySew_4_2_7};
  wire [63:0]      dataInMem_hi_hi_428;
  assign dataInMem_hi_hi_428 = _GEN_556;
  wire [63:0]      dataInMem_hi_lo_238;
  assign dataInMem_hi_lo_238 = _GEN_556;
  wire [95:0]      dataInMem_hi_652 = {dataInMem_hi_hi_428, dataRegroupBySew_3_2_7};
  wire [95:0]      dataInMem_lo_541 = {dataInMem_lo_hi_317, dataRegroupBySew_0_2_8};
  wire [63:0]      _GEN_557 = {dataRegroupBySew_5_2_8, dataRegroupBySew_4_2_8};
  wire [63:0]      dataInMem_hi_hi_429;
  assign dataInMem_hi_hi_429 = _GEN_557;
  wire [63:0]      dataInMem_hi_lo_239;
  assign dataInMem_hi_lo_239 = _GEN_557;
  wire [95:0]      dataInMem_hi_653 = {dataInMem_hi_hi_429, dataRegroupBySew_3_2_8};
  wire [95:0]      dataInMem_lo_542 = {dataInMem_lo_hi_318, dataRegroupBySew_0_2_9};
  wire [63:0]      _GEN_558 = {dataRegroupBySew_5_2_9, dataRegroupBySew_4_2_9};
  wire [63:0]      dataInMem_hi_hi_430;
  assign dataInMem_hi_hi_430 = _GEN_558;
  wire [63:0]      dataInMem_hi_lo_240;
  assign dataInMem_hi_lo_240 = _GEN_558;
  wire [95:0]      dataInMem_hi_654 = {dataInMem_hi_hi_430, dataRegroupBySew_3_2_9};
  wire [95:0]      dataInMem_lo_543 = {dataInMem_lo_hi_319, dataRegroupBySew_0_2_10};
  wire [63:0]      _GEN_559 = {dataRegroupBySew_5_2_10, dataRegroupBySew_4_2_10};
  wire [63:0]      dataInMem_hi_hi_431;
  assign dataInMem_hi_hi_431 = _GEN_559;
  wire [63:0]      dataInMem_hi_lo_241;
  assign dataInMem_hi_lo_241 = _GEN_559;
  wire [95:0]      dataInMem_hi_655 = {dataInMem_hi_hi_431, dataRegroupBySew_3_2_10};
  wire [95:0]      dataInMem_lo_544 = {dataInMem_lo_hi_320, dataRegroupBySew_0_2_11};
  wire [63:0]      _GEN_560 = {dataRegroupBySew_5_2_11, dataRegroupBySew_4_2_11};
  wire [63:0]      dataInMem_hi_hi_432;
  assign dataInMem_hi_hi_432 = _GEN_560;
  wire [63:0]      dataInMem_hi_lo_242;
  assign dataInMem_hi_lo_242 = _GEN_560;
  wire [95:0]      dataInMem_hi_656 = {dataInMem_hi_hi_432, dataRegroupBySew_3_2_11};
  wire [95:0]      dataInMem_lo_545 = {dataInMem_lo_hi_321, dataRegroupBySew_0_2_12};
  wire [63:0]      _GEN_561 = {dataRegroupBySew_5_2_12, dataRegroupBySew_4_2_12};
  wire [63:0]      dataInMem_hi_hi_433;
  assign dataInMem_hi_hi_433 = _GEN_561;
  wire [63:0]      dataInMem_hi_lo_243;
  assign dataInMem_hi_lo_243 = _GEN_561;
  wire [95:0]      dataInMem_hi_657 = {dataInMem_hi_hi_433, dataRegroupBySew_3_2_12};
  wire [95:0]      dataInMem_lo_546 = {dataInMem_lo_hi_322, dataRegroupBySew_0_2_13};
  wire [63:0]      _GEN_562 = {dataRegroupBySew_5_2_13, dataRegroupBySew_4_2_13};
  wire [63:0]      dataInMem_hi_hi_434;
  assign dataInMem_hi_hi_434 = _GEN_562;
  wire [63:0]      dataInMem_hi_lo_244;
  assign dataInMem_hi_lo_244 = _GEN_562;
  wire [95:0]      dataInMem_hi_658 = {dataInMem_hi_hi_434, dataRegroupBySew_3_2_13};
  wire [95:0]      dataInMem_lo_547 = {dataInMem_lo_hi_323, dataRegroupBySew_0_2_14};
  wire [63:0]      _GEN_563 = {dataRegroupBySew_5_2_14, dataRegroupBySew_4_2_14};
  wire [63:0]      dataInMem_hi_hi_435;
  assign dataInMem_hi_hi_435 = _GEN_563;
  wire [63:0]      dataInMem_hi_lo_245;
  assign dataInMem_hi_lo_245 = _GEN_563;
  wire [95:0]      dataInMem_hi_659 = {dataInMem_hi_hi_435, dataRegroupBySew_3_2_14};
  wire [95:0]      dataInMem_lo_548 = {dataInMem_lo_hi_324, dataRegroupBySew_0_2_15};
  wire [63:0]      _GEN_564 = {dataRegroupBySew_5_2_15, dataRegroupBySew_4_2_15};
  wire [63:0]      dataInMem_hi_hi_436;
  assign dataInMem_hi_hi_436 = _GEN_564;
  wire [63:0]      dataInMem_hi_lo_246;
  assign dataInMem_hi_lo_246 = _GEN_564;
  wire [95:0]      dataInMem_hi_660 = {dataInMem_hi_hi_436, dataRegroupBySew_3_2_15};
  wire [383:0]     dataInMem_lo_lo_lo_21 = {dataInMem_hi_646, dataInMem_lo_534, dataInMem_hi_645, dataInMem_lo_533};
  wire [383:0]     dataInMem_lo_lo_hi_21 = {dataInMem_hi_648, dataInMem_lo_536, dataInMem_hi_647, dataInMem_lo_535};
  wire [767:0]     dataInMem_lo_lo_117 = {dataInMem_lo_lo_hi_21, dataInMem_lo_lo_lo_21};
  wire [383:0]     dataInMem_lo_hi_lo_21 = {dataInMem_hi_650, dataInMem_lo_538, dataInMem_hi_649, dataInMem_lo_537};
  wire [383:0]     dataInMem_lo_hi_hi_21 = {dataInMem_hi_652, dataInMem_lo_540, dataInMem_hi_651, dataInMem_lo_539};
  wire [767:0]     dataInMem_lo_hi_325 = {dataInMem_lo_hi_hi_21, dataInMem_lo_hi_lo_21};
  wire [1535:0]    dataInMem_lo_549 = {dataInMem_lo_hi_325, dataInMem_lo_lo_117};
  wire [383:0]     dataInMem_hi_lo_lo_21 = {dataInMem_hi_654, dataInMem_lo_542, dataInMem_hi_653, dataInMem_lo_541};
  wire [383:0]     dataInMem_hi_lo_hi_21 = {dataInMem_hi_656, dataInMem_lo_544, dataInMem_hi_655, dataInMem_lo_543};
  wire [767:0]     dataInMem_hi_lo_213 = {dataInMem_hi_lo_hi_21, dataInMem_hi_lo_lo_21};
  wire [383:0]     dataInMem_hi_hi_lo_21 = {dataInMem_hi_658, dataInMem_lo_546, dataInMem_hi_657, dataInMem_lo_545};
  wire [383:0]     dataInMem_hi_hi_hi_21 = {dataInMem_hi_660, dataInMem_lo_548, dataInMem_hi_659, dataInMem_lo_547};
  wire [767:0]     dataInMem_hi_hi_437 = {dataInMem_hi_hi_hi_21, dataInMem_hi_hi_lo_21};
  wire [1535:0]    dataInMem_hi_661 = {dataInMem_hi_hi_437, dataInMem_hi_lo_213};
  wire [3071:0]    dataInMem_21 = {dataInMem_hi_661, dataInMem_lo_549};
  wire [511:0]     regroupCacheLine_21_0 = dataInMem_21[511:0];
  wire [511:0]     regroupCacheLine_21_1 = dataInMem_21[1023:512];
  wire [511:0]     regroupCacheLine_21_2 = dataInMem_21[1535:1024];
  wire [511:0]     regroupCacheLine_21_3 = dataInMem_21[2047:1536];
  wire [511:0]     regroupCacheLine_21_4 = dataInMem_21[2559:2048];
  wire [511:0]     regroupCacheLine_21_5 = dataInMem_21[3071:2560];
  wire [511:0]     res_168 = regroupCacheLine_21_0;
  wire [511:0]     res_169 = regroupCacheLine_21_1;
  wire [511:0]     res_170 = regroupCacheLine_21_2;
  wire [511:0]     res_171 = regroupCacheLine_21_3;
  wire [511:0]     res_172 = regroupCacheLine_21_4;
  wire [511:0]     res_173 = regroupCacheLine_21_5;
  wire [1023:0]    lo_lo_21 = {res_169, res_168};
  wire [1023:0]    lo_hi_21 = {res_171, res_170};
  wire [2047:0]    lo_21 = {lo_hi_21, lo_lo_21};
  wire [1023:0]    hi_lo_21 = {res_173, res_172};
  wire [2047:0]    hi_21 = {1024'h0, hi_lo_21};
  wire [4095:0]    regroupLoadData_2_5 = {hi_21, lo_21};
  wire [95:0]      dataInMem_lo_550 = {dataInMem_lo_hi_326, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_hi_hi_438 = {dataRegroupBySew_6_2_0, dataRegroupBySew_5_2_0};
  wire [127:0]     dataInMem_hi_662 = {dataInMem_hi_hi_438, dataInMem_hi_lo_214};
  wire [95:0]      dataInMem_lo_551 = {dataInMem_lo_hi_327, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_hi_hi_439 = {dataRegroupBySew_6_2_1, dataRegroupBySew_5_2_1};
  wire [127:0]     dataInMem_hi_663 = {dataInMem_hi_hi_439, dataInMem_hi_lo_215};
  wire [95:0]      dataInMem_lo_552 = {dataInMem_lo_hi_328, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_hi_hi_440 = {dataRegroupBySew_6_2_2, dataRegroupBySew_5_2_2};
  wire [127:0]     dataInMem_hi_664 = {dataInMem_hi_hi_440, dataInMem_hi_lo_216};
  wire [95:0]      dataInMem_lo_553 = {dataInMem_lo_hi_329, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_hi_hi_441 = {dataRegroupBySew_6_2_3, dataRegroupBySew_5_2_3};
  wire [127:0]     dataInMem_hi_665 = {dataInMem_hi_hi_441, dataInMem_hi_lo_217};
  wire [95:0]      dataInMem_lo_554 = {dataInMem_lo_hi_330, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_hi_hi_442 = {dataRegroupBySew_6_2_4, dataRegroupBySew_5_2_4};
  wire [127:0]     dataInMem_hi_666 = {dataInMem_hi_hi_442, dataInMem_hi_lo_218};
  wire [95:0]      dataInMem_lo_555 = {dataInMem_lo_hi_331, dataRegroupBySew_0_2_5};
  wire [63:0]      dataInMem_hi_hi_443 = {dataRegroupBySew_6_2_5, dataRegroupBySew_5_2_5};
  wire [127:0]     dataInMem_hi_667 = {dataInMem_hi_hi_443, dataInMem_hi_lo_219};
  wire [95:0]      dataInMem_lo_556 = {dataInMem_lo_hi_332, dataRegroupBySew_0_2_6};
  wire [63:0]      dataInMem_hi_hi_444 = {dataRegroupBySew_6_2_6, dataRegroupBySew_5_2_6};
  wire [127:0]     dataInMem_hi_668 = {dataInMem_hi_hi_444, dataInMem_hi_lo_220};
  wire [95:0]      dataInMem_lo_557 = {dataInMem_lo_hi_333, dataRegroupBySew_0_2_7};
  wire [63:0]      dataInMem_hi_hi_445 = {dataRegroupBySew_6_2_7, dataRegroupBySew_5_2_7};
  wire [127:0]     dataInMem_hi_669 = {dataInMem_hi_hi_445, dataInMem_hi_lo_221};
  wire [95:0]      dataInMem_lo_558 = {dataInMem_lo_hi_334, dataRegroupBySew_0_2_8};
  wire [63:0]      dataInMem_hi_hi_446 = {dataRegroupBySew_6_2_8, dataRegroupBySew_5_2_8};
  wire [127:0]     dataInMem_hi_670 = {dataInMem_hi_hi_446, dataInMem_hi_lo_222};
  wire [95:0]      dataInMem_lo_559 = {dataInMem_lo_hi_335, dataRegroupBySew_0_2_9};
  wire [63:0]      dataInMem_hi_hi_447 = {dataRegroupBySew_6_2_9, dataRegroupBySew_5_2_9};
  wire [127:0]     dataInMem_hi_671 = {dataInMem_hi_hi_447, dataInMem_hi_lo_223};
  wire [95:0]      dataInMem_lo_560 = {dataInMem_lo_hi_336, dataRegroupBySew_0_2_10};
  wire [63:0]      dataInMem_hi_hi_448 = {dataRegroupBySew_6_2_10, dataRegroupBySew_5_2_10};
  wire [127:0]     dataInMem_hi_672 = {dataInMem_hi_hi_448, dataInMem_hi_lo_224};
  wire [95:0]      dataInMem_lo_561 = {dataInMem_lo_hi_337, dataRegroupBySew_0_2_11};
  wire [63:0]      dataInMem_hi_hi_449 = {dataRegroupBySew_6_2_11, dataRegroupBySew_5_2_11};
  wire [127:0]     dataInMem_hi_673 = {dataInMem_hi_hi_449, dataInMem_hi_lo_225};
  wire [95:0]      dataInMem_lo_562 = {dataInMem_lo_hi_338, dataRegroupBySew_0_2_12};
  wire [63:0]      dataInMem_hi_hi_450 = {dataRegroupBySew_6_2_12, dataRegroupBySew_5_2_12};
  wire [127:0]     dataInMem_hi_674 = {dataInMem_hi_hi_450, dataInMem_hi_lo_226};
  wire [95:0]      dataInMem_lo_563 = {dataInMem_lo_hi_339, dataRegroupBySew_0_2_13};
  wire [63:0]      dataInMem_hi_hi_451 = {dataRegroupBySew_6_2_13, dataRegroupBySew_5_2_13};
  wire [127:0]     dataInMem_hi_675 = {dataInMem_hi_hi_451, dataInMem_hi_lo_227};
  wire [95:0]      dataInMem_lo_564 = {dataInMem_lo_hi_340, dataRegroupBySew_0_2_14};
  wire [63:0]      dataInMem_hi_hi_452 = {dataRegroupBySew_6_2_14, dataRegroupBySew_5_2_14};
  wire [127:0]     dataInMem_hi_676 = {dataInMem_hi_hi_452, dataInMem_hi_lo_228};
  wire [95:0]      dataInMem_lo_565 = {dataInMem_lo_hi_341, dataRegroupBySew_0_2_15};
  wire [63:0]      dataInMem_hi_hi_453 = {dataRegroupBySew_6_2_15, dataRegroupBySew_5_2_15};
  wire [127:0]     dataInMem_hi_677 = {dataInMem_hi_hi_453, dataInMem_hi_lo_229};
  wire [447:0]     dataInMem_lo_lo_lo_22 = {dataInMem_hi_663, dataInMem_lo_551, dataInMem_hi_662, dataInMem_lo_550};
  wire [447:0]     dataInMem_lo_lo_hi_22 = {dataInMem_hi_665, dataInMem_lo_553, dataInMem_hi_664, dataInMem_lo_552};
  wire [895:0]     dataInMem_lo_lo_118 = {dataInMem_lo_lo_hi_22, dataInMem_lo_lo_lo_22};
  wire [447:0]     dataInMem_lo_hi_lo_22 = {dataInMem_hi_667, dataInMem_lo_555, dataInMem_hi_666, dataInMem_lo_554};
  wire [447:0]     dataInMem_lo_hi_hi_22 = {dataInMem_hi_669, dataInMem_lo_557, dataInMem_hi_668, dataInMem_lo_556};
  wire [895:0]     dataInMem_lo_hi_342 = {dataInMem_lo_hi_hi_22, dataInMem_lo_hi_lo_22};
  wire [1791:0]    dataInMem_lo_566 = {dataInMem_lo_hi_342, dataInMem_lo_lo_118};
  wire [447:0]     dataInMem_hi_lo_lo_22 = {dataInMem_hi_671, dataInMem_lo_559, dataInMem_hi_670, dataInMem_lo_558};
  wire [447:0]     dataInMem_hi_lo_hi_22 = {dataInMem_hi_673, dataInMem_lo_561, dataInMem_hi_672, dataInMem_lo_560};
  wire [895:0]     dataInMem_hi_lo_230 = {dataInMem_hi_lo_hi_22, dataInMem_hi_lo_lo_22};
  wire [447:0]     dataInMem_hi_hi_lo_22 = {dataInMem_hi_675, dataInMem_lo_563, dataInMem_hi_674, dataInMem_lo_562};
  wire [447:0]     dataInMem_hi_hi_hi_22 = {dataInMem_hi_677, dataInMem_lo_565, dataInMem_hi_676, dataInMem_lo_564};
  wire [895:0]     dataInMem_hi_hi_454 = {dataInMem_hi_hi_hi_22, dataInMem_hi_hi_lo_22};
  wire [1791:0]    dataInMem_hi_678 = {dataInMem_hi_hi_454, dataInMem_hi_lo_230};
  wire [3583:0]    dataInMem_22 = {dataInMem_hi_678, dataInMem_lo_566};
  wire [511:0]     regroupCacheLine_22_0 = dataInMem_22[511:0];
  wire [511:0]     regroupCacheLine_22_1 = dataInMem_22[1023:512];
  wire [511:0]     regroupCacheLine_22_2 = dataInMem_22[1535:1024];
  wire [511:0]     regroupCacheLine_22_3 = dataInMem_22[2047:1536];
  wire [511:0]     regroupCacheLine_22_4 = dataInMem_22[2559:2048];
  wire [511:0]     regroupCacheLine_22_5 = dataInMem_22[3071:2560];
  wire [511:0]     regroupCacheLine_22_6 = dataInMem_22[3583:3072];
  wire [511:0]     res_176 = regroupCacheLine_22_0;
  wire [511:0]     res_177 = regroupCacheLine_22_1;
  wire [511:0]     res_178 = regroupCacheLine_22_2;
  wire [511:0]     res_179 = regroupCacheLine_22_3;
  wire [511:0]     res_180 = regroupCacheLine_22_4;
  wire [511:0]     res_181 = regroupCacheLine_22_5;
  wire [511:0]     res_182 = regroupCacheLine_22_6;
  wire [1023:0]    lo_lo_22 = {res_177, res_176};
  wire [1023:0]    lo_hi_22 = {res_179, res_178};
  wire [2047:0]    lo_22 = {lo_hi_22, lo_lo_22};
  wire [1023:0]    hi_lo_22 = {res_181, res_180};
  wire [1023:0]    hi_hi_22 = {512'h0, res_182};
  wire [2047:0]    hi_22 = {hi_hi_22, hi_lo_22};
  wire [4095:0]    regroupLoadData_2_6 = {hi_22, lo_22};
  wire [127:0]     dataInMem_lo_567 = {dataInMem_lo_hi_343, dataInMem_lo_lo_119};
  wire [63:0]      dataInMem_hi_hi_455 = {dataRegroupBySew_7_2_0, dataRegroupBySew_6_2_0};
  wire [127:0]     dataInMem_hi_679 = {dataInMem_hi_hi_455, dataInMem_hi_lo_231};
  wire [127:0]     dataInMem_lo_568 = {dataInMem_lo_hi_344, dataInMem_lo_lo_120};
  wire [63:0]      dataInMem_hi_hi_456 = {dataRegroupBySew_7_2_1, dataRegroupBySew_6_2_1};
  wire [127:0]     dataInMem_hi_680 = {dataInMem_hi_hi_456, dataInMem_hi_lo_232};
  wire [127:0]     dataInMem_lo_569 = {dataInMem_lo_hi_345, dataInMem_lo_lo_121};
  wire [63:0]      dataInMem_hi_hi_457 = {dataRegroupBySew_7_2_2, dataRegroupBySew_6_2_2};
  wire [127:0]     dataInMem_hi_681 = {dataInMem_hi_hi_457, dataInMem_hi_lo_233};
  wire [127:0]     dataInMem_lo_570 = {dataInMem_lo_hi_346, dataInMem_lo_lo_122};
  wire [63:0]      dataInMem_hi_hi_458 = {dataRegroupBySew_7_2_3, dataRegroupBySew_6_2_3};
  wire [127:0]     dataInMem_hi_682 = {dataInMem_hi_hi_458, dataInMem_hi_lo_234};
  wire [127:0]     dataInMem_lo_571 = {dataInMem_lo_hi_347, dataInMem_lo_lo_123};
  wire [63:0]      dataInMem_hi_hi_459 = {dataRegroupBySew_7_2_4, dataRegroupBySew_6_2_4};
  wire [127:0]     dataInMem_hi_683 = {dataInMem_hi_hi_459, dataInMem_hi_lo_235};
  wire [127:0]     dataInMem_lo_572 = {dataInMem_lo_hi_348, dataInMem_lo_lo_124};
  wire [63:0]      dataInMem_hi_hi_460 = {dataRegroupBySew_7_2_5, dataRegroupBySew_6_2_5};
  wire [127:0]     dataInMem_hi_684 = {dataInMem_hi_hi_460, dataInMem_hi_lo_236};
  wire [127:0]     dataInMem_lo_573 = {dataInMem_lo_hi_349, dataInMem_lo_lo_125};
  wire [63:0]      dataInMem_hi_hi_461 = {dataRegroupBySew_7_2_6, dataRegroupBySew_6_2_6};
  wire [127:0]     dataInMem_hi_685 = {dataInMem_hi_hi_461, dataInMem_hi_lo_237};
  wire [127:0]     dataInMem_lo_574 = {dataInMem_lo_hi_350, dataInMem_lo_lo_126};
  wire [63:0]      dataInMem_hi_hi_462 = {dataRegroupBySew_7_2_7, dataRegroupBySew_6_2_7};
  wire [127:0]     dataInMem_hi_686 = {dataInMem_hi_hi_462, dataInMem_hi_lo_238};
  wire [127:0]     dataInMem_lo_575 = {dataInMem_lo_hi_351, dataInMem_lo_lo_127};
  wire [63:0]      dataInMem_hi_hi_463 = {dataRegroupBySew_7_2_8, dataRegroupBySew_6_2_8};
  wire [127:0]     dataInMem_hi_687 = {dataInMem_hi_hi_463, dataInMem_hi_lo_239};
  wire [127:0]     dataInMem_lo_576 = {dataInMem_lo_hi_352, dataInMem_lo_lo_128};
  wire [63:0]      dataInMem_hi_hi_464 = {dataRegroupBySew_7_2_9, dataRegroupBySew_6_2_9};
  wire [127:0]     dataInMem_hi_688 = {dataInMem_hi_hi_464, dataInMem_hi_lo_240};
  wire [127:0]     dataInMem_lo_577 = {dataInMem_lo_hi_353, dataInMem_lo_lo_129};
  wire [63:0]      dataInMem_hi_hi_465 = {dataRegroupBySew_7_2_10, dataRegroupBySew_6_2_10};
  wire [127:0]     dataInMem_hi_689 = {dataInMem_hi_hi_465, dataInMem_hi_lo_241};
  wire [127:0]     dataInMem_lo_578 = {dataInMem_lo_hi_354, dataInMem_lo_lo_130};
  wire [63:0]      dataInMem_hi_hi_466 = {dataRegroupBySew_7_2_11, dataRegroupBySew_6_2_11};
  wire [127:0]     dataInMem_hi_690 = {dataInMem_hi_hi_466, dataInMem_hi_lo_242};
  wire [127:0]     dataInMem_lo_579 = {dataInMem_lo_hi_355, dataInMem_lo_lo_131};
  wire [63:0]      dataInMem_hi_hi_467 = {dataRegroupBySew_7_2_12, dataRegroupBySew_6_2_12};
  wire [127:0]     dataInMem_hi_691 = {dataInMem_hi_hi_467, dataInMem_hi_lo_243};
  wire [127:0]     dataInMem_lo_580 = {dataInMem_lo_hi_356, dataInMem_lo_lo_132};
  wire [63:0]      dataInMem_hi_hi_468 = {dataRegroupBySew_7_2_13, dataRegroupBySew_6_2_13};
  wire [127:0]     dataInMem_hi_692 = {dataInMem_hi_hi_468, dataInMem_hi_lo_244};
  wire [127:0]     dataInMem_lo_581 = {dataInMem_lo_hi_357, dataInMem_lo_lo_133};
  wire [63:0]      dataInMem_hi_hi_469 = {dataRegroupBySew_7_2_14, dataRegroupBySew_6_2_14};
  wire [127:0]     dataInMem_hi_693 = {dataInMem_hi_hi_469, dataInMem_hi_lo_245};
  wire [127:0]     dataInMem_lo_582 = {dataInMem_lo_hi_358, dataInMem_lo_lo_134};
  wire [63:0]      dataInMem_hi_hi_470 = {dataRegroupBySew_7_2_15, dataRegroupBySew_6_2_15};
  wire [127:0]     dataInMem_hi_694 = {dataInMem_hi_hi_470, dataInMem_hi_lo_246};
  wire [511:0]     dataInMem_lo_lo_lo_23 = {dataInMem_hi_680, dataInMem_lo_568, dataInMem_hi_679, dataInMem_lo_567};
  wire [511:0]     dataInMem_lo_lo_hi_23 = {dataInMem_hi_682, dataInMem_lo_570, dataInMem_hi_681, dataInMem_lo_569};
  wire [1023:0]    dataInMem_lo_lo_135 = {dataInMem_lo_lo_hi_23, dataInMem_lo_lo_lo_23};
  wire [511:0]     dataInMem_lo_hi_lo_23 = {dataInMem_hi_684, dataInMem_lo_572, dataInMem_hi_683, dataInMem_lo_571};
  wire [511:0]     dataInMem_lo_hi_hi_23 = {dataInMem_hi_686, dataInMem_lo_574, dataInMem_hi_685, dataInMem_lo_573};
  wire [1023:0]    dataInMem_lo_hi_359 = {dataInMem_lo_hi_hi_23, dataInMem_lo_hi_lo_23};
  wire [2047:0]    dataInMem_lo_583 = {dataInMem_lo_hi_359, dataInMem_lo_lo_135};
  wire [511:0]     dataInMem_hi_lo_lo_23 = {dataInMem_hi_688, dataInMem_lo_576, dataInMem_hi_687, dataInMem_lo_575};
  wire [511:0]     dataInMem_hi_lo_hi_23 = {dataInMem_hi_690, dataInMem_lo_578, dataInMem_hi_689, dataInMem_lo_577};
  wire [1023:0]    dataInMem_hi_lo_247 = {dataInMem_hi_lo_hi_23, dataInMem_hi_lo_lo_23};
  wire [511:0]     dataInMem_hi_hi_lo_23 = {dataInMem_hi_692, dataInMem_lo_580, dataInMem_hi_691, dataInMem_lo_579};
  wire [511:0]     dataInMem_hi_hi_hi_23 = {dataInMem_hi_694, dataInMem_lo_582, dataInMem_hi_693, dataInMem_lo_581};
  wire [1023:0]    dataInMem_hi_hi_471 = {dataInMem_hi_hi_hi_23, dataInMem_hi_hi_lo_23};
  wire [2047:0]    dataInMem_hi_695 = {dataInMem_hi_hi_471, dataInMem_hi_lo_247};
  wire [4095:0]    dataInMem_23 = {dataInMem_hi_695, dataInMem_lo_583};
  wire [511:0]     regroupCacheLine_23_0 = dataInMem_23[511:0];
  wire [511:0]     regroupCacheLine_23_1 = dataInMem_23[1023:512];
  wire [511:0]     regroupCacheLine_23_2 = dataInMem_23[1535:1024];
  wire [511:0]     regroupCacheLine_23_3 = dataInMem_23[2047:1536];
  wire [511:0]     regroupCacheLine_23_4 = dataInMem_23[2559:2048];
  wire [511:0]     regroupCacheLine_23_5 = dataInMem_23[3071:2560];
  wire [511:0]     regroupCacheLine_23_6 = dataInMem_23[3583:3072];
  wire [511:0]     regroupCacheLine_23_7 = dataInMem_23[4095:3584];
  wire [511:0]     res_184 = regroupCacheLine_23_0;
  wire [511:0]     res_185 = regroupCacheLine_23_1;
  wire [511:0]     res_186 = regroupCacheLine_23_2;
  wire [511:0]     res_187 = regroupCacheLine_23_3;
  wire [511:0]     res_188 = regroupCacheLine_23_4;
  wire [511:0]     res_189 = regroupCacheLine_23_5;
  wire [511:0]     res_190 = regroupCacheLine_23_6;
  wire [511:0]     res_191 = regroupCacheLine_23_7;
  wire [1023:0]    lo_lo_23 = {res_185, res_184};
  wire [1023:0]    lo_hi_23 = {res_187, res_186};
  wire [2047:0]    lo_23 = {lo_hi_23, lo_lo_23};
  wire [1023:0]    hi_lo_23 = {res_189, res_188};
  wire [1023:0]    hi_hi_23 = {res_191, res_190};
  wire [2047:0]    hi_23 = {hi_hi_23, hi_lo_23};
  wire [4095:0]    regroupLoadData_2_7 = {hi_23, lo_23};
  wire             _GEN_565 = lsuRequest_valid | accessBufferDequeueFire;
  wire             _GEN_566 = isLastDataGroup & ~isLastMaskGroup;
  wire             _maskSelect_valid_output = _GEN_565 & _GEN_566;
  wire [7:0][63:0] _GEN_567 = {{maskForBufferData_7}, {maskForBufferData_6}, {maskForBufferData_5}, {maskForBufferData_4}, {maskForBufferData_3}, {maskForBufferData_2}, {maskForBufferData_1}, {maskForBufferData_0}};
  wire [63:0]      _GEN_568 = _GEN_567[cacheLineIndexInBuffer];
  wire             needSendTail = {7'h0, bufferBaseCacheLineIndex} == cacheLineNumberReg;
  assign memRequest_valid_0 = (bufferValid | canSendTail & needSendTail) & addressQueueFree;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo = {cacheLineTemp[8], cacheLineTemp[0]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi = {cacheLineTemp[24], cacheLineTemp[16]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo = {cacheLineTemp[40], cacheLineTemp[32]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi = {cacheLineTemp[56], cacheLineTemp[48]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo = {cacheLineTemp[72], cacheLineTemp[64]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi = {cacheLineTemp[88], cacheLineTemp[80]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo = {cacheLineTemp[104], cacheLineTemp[96]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi = {cacheLineTemp[120], cacheLineTemp[112]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo = {cacheLineTemp[136], cacheLineTemp[128]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi = {cacheLineTemp[152], cacheLineTemp[144]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo = {memRequest_bits_data_lo_lo_hi_lo_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo = {cacheLineTemp[168], cacheLineTemp[160]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi = {cacheLineTemp[184], cacheLineTemp[176]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi = {memRequest_bits_data_lo_lo_hi_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo = {cacheLineTemp[200], cacheLineTemp[192]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi = {cacheLineTemp[216], cacheLineTemp[208]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo = {memRequest_bits_data_lo_lo_hi_hi_lo_hi, memRequest_bits_data_lo_lo_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo = {cacheLineTemp[232], cacheLineTemp[224]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi = {cacheLineTemp[248], cacheLineTemp[240]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_lo_hi = {memRequest_bits_data_lo_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo};
  wire [31:0]      memRequest_bits_data_lo_lo = {memRequest_bits_data_lo_lo_hi, memRequest_bits_data_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo = {cacheLineTemp[264], cacheLineTemp[256]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi = {cacheLineTemp[280], cacheLineTemp[272]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo = {cacheLineTemp[296], cacheLineTemp[288]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi = {cacheLineTemp[312], cacheLineTemp[304]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi = {memRequest_bits_data_lo_hi_lo_lo_hi_hi, memRequest_bits_data_lo_hi_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo = {cacheLineTemp[328], cacheLineTemp[320]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi = {cacheLineTemp[344], cacheLineTemp[336]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo = {cacheLineTemp[360], cacheLineTemp[352]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi = {cacheLineTemp[376], cacheLineTemp[368]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi = {memRequest_bits_data_lo_hi_lo_hi_hi_hi, memRequest_bits_data_lo_hi_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi = {memRequest_bits_data_lo_hi_lo_hi_hi, memRequest_bits_data_lo_hi_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo = {cacheLineTemp[392], cacheLineTemp[384]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi = {cacheLineTemp[408], cacheLineTemp[400]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo = {memRequest_bits_data_lo_hi_hi_lo_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo = {cacheLineTemp[424], cacheLineTemp[416]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi = {cacheLineTemp[440], cacheLineTemp[432]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi = {memRequest_bits_data_lo_hi_hi_lo_hi_hi, memRequest_bits_data_lo_hi_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo = {cacheLineTemp[456], cacheLineTemp[448]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi = {cacheLineTemp[472], cacheLineTemp[464]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo = {cacheLineTemp[488], cacheLineTemp[480]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi = {cacheLineTemp[504], cacheLineTemp[496]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_hi_hi = {memRequest_bits_data_lo_hi_hi_hi, memRequest_bits_data_lo_hi_hi_lo};
  wire [31:0]      memRequest_bits_data_lo_hi = {memRequest_bits_data_lo_hi_hi, memRequest_bits_data_lo_hi_lo};
  wire [63:0]      memRequest_bits_data_lo = {memRequest_bits_data_lo_hi, memRequest_bits_data_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo = {dataBuffer_0[8], dataBuffer_0[0]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi = {dataBuffer_0[24], dataBuffer_0[16]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo = {dataBuffer_0[40], dataBuffer_0[32]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi = {dataBuffer_0[56], dataBuffer_0[48]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo = {dataBuffer_0[72], dataBuffer_0[64]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi = {dataBuffer_0[88], dataBuffer_0[80]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo = {memRequest_bits_data_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_lo_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo = {dataBuffer_0[104], dataBuffer_0[96]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi = {dataBuffer_0[120], dataBuffer_0[112]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_lo_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_lo_lo = {memRequest_bits_data_hi_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo = {dataBuffer_0[136], dataBuffer_0[128]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi = {dataBuffer_0[152], dataBuffer_0[144]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo = {memRequest_bits_data_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo = {dataBuffer_0[168], dataBuffer_0[160]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi = {dataBuffer_0[184], dataBuffer_0[176]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo = {memRequest_bits_data_hi_lo_hi_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo = {dataBuffer_0[200], dataBuffer_0[192]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi = {dataBuffer_0[216], dataBuffer_0[208]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo = {memRequest_bits_data_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_lo_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo = {dataBuffer_0[232], dataBuffer_0[224]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi = {dataBuffer_0[248], dataBuffer_0[240]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo};
  wire [31:0]      memRequest_bits_data_hi_lo = {memRequest_bits_data_hi_lo_hi, memRequest_bits_data_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo = {dataBuffer_0[264], dataBuffer_0[256]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi = {dataBuffer_0[280], dataBuffer_0[272]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo = {dataBuffer_0[296], dataBuffer_0[288]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi = {dataBuffer_0[312], dataBuffer_0[304]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_hi_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo = {dataBuffer_0[328], dataBuffer_0[320]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi = {dataBuffer_0[344], dataBuffer_0[336]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo = {memRequest_bits_data_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_hi_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo = {dataBuffer_0[360], dataBuffer_0[352]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi = {dataBuffer_0[376], dataBuffer_0[368]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_hi_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_hi_lo = {memRequest_bits_data_hi_hi_lo_hi, memRequest_bits_data_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo = {dataBuffer_0[392], dataBuffer_0[384]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi = {dataBuffer_0[408], dataBuffer_0[400]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo = {dataBuffer_0[424], dataBuffer_0[416]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi = {dataBuffer_0[440], dataBuffer_0[432]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo = {dataBuffer_0[456], dataBuffer_0[448]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi = {dataBuffer_0[472], dataBuffer_0[464]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo = {dataBuffer_0[488], dataBuffer_0[480]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi = {dataBuffer_0[504], dataBuffer_0[496]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_lo};
  wire [31:0]      memRequest_bits_data_hi_hi = {memRequest_bits_data_hi_hi_hi, memRequest_bits_data_hi_hi_lo};
  wire [63:0]      memRequest_bits_data_hi = {memRequest_bits_data_hi_hi, memRequest_bits_data_hi_lo};
  wire [190:0]     _GEN_569 = {185'h0, initOffset};
  wire [190:0]     _memRequest_bits_data_T_1026 = {63'h0, memRequest_bits_data_hi, memRequest_bits_data_lo} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_1 = {cacheLineTemp[9], cacheLineTemp[1]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_1 = {cacheLineTemp[25], cacheLineTemp[17]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_1 = {cacheLineTemp[41], cacheLineTemp[33]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_1 = {cacheLineTemp[57], cacheLineTemp[49]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_1 = {cacheLineTemp[73], cacheLineTemp[65]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_1 = {cacheLineTemp[89], cacheLineTemp[81]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_1 = {cacheLineTemp[105], cacheLineTemp[97]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_1 = {cacheLineTemp[121], cacheLineTemp[113]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_1 = {cacheLineTemp[137], cacheLineTemp[129]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_1 = {cacheLineTemp[153], cacheLineTemp[145]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_1 = {cacheLineTemp[169], cacheLineTemp[161]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_1 = {cacheLineTemp[185], cacheLineTemp[177]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_1 = {cacheLineTemp[201], cacheLineTemp[193]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_1 = {cacheLineTemp[217], cacheLineTemp[209]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_1 = {cacheLineTemp[233], cacheLineTemp[225]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_1 = {cacheLineTemp[249], cacheLineTemp[241]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_1};
  wire [31:0]      memRequest_bits_data_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_1 = {cacheLineTemp[265], cacheLineTemp[257]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_1 = {cacheLineTemp[281], cacheLineTemp[273]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_1 = {cacheLineTemp[297], cacheLineTemp[289]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_1 = {cacheLineTemp[313], cacheLineTemp[305]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_1 = {cacheLineTemp[329], cacheLineTemp[321]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_1 = {cacheLineTemp[345], cacheLineTemp[337]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_1 = {cacheLineTemp[361], cacheLineTemp[353]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_1 = {cacheLineTemp[377], cacheLineTemp[369]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_1 = {cacheLineTemp[393], cacheLineTemp[385]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_1 = {cacheLineTemp[409], cacheLineTemp[401]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_1 = {cacheLineTemp[425], cacheLineTemp[417]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_1 = {cacheLineTemp[441], cacheLineTemp[433]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_1 = {cacheLineTemp[457], cacheLineTemp[449]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_1 = {cacheLineTemp[473], cacheLineTemp[465]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_1 = {cacheLineTemp[489], cacheLineTemp[481]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_1 = {cacheLineTemp[505], cacheLineTemp[497]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_1};
  wire [31:0]      memRequest_bits_data_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_1};
  wire [63:0]      memRequest_bits_data_lo_1 = {memRequest_bits_data_lo_hi_1, memRequest_bits_data_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_1 = {dataBuffer_0[9], dataBuffer_0[1]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_1 = {dataBuffer_0[25], dataBuffer_0[17]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_1 = {dataBuffer_0[41], dataBuffer_0[33]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_1 = {dataBuffer_0[57], dataBuffer_0[49]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_1 = {dataBuffer_0[73], dataBuffer_0[65]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_1 = {dataBuffer_0[89], dataBuffer_0[81]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_1 = {dataBuffer_0[105], dataBuffer_0[97]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_1 = {dataBuffer_0[121], dataBuffer_0[113]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_1 = {dataBuffer_0[137], dataBuffer_0[129]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_1 = {dataBuffer_0[153], dataBuffer_0[145]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_1 = {dataBuffer_0[169], dataBuffer_0[161]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_1 = {dataBuffer_0[185], dataBuffer_0[177]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_1 = {dataBuffer_0[201], dataBuffer_0[193]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_1 = {dataBuffer_0[217], dataBuffer_0[209]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_1 = {dataBuffer_0[233], dataBuffer_0[225]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_1 = {dataBuffer_0[249], dataBuffer_0[241]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_1};
  wire [31:0]      memRequest_bits_data_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_1 = {dataBuffer_0[265], dataBuffer_0[257]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_1 = {dataBuffer_0[281], dataBuffer_0[273]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_1 = {dataBuffer_0[297], dataBuffer_0[289]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_1 = {dataBuffer_0[313], dataBuffer_0[305]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_1 = {dataBuffer_0[329], dataBuffer_0[321]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_1 = {dataBuffer_0[345], dataBuffer_0[337]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_1 = {dataBuffer_0[361], dataBuffer_0[353]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_1 = {dataBuffer_0[377], dataBuffer_0[369]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_1 = {dataBuffer_0[393], dataBuffer_0[385]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_1 = {dataBuffer_0[409], dataBuffer_0[401]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_1 = {dataBuffer_0[425], dataBuffer_0[417]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_1 = {dataBuffer_0[441], dataBuffer_0[433]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_1 = {dataBuffer_0[457], dataBuffer_0[449]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_1 = {dataBuffer_0[473], dataBuffer_0[465]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_1 = {dataBuffer_0[489], dataBuffer_0[481]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_1 = {dataBuffer_0[505], dataBuffer_0[497]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_1};
  wire [31:0]      memRequest_bits_data_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_1};
  wire [63:0]      memRequest_bits_data_hi_1 = {memRequest_bits_data_hi_hi_1, memRequest_bits_data_hi_lo_1};
  wire [190:0]     _memRequest_bits_data_T_1219 = {63'h0, memRequest_bits_data_hi_1, memRequest_bits_data_lo_1} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_2 = {cacheLineTemp[10], cacheLineTemp[2]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_2 = {cacheLineTemp[26], cacheLineTemp[18]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_2 = {cacheLineTemp[42], cacheLineTemp[34]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_2 = {cacheLineTemp[58], cacheLineTemp[50]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_2 = {cacheLineTemp[74], cacheLineTemp[66]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_2 = {cacheLineTemp[90], cacheLineTemp[82]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_2 = {cacheLineTemp[106], cacheLineTemp[98]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_2 = {cacheLineTemp[122], cacheLineTemp[114]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_2 = {cacheLineTemp[138], cacheLineTemp[130]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_2 = {cacheLineTemp[154], cacheLineTemp[146]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_2 = {cacheLineTemp[170], cacheLineTemp[162]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_2 = {cacheLineTemp[186], cacheLineTemp[178]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_2 = {cacheLineTemp[202], cacheLineTemp[194]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_2 = {cacheLineTemp[218], cacheLineTemp[210]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_2 = {cacheLineTemp[234], cacheLineTemp[226]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_2 = {cacheLineTemp[250], cacheLineTemp[242]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_2};
  wire [31:0]      memRequest_bits_data_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_2 = {cacheLineTemp[266], cacheLineTemp[258]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_2 = {cacheLineTemp[282], cacheLineTemp[274]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_2 = {cacheLineTemp[298], cacheLineTemp[290]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_2 = {cacheLineTemp[314], cacheLineTemp[306]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_2 = {cacheLineTemp[330], cacheLineTemp[322]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_2 = {cacheLineTemp[346], cacheLineTemp[338]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_2 = {cacheLineTemp[362], cacheLineTemp[354]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_2 = {cacheLineTemp[378], cacheLineTemp[370]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_2 = {cacheLineTemp[394], cacheLineTemp[386]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_2 = {cacheLineTemp[410], cacheLineTemp[402]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_2 = {cacheLineTemp[426], cacheLineTemp[418]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_2 = {cacheLineTemp[442], cacheLineTemp[434]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_2 = {cacheLineTemp[458], cacheLineTemp[450]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_2 = {cacheLineTemp[474], cacheLineTemp[466]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_2 = {cacheLineTemp[490], cacheLineTemp[482]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_2 = {cacheLineTemp[506], cacheLineTemp[498]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_2};
  wire [31:0]      memRequest_bits_data_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_2};
  wire [63:0]      memRequest_bits_data_lo_2 = {memRequest_bits_data_lo_hi_2, memRequest_bits_data_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_2 = {dataBuffer_0[10], dataBuffer_0[2]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_2 = {dataBuffer_0[26], dataBuffer_0[18]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_2 = {dataBuffer_0[42], dataBuffer_0[34]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_2 = {dataBuffer_0[58], dataBuffer_0[50]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_2 = {dataBuffer_0[74], dataBuffer_0[66]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_2 = {dataBuffer_0[90], dataBuffer_0[82]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_2 = {dataBuffer_0[106], dataBuffer_0[98]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_2 = {dataBuffer_0[122], dataBuffer_0[114]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_2 = {dataBuffer_0[138], dataBuffer_0[130]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_2 = {dataBuffer_0[154], dataBuffer_0[146]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_2 = {dataBuffer_0[170], dataBuffer_0[162]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_2 = {dataBuffer_0[186], dataBuffer_0[178]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_2 = {dataBuffer_0[202], dataBuffer_0[194]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_2 = {dataBuffer_0[218], dataBuffer_0[210]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_2 = {dataBuffer_0[234], dataBuffer_0[226]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_2 = {dataBuffer_0[250], dataBuffer_0[242]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_2};
  wire [31:0]      memRequest_bits_data_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_2 = {dataBuffer_0[266], dataBuffer_0[258]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_2 = {dataBuffer_0[282], dataBuffer_0[274]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_2 = {dataBuffer_0[298], dataBuffer_0[290]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_2 = {dataBuffer_0[314], dataBuffer_0[306]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_2 = {dataBuffer_0[330], dataBuffer_0[322]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_2 = {dataBuffer_0[346], dataBuffer_0[338]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_2 = {dataBuffer_0[362], dataBuffer_0[354]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_2 = {dataBuffer_0[378], dataBuffer_0[370]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_2 = {dataBuffer_0[394], dataBuffer_0[386]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_2 = {dataBuffer_0[410], dataBuffer_0[402]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_2 = {dataBuffer_0[426], dataBuffer_0[418]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_2 = {dataBuffer_0[442], dataBuffer_0[434]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_2 = {dataBuffer_0[458], dataBuffer_0[450]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_2 = {dataBuffer_0[474], dataBuffer_0[466]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_2 = {dataBuffer_0[490], dataBuffer_0[482]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_2 = {dataBuffer_0[506], dataBuffer_0[498]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_2};
  wire [31:0]      memRequest_bits_data_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_2};
  wire [63:0]      memRequest_bits_data_hi_2 = {memRequest_bits_data_hi_hi_2, memRequest_bits_data_hi_lo_2};
  wire [190:0]     _memRequest_bits_data_T_1412 = {63'h0, memRequest_bits_data_hi_2, memRequest_bits_data_lo_2} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_3 = {cacheLineTemp[11], cacheLineTemp[3]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_3 = {cacheLineTemp[27], cacheLineTemp[19]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_3 = {cacheLineTemp[43], cacheLineTemp[35]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_3 = {cacheLineTemp[59], cacheLineTemp[51]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_3 = {cacheLineTemp[75], cacheLineTemp[67]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_3 = {cacheLineTemp[91], cacheLineTemp[83]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_3 = {cacheLineTemp[107], cacheLineTemp[99]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_3 = {cacheLineTemp[123], cacheLineTemp[115]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_3 = {cacheLineTemp[139], cacheLineTemp[131]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_3 = {cacheLineTemp[155], cacheLineTemp[147]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_3 = {cacheLineTemp[171], cacheLineTemp[163]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_3 = {cacheLineTemp[187], cacheLineTemp[179]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_3 = {cacheLineTemp[203], cacheLineTemp[195]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_3 = {cacheLineTemp[219], cacheLineTemp[211]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_3 = {cacheLineTemp[235], cacheLineTemp[227]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_3 = {cacheLineTemp[251], cacheLineTemp[243]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_3};
  wire [31:0]      memRequest_bits_data_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_3 = {cacheLineTemp[267], cacheLineTemp[259]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_3 = {cacheLineTemp[283], cacheLineTemp[275]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_3 = {cacheLineTemp[299], cacheLineTemp[291]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_3 = {cacheLineTemp[315], cacheLineTemp[307]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_3 = {cacheLineTemp[331], cacheLineTemp[323]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_3 = {cacheLineTemp[347], cacheLineTemp[339]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_3 = {cacheLineTemp[363], cacheLineTemp[355]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_3 = {cacheLineTemp[379], cacheLineTemp[371]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_3 = {cacheLineTemp[395], cacheLineTemp[387]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_3 = {cacheLineTemp[411], cacheLineTemp[403]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_3 = {cacheLineTemp[427], cacheLineTemp[419]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_3 = {cacheLineTemp[443], cacheLineTemp[435]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_3 = {cacheLineTemp[459], cacheLineTemp[451]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_3 = {cacheLineTemp[475], cacheLineTemp[467]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_3 = {cacheLineTemp[491], cacheLineTemp[483]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_3 = {cacheLineTemp[507], cacheLineTemp[499]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_3};
  wire [31:0]      memRequest_bits_data_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_3};
  wire [63:0]      memRequest_bits_data_lo_3 = {memRequest_bits_data_lo_hi_3, memRequest_bits_data_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_3 = {dataBuffer_0[11], dataBuffer_0[3]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_3 = {dataBuffer_0[27], dataBuffer_0[19]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_3 = {dataBuffer_0[43], dataBuffer_0[35]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_3 = {dataBuffer_0[59], dataBuffer_0[51]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_3 = {dataBuffer_0[75], dataBuffer_0[67]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_3 = {dataBuffer_0[91], dataBuffer_0[83]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_3 = {dataBuffer_0[107], dataBuffer_0[99]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_3 = {dataBuffer_0[123], dataBuffer_0[115]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_3 = {dataBuffer_0[139], dataBuffer_0[131]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_3 = {dataBuffer_0[155], dataBuffer_0[147]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_3 = {dataBuffer_0[171], dataBuffer_0[163]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_3 = {dataBuffer_0[187], dataBuffer_0[179]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_3 = {dataBuffer_0[203], dataBuffer_0[195]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_3 = {dataBuffer_0[219], dataBuffer_0[211]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_3 = {dataBuffer_0[235], dataBuffer_0[227]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_3 = {dataBuffer_0[251], dataBuffer_0[243]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_3};
  wire [31:0]      memRequest_bits_data_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_3 = {dataBuffer_0[267], dataBuffer_0[259]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_3 = {dataBuffer_0[283], dataBuffer_0[275]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_3 = {dataBuffer_0[299], dataBuffer_0[291]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_3 = {dataBuffer_0[315], dataBuffer_0[307]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_3 = {dataBuffer_0[331], dataBuffer_0[323]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_3 = {dataBuffer_0[347], dataBuffer_0[339]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_3 = {dataBuffer_0[363], dataBuffer_0[355]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_3 = {dataBuffer_0[379], dataBuffer_0[371]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_3 = {dataBuffer_0[395], dataBuffer_0[387]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_3 = {dataBuffer_0[411], dataBuffer_0[403]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_3 = {dataBuffer_0[427], dataBuffer_0[419]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_3 = {dataBuffer_0[443], dataBuffer_0[435]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_3 = {dataBuffer_0[459], dataBuffer_0[451]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_3 = {dataBuffer_0[475], dataBuffer_0[467]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_3 = {dataBuffer_0[491], dataBuffer_0[483]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_3 = {dataBuffer_0[507], dataBuffer_0[499]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_3};
  wire [31:0]      memRequest_bits_data_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_3};
  wire [63:0]      memRequest_bits_data_hi_3 = {memRequest_bits_data_hi_hi_3, memRequest_bits_data_hi_lo_3};
  wire [190:0]     _memRequest_bits_data_T_1605 = {63'h0, memRequest_bits_data_hi_3, memRequest_bits_data_lo_3} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_4 = {cacheLineTemp[12], cacheLineTemp[4]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_4 = {cacheLineTemp[28], cacheLineTemp[20]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_4 = {cacheLineTemp[44], cacheLineTemp[36]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_4 = {cacheLineTemp[60], cacheLineTemp[52]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_4 = {cacheLineTemp[76], cacheLineTemp[68]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_4 = {cacheLineTemp[92], cacheLineTemp[84]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_4 = {cacheLineTemp[108], cacheLineTemp[100]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_4 = {cacheLineTemp[124], cacheLineTemp[116]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_4 = {cacheLineTemp[140], cacheLineTemp[132]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_4 = {cacheLineTemp[156], cacheLineTemp[148]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_4 = {cacheLineTemp[172], cacheLineTemp[164]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_4 = {cacheLineTemp[188], cacheLineTemp[180]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_4 = {cacheLineTemp[204], cacheLineTemp[196]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_4 = {cacheLineTemp[220], cacheLineTemp[212]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_4 = {cacheLineTemp[236], cacheLineTemp[228]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_4 = {cacheLineTemp[252], cacheLineTemp[244]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_4};
  wire [31:0]      memRequest_bits_data_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_4 = {cacheLineTemp[268], cacheLineTemp[260]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_4 = {cacheLineTemp[284], cacheLineTemp[276]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_4 = {cacheLineTemp[300], cacheLineTemp[292]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_4 = {cacheLineTemp[316], cacheLineTemp[308]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_4 = {cacheLineTemp[332], cacheLineTemp[324]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_4 = {cacheLineTemp[348], cacheLineTemp[340]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_4 = {cacheLineTemp[364], cacheLineTemp[356]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_4 = {cacheLineTemp[380], cacheLineTemp[372]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_4 = {cacheLineTemp[396], cacheLineTemp[388]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_4 = {cacheLineTemp[412], cacheLineTemp[404]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_4 = {cacheLineTemp[428], cacheLineTemp[420]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_4 = {cacheLineTemp[444], cacheLineTemp[436]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_4 = {cacheLineTemp[460], cacheLineTemp[452]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_4 = {cacheLineTemp[476], cacheLineTemp[468]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_4 = {cacheLineTemp[492], cacheLineTemp[484]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_4 = {cacheLineTemp[508], cacheLineTemp[500]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_4};
  wire [31:0]      memRequest_bits_data_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_4};
  wire [63:0]      memRequest_bits_data_lo_4 = {memRequest_bits_data_lo_hi_4, memRequest_bits_data_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_4 = {dataBuffer_0[12], dataBuffer_0[4]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_4 = {dataBuffer_0[28], dataBuffer_0[20]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_4 = {dataBuffer_0[44], dataBuffer_0[36]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_4 = {dataBuffer_0[60], dataBuffer_0[52]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_4 = {dataBuffer_0[76], dataBuffer_0[68]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_4 = {dataBuffer_0[92], dataBuffer_0[84]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_4 = {dataBuffer_0[108], dataBuffer_0[100]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_4 = {dataBuffer_0[124], dataBuffer_0[116]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_4 = {dataBuffer_0[140], dataBuffer_0[132]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_4 = {dataBuffer_0[156], dataBuffer_0[148]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_4 = {dataBuffer_0[172], dataBuffer_0[164]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_4 = {dataBuffer_0[188], dataBuffer_0[180]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_4 = {dataBuffer_0[204], dataBuffer_0[196]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_4 = {dataBuffer_0[220], dataBuffer_0[212]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_4 = {dataBuffer_0[236], dataBuffer_0[228]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_4 = {dataBuffer_0[252], dataBuffer_0[244]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_4};
  wire [31:0]      memRequest_bits_data_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_4 = {dataBuffer_0[268], dataBuffer_0[260]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_4 = {dataBuffer_0[284], dataBuffer_0[276]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_4 = {dataBuffer_0[300], dataBuffer_0[292]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_4 = {dataBuffer_0[316], dataBuffer_0[308]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_4 = {dataBuffer_0[332], dataBuffer_0[324]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_4 = {dataBuffer_0[348], dataBuffer_0[340]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_4 = {dataBuffer_0[364], dataBuffer_0[356]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_4 = {dataBuffer_0[380], dataBuffer_0[372]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_4 = {dataBuffer_0[396], dataBuffer_0[388]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_4 = {dataBuffer_0[412], dataBuffer_0[404]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_4 = {dataBuffer_0[428], dataBuffer_0[420]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_4 = {dataBuffer_0[444], dataBuffer_0[436]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_4 = {dataBuffer_0[460], dataBuffer_0[452]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_4 = {dataBuffer_0[476], dataBuffer_0[468]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_4 = {dataBuffer_0[492], dataBuffer_0[484]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_4 = {dataBuffer_0[508], dataBuffer_0[500]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_4};
  wire [31:0]      memRequest_bits_data_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_4};
  wire [63:0]      memRequest_bits_data_hi_4 = {memRequest_bits_data_hi_hi_4, memRequest_bits_data_hi_lo_4};
  wire [190:0]     _memRequest_bits_data_T_1798 = {63'h0, memRequest_bits_data_hi_4, memRequest_bits_data_lo_4} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_5 = {cacheLineTemp[13], cacheLineTemp[5]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_5 = {cacheLineTemp[29], cacheLineTemp[21]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_5 = {cacheLineTemp[45], cacheLineTemp[37]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_5 = {cacheLineTemp[61], cacheLineTemp[53]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_5 = {cacheLineTemp[77], cacheLineTemp[69]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_5 = {cacheLineTemp[93], cacheLineTemp[85]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_5 = {cacheLineTemp[109], cacheLineTemp[101]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_5 = {cacheLineTemp[125], cacheLineTemp[117]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_5 = {cacheLineTemp[141], cacheLineTemp[133]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_5 = {cacheLineTemp[157], cacheLineTemp[149]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_5 = {cacheLineTemp[173], cacheLineTemp[165]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_5 = {cacheLineTemp[189], cacheLineTemp[181]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_5 = {cacheLineTemp[205], cacheLineTemp[197]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_5 = {cacheLineTemp[221], cacheLineTemp[213]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_5 = {cacheLineTemp[237], cacheLineTemp[229]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_5 = {cacheLineTemp[253], cacheLineTemp[245]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_5};
  wire [31:0]      memRequest_bits_data_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_5 = {cacheLineTemp[269], cacheLineTemp[261]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_5 = {cacheLineTemp[285], cacheLineTemp[277]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_5 = {cacheLineTemp[301], cacheLineTemp[293]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_5 = {cacheLineTemp[317], cacheLineTemp[309]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_5 = {cacheLineTemp[333], cacheLineTemp[325]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_5 = {cacheLineTemp[349], cacheLineTemp[341]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_5 = {cacheLineTemp[365], cacheLineTemp[357]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_5 = {cacheLineTemp[381], cacheLineTemp[373]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_5 = {cacheLineTemp[397], cacheLineTemp[389]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_5 = {cacheLineTemp[413], cacheLineTemp[405]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_5 = {cacheLineTemp[429], cacheLineTemp[421]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_5 = {cacheLineTemp[445], cacheLineTemp[437]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_5 = {cacheLineTemp[461], cacheLineTemp[453]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_5 = {cacheLineTemp[477], cacheLineTemp[469]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_5 = {cacheLineTemp[493], cacheLineTemp[485]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_5 = {cacheLineTemp[509], cacheLineTemp[501]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_5};
  wire [31:0]      memRequest_bits_data_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_5};
  wire [63:0]      memRequest_bits_data_lo_5 = {memRequest_bits_data_lo_hi_5, memRequest_bits_data_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_5 = {dataBuffer_0[13], dataBuffer_0[5]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_5 = {dataBuffer_0[29], dataBuffer_0[21]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_5 = {dataBuffer_0[45], dataBuffer_0[37]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_5 = {dataBuffer_0[61], dataBuffer_0[53]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_5 = {dataBuffer_0[77], dataBuffer_0[69]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_5 = {dataBuffer_0[93], dataBuffer_0[85]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_5 = {dataBuffer_0[109], dataBuffer_0[101]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_5 = {dataBuffer_0[125], dataBuffer_0[117]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_5 = {dataBuffer_0[141], dataBuffer_0[133]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_5 = {dataBuffer_0[157], dataBuffer_0[149]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_5 = {dataBuffer_0[173], dataBuffer_0[165]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_5 = {dataBuffer_0[189], dataBuffer_0[181]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_5 = {dataBuffer_0[205], dataBuffer_0[197]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_5 = {dataBuffer_0[221], dataBuffer_0[213]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_5 = {dataBuffer_0[237], dataBuffer_0[229]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_5 = {dataBuffer_0[253], dataBuffer_0[245]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_5};
  wire [31:0]      memRequest_bits_data_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_5 = {dataBuffer_0[269], dataBuffer_0[261]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_5 = {dataBuffer_0[285], dataBuffer_0[277]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_5 = {dataBuffer_0[301], dataBuffer_0[293]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_5 = {dataBuffer_0[317], dataBuffer_0[309]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_5 = {dataBuffer_0[333], dataBuffer_0[325]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_5 = {dataBuffer_0[349], dataBuffer_0[341]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_5 = {dataBuffer_0[365], dataBuffer_0[357]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_5 = {dataBuffer_0[381], dataBuffer_0[373]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_5 = {dataBuffer_0[397], dataBuffer_0[389]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_5 = {dataBuffer_0[413], dataBuffer_0[405]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_5 = {dataBuffer_0[429], dataBuffer_0[421]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_5 = {dataBuffer_0[445], dataBuffer_0[437]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_5 = {dataBuffer_0[461], dataBuffer_0[453]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_5 = {dataBuffer_0[477], dataBuffer_0[469]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_5 = {dataBuffer_0[493], dataBuffer_0[485]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_5 = {dataBuffer_0[509], dataBuffer_0[501]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_5};
  wire [31:0]      memRequest_bits_data_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_5};
  wire [63:0]      memRequest_bits_data_hi_5 = {memRequest_bits_data_hi_hi_5, memRequest_bits_data_hi_lo_5};
  wire [190:0]     _memRequest_bits_data_T_1991 = {63'h0, memRequest_bits_data_hi_5, memRequest_bits_data_lo_5} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_6 = {cacheLineTemp[14], cacheLineTemp[6]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_6 = {cacheLineTemp[30], cacheLineTemp[22]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_6 = {cacheLineTemp[46], cacheLineTemp[38]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_6 = {cacheLineTemp[62], cacheLineTemp[54]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_6 = {cacheLineTemp[78], cacheLineTemp[70]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_6 = {cacheLineTemp[94], cacheLineTemp[86]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_6 = {cacheLineTemp[110], cacheLineTemp[102]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_6 = {cacheLineTemp[126], cacheLineTemp[118]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_6 = {cacheLineTemp[142], cacheLineTemp[134]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_6 = {cacheLineTemp[158], cacheLineTemp[150]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_6 = {cacheLineTemp[174], cacheLineTemp[166]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_6 = {cacheLineTemp[190], cacheLineTemp[182]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_6 = {cacheLineTemp[206], cacheLineTemp[198]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_6 = {cacheLineTemp[222], cacheLineTemp[214]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_6 = {cacheLineTemp[238], cacheLineTemp[230]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_6 = {cacheLineTemp[254], cacheLineTemp[246]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_6};
  wire [31:0]      memRequest_bits_data_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_6 = {cacheLineTemp[270], cacheLineTemp[262]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_6 = {cacheLineTemp[286], cacheLineTemp[278]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_6 = {cacheLineTemp[302], cacheLineTemp[294]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_6 = {cacheLineTemp[318], cacheLineTemp[310]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_6 = {cacheLineTemp[334], cacheLineTemp[326]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_6 = {cacheLineTemp[350], cacheLineTemp[342]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_6 = {cacheLineTemp[366], cacheLineTemp[358]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_6 = {cacheLineTemp[382], cacheLineTemp[374]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_6 = {cacheLineTemp[398], cacheLineTemp[390]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_6 = {cacheLineTemp[414], cacheLineTemp[406]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_6 = {cacheLineTemp[430], cacheLineTemp[422]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_6 = {cacheLineTemp[446], cacheLineTemp[438]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_6 = {cacheLineTemp[462], cacheLineTemp[454]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_6 = {cacheLineTemp[478], cacheLineTemp[470]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_6 = {cacheLineTemp[494], cacheLineTemp[486]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_6 = {cacheLineTemp[510], cacheLineTemp[502]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_6};
  wire [31:0]      memRequest_bits_data_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_6};
  wire [63:0]      memRequest_bits_data_lo_6 = {memRequest_bits_data_lo_hi_6, memRequest_bits_data_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_6 = {dataBuffer_0[14], dataBuffer_0[6]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_6 = {dataBuffer_0[30], dataBuffer_0[22]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_6 = {dataBuffer_0[46], dataBuffer_0[38]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_6 = {dataBuffer_0[62], dataBuffer_0[54]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_6 = {dataBuffer_0[78], dataBuffer_0[70]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_6 = {dataBuffer_0[94], dataBuffer_0[86]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_6 = {dataBuffer_0[110], dataBuffer_0[102]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_6 = {dataBuffer_0[126], dataBuffer_0[118]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_6 = {dataBuffer_0[142], dataBuffer_0[134]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_6 = {dataBuffer_0[158], dataBuffer_0[150]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_6 = {dataBuffer_0[174], dataBuffer_0[166]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_6 = {dataBuffer_0[190], dataBuffer_0[182]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_6 = {dataBuffer_0[206], dataBuffer_0[198]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_6 = {dataBuffer_0[222], dataBuffer_0[214]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_6 = {dataBuffer_0[238], dataBuffer_0[230]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_6 = {dataBuffer_0[254], dataBuffer_0[246]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_6};
  wire [31:0]      memRequest_bits_data_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_6 = {dataBuffer_0[270], dataBuffer_0[262]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_6 = {dataBuffer_0[286], dataBuffer_0[278]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_6 = {dataBuffer_0[302], dataBuffer_0[294]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_6 = {dataBuffer_0[318], dataBuffer_0[310]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_6 = {dataBuffer_0[334], dataBuffer_0[326]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_6 = {dataBuffer_0[350], dataBuffer_0[342]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_6 = {dataBuffer_0[366], dataBuffer_0[358]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_6 = {dataBuffer_0[382], dataBuffer_0[374]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_6 = {dataBuffer_0[398], dataBuffer_0[390]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_6 = {dataBuffer_0[414], dataBuffer_0[406]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_6 = {dataBuffer_0[430], dataBuffer_0[422]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_6 = {dataBuffer_0[446], dataBuffer_0[438]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_6 = {dataBuffer_0[462], dataBuffer_0[454]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_6 = {dataBuffer_0[478], dataBuffer_0[470]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_6 = {dataBuffer_0[494], dataBuffer_0[486]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_6 = {dataBuffer_0[510], dataBuffer_0[502]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_6};
  wire [31:0]      memRequest_bits_data_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_6};
  wire [63:0]      memRequest_bits_data_hi_6 = {memRequest_bits_data_hi_hi_6, memRequest_bits_data_hi_lo_6};
  wire [190:0]     _memRequest_bits_data_T_2184 = {63'h0, memRequest_bits_data_hi_6, memRequest_bits_data_lo_6} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_7 = {cacheLineTemp[15], cacheLineTemp[7]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_7 = {cacheLineTemp[31], cacheLineTemp[23]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_7 = {cacheLineTemp[47], cacheLineTemp[39]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_7 = {cacheLineTemp[63], cacheLineTemp[55]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_7 = {cacheLineTemp[79], cacheLineTemp[71]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_7 = {cacheLineTemp[95], cacheLineTemp[87]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_7 = {cacheLineTemp[111], cacheLineTemp[103]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_7 = {cacheLineTemp[127], cacheLineTemp[119]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_7 = {cacheLineTemp[143], cacheLineTemp[135]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_7 = {cacheLineTemp[159], cacheLineTemp[151]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_7 = {cacheLineTemp[175], cacheLineTemp[167]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_7 = {cacheLineTemp[191], cacheLineTemp[183]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_7 = {cacheLineTemp[207], cacheLineTemp[199]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_7 = {cacheLineTemp[223], cacheLineTemp[215]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_7 = {cacheLineTemp[239], cacheLineTemp[231]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_7 = {cacheLineTemp[255], cacheLineTemp[247]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_7};
  wire [31:0]      memRequest_bits_data_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_7 = {cacheLineTemp[271], cacheLineTemp[263]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_7 = {cacheLineTemp[287], cacheLineTemp[279]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_7 = {cacheLineTemp[303], cacheLineTemp[295]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_7 = {cacheLineTemp[319], cacheLineTemp[311]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_7 = {cacheLineTemp[335], cacheLineTemp[327]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_7 = {cacheLineTemp[351], cacheLineTemp[343]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_7 = {cacheLineTemp[367], cacheLineTemp[359]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_7 = {cacheLineTemp[383], cacheLineTemp[375]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_7 = {cacheLineTemp[399], cacheLineTemp[391]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_7 = {cacheLineTemp[415], cacheLineTemp[407]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_7 = {cacheLineTemp[431], cacheLineTemp[423]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_7 = {cacheLineTemp[447], cacheLineTemp[439]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_7 = {cacheLineTemp[463], cacheLineTemp[455]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_7 = {cacheLineTemp[479], cacheLineTemp[471]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_7 = {cacheLineTemp[495], cacheLineTemp[487]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_7 = {cacheLineTemp[511], cacheLineTemp[503]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_7};
  wire [31:0]      memRequest_bits_data_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_7};
  wire [63:0]      memRequest_bits_data_lo_7 = {memRequest_bits_data_lo_hi_7, memRequest_bits_data_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_7 = {dataBuffer_0[15], dataBuffer_0[7]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_7 = {dataBuffer_0[31], dataBuffer_0[23]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_7 = {dataBuffer_0[47], dataBuffer_0[39]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_7 = {dataBuffer_0[63], dataBuffer_0[55]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_7 = {dataBuffer_0[79], dataBuffer_0[71]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_7 = {dataBuffer_0[95], dataBuffer_0[87]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_7 = {dataBuffer_0[111], dataBuffer_0[103]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_7 = {dataBuffer_0[127], dataBuffer_0[119]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_7 = {dataBuffer_0[143], dataBuffer_0[135]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_7 = {dataBuffer_0[159], dataBuffer_0[151]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_7 = {dataBuffer_0[175], dataBuffer_0[167]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_7 = {dataBuffer_0[191], dataBuffer_0[183]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_7 = {dataBuffer_0[207], dataBuffer_0[199]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_7 = {dataBuffer_0[223], dataBuffer_0[215]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_7 = {dataBuffer_0[239], dataBuffer_0[231]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_7 = {dataBuffer_0[255], dataBuffer_0[247]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_7};
  wire [31:0]      memRequest_bits_data_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_7 = {dataBuffer_0[271], dataBuffer_0[263]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_7 = {dataBuffer_0[287], dataBuffer_0[279]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_7 = {dataBuffer_0[303], dataBuffer_0[295]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_7 = {dataBuffer_0[319], dataBuffer_0[311]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_7 = {dataBuffer_0[335], dataBuffer_0[327]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_7 = {dataBuffer_0[351], dataBuffer_0[343]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_7 = {dataBuffer_0[367], dataBuffer_0[359]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_7 = {dataBuffer_0[383], dataBuffer_0[375]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_7 = {dataBuffer_0[399], dataBuffer_0[391]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_7 = {dataBuffer_0[415], dataBuffer_0[407]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_7 = {dataBuffer_0[431], dataBuffer_0[423]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_7 = {dataBuffer_0[447], dataBuffer_0[439]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_7 = {dataBuffer_0[463], dataBuffer_0[455]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_7 = {dataBuffer_0[479], dataBuffer_0[471]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_7 = {dataBuffer_0[495], dataBuffer_0[487]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_7 = {dataBuffer_0[511], dataBuffer_0[503]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_7};
  wire [31:0]      memRequest_bits_data_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_7};
  wire [63:0]      memRequest_bits_data_hi_7 = {memRequest_bits_data_hi_hi_7, memRequest_bits_data_hi_lo_7};
  wire [190:0]     _memRequest_bits_data_T_2377 = {63'h0, memRequest_bits_data_hi_7, memRequest_bits_data_lo_7} << _GEN_569;
  wire [1:0]       memRequest_bits_data_lo_lo_8 = {_memRequest_bits_data_T_1219[0], _memRequest_bits_data_T_1026[0]};
  wire [1:0]       memRequest_bits_data_lo_hi_8 = {_memRequest_bits_data_T_1605[0], _memRequest_bits_data_T_1412[0]};
  wire [3:0]       memRequest_bits_data_lo_8 = {memRequest_bits_data_lo_hi_8, memRequest_bits_data_lo_lo_8};
  wire [1:0]       memRequest_bits_data_hi_lo_8 = {_memRequest_bits_data_T_1991[0], _memRequest_bits_data_T_1798[0]};
  wire [1:0]       memRequest_bits_data_hi_hi_8 = {_memRequest_bits_data_T_2377[0], _memRequest_bits_data_T_2184[0]};
  wire [3:0]       memRequest_bits_data_hi_8 = {memRequest_bits_data_hi_hi_8, memRequest_bits_data_hi_lo_8};
  wire [1:0]       memRequest_bits_data_lo_lo_9 = {_memRequest_bits_data_T_1219[1], _memRequest_bits_data_T_1026[1]};
  wire [1:0]       memRequest_bits_data_lo_hi_9 = {_memRequest_bits_data_T_1605[1], _memRequest_bits_data_T_1412[1]};
  wire [3:0]       memRequest_bits_data_lo_9 = {memRequest_bits_data_lo_hi_9, memRequest_bits_data_lo_lo_9};
  wire [1:0]       memRequest_bits_data_hi_lo_9 = {_memRequest_bits_data_T_1991[1], _memRequest_bits_data_T_1798[1]};
  wire [1:0]       memRequest_bits_data_hi_hi_9 = {_memRequest_bits_data_T_2377[1], _memRequest_bits_data_T_2184[1]};
  wire [3:0]       memRequest_bits_data_hi_9 = {memRequest_bits_data_hi_hi_9, memRequest_bits_data_hi_lo_9};
  wire [1:0]       memRequest_bits_data_lo_lo_10 = {_memRequest_bits_data_T_1219[2], _memRequest_bits_data_T_1026[2]};
  wire [1:0]       memRequest_bits_data_lo_hi_10 = {_memRequest_bits_data_T_1605[2], _memRequest_bits_data_T_1412[2]};
  wire [3:0]       memRequest_bits_data_lo_10 = {memRequest_bits_data_lo_hi_10, memRequest_bits_data_lo_lo_10};
  wire [1:0]       memRequest_bits_data_hi_lo_10 = {_memRequest_bits_data_T_1991[2], _memRequest_bits_data_T_1798[2]};
  wire [1:0]       memRequest_bits_data_hi_hi_10 = {_memRequest_bits_data_T_2377[2], _memRequest_bits_data_T_2184[2]};
  wire [3:0]       memRequest_bits_data_hi_10 = {memRequest_bits_data_hi_hi_10, memRequest_bits_data_hi_lo_10};
  wire [1:0]       memRequest_bits_data_lo_lo_11 = {_memRequest_bits_data_T_1219[3], _memRequest_bits_data_T_1026[3]};
  wire [1:0]       memRequest_bits_data_lo_hi_11 = {_memRequest_bits_data_T_1605[3], _memRequest_bits_data_T_1412[3]};
  wire [3:0]       memRequest_bits_data_lo_11 = {memRequest_bits_data_lo_hi_11, memRequest_bits_data_lo_lo_11};
  wire [1:0]       memRequest_bits_data_hi_lo_11 = {_memRequest_bits_data_T_1991[3], _memRequest_bits_data_T_1798[3]};
  wire [1:0]       memRequest_bits_data_hi_hi_11 = {_memRequest_bits_data_T_2377[3], _memRequest_bits_data_T_2184[3]};
  wire [3:0]       memRequest_bits_data_hi_11 = {memRequest_bits_data_hi_hi_11, memRequest_bits_data_hi_lo_11};
  wire [1:0]       memRequest_bits_data_lo_lo_12 = {_memRequest_bits_data_T_1219[4], _memRequest_bits_data_T_1026[4]};
  wire [1:0]       memRequest_bits_data_lo_hi_12 = {_memRequest_bits_data_T_1605[4], _memRequest_bits_data_T_1412[4]};
  wire [3:0]       memRequest_bits_data_lo_12 = {memRequest_bits_data_lo_hi_12, memRequest_bits_data_lo_lo_12};
  wire [1:0]       memRequest_bits_data_hi_lo_12 = {_memRequest_bits_data_T_1991[4], _memRequest_bits_data_T_1798[4]};
  wire [1:0]       memRequest_bits_data_hi_hi_12 = {_memRequest_bits_data_T_2377[4], _memRequest_bits_data_T_2184[4]};
  wire [3:0]       memRequest_bits_data_hi_12 = {memRequest_bits_data_hi_hi_12, memRequest_bits_data_hi_lo_12};
  wire [1:0]       memRequest_bits_data_lo_lo_13 = {_memRequest_bits_data_T_1219[5], _memRequest_bits_data_T_1026[5]};
  wire [1:0]       memRequest_bits_data_lo_hi_13 = {_memRequest_bits_data_T_1605[5], _memRequest_bits_data_T_1412[5]};
  wire [3:0]       memRequest_bits_data_lo_13 = {memRequest_bits_data_lo_hi_13, memRequest_bits_data_lo_lo_13};
  wire [1:0]       memRequest_bits_data_hi_lo_13 = {_memRequest_bits_data_T_1991[5], _memRequest_bits_data_T_1798[5]};
  wire [1:0]       memRequest_bits_data_hi_hi_13 = {_memRequest_bits_data_T_2377[5], _memRequest_bits_data_T_2184[5]};
  wire [3:0]       memRequest_bits_data_hi_13 = {memRequest_bits_data_hi_hi_13, memRequest_bits_data_hi_lo_13};
  wire [1:0]       memRequest_bits_data_lo_lo_14 = {_memRequest_bits_data_T_1219[6], _memRequest_bits_data_T_1026[6]};
  wire [1:0]       memRequest_bits_data_lo_hi_14 = {_memRequest_bits_data_T_1605[6], _memRequest_bits_data_T_1412[6]};
  wire [3:0]       memRequest_bits_data_lo_14 = {memRequest_bits_data_lo_hi_14, memRequest_bits_data_lo_lo_14};
  wire [1:0]       memRequest_bits_data_hi_lo_14 = {_memRequest_bits_data_T_1991[6], _memRequest_bits_data_T_1798[6]};
  wire [1:0]       memRequest_bits_data_hi_hi_14 = {_memRequest_bits_data_T_2377[6], _memRequest_bits_data_T_2184[6]};
  wire [3:0]       memRequest_bits_data_hi_14 = {memRequest_bits_data_hi_hi_14, memRequest_bits_data_hi_lo_14};
  wire [1:0]       memRequest_bits_data_lo_lo_15 = {_memRequest_bits_data_T_1219[7], _memRequest_bits_data_T_1026[7]};
  wire [1:0]       memRequest_bits_data_lo_hi_15 = {_memRequest_bits_data_T_1605[7], _memRequest_bits_data_T_1412[7]};
  wire [3:0]       memRequest_bits_data_lo_15 = {memRequest_bits_data_lo_hi_15, memRequest_bits_data_lo_lo_15};
  wire [1:0]       memRequest_bits_data_hi_lo_15 = {_memRequest_bits_data_T_1991[7], _memRequest_bits_data_T_1798[7]};
  wire [1:0]       memRequest_bits_data_hi_hi_15 = {_memRequest_bits_data_T_2377[7], _memRequest_bits_data_T_2184[7]};
  wire [3:0]       memRequest_bits_data_hi_15 = {memRequest_bits_data_hi_hi_15, memRequest_bits_data_hi_lo_15};
  wire [1:0]       memRequest_bits_data_lo_lo_16 = {_memRequest_bits_data_T_1219[8], _memRequest_bits_data_T_1026[8]};
  wire [1:0]       memRequest_bits_data_lo_hi_16 = {_memRequest_bits_data_T_1605[8], _memRequest_bits_data_T_1412[8]};
  wire [3:0]       memRequest_bits_data_lo_16 = {memRequest_bits_data_lo_hi_16, memRequest_bits_data_lo_lo_16};
  wire [1:0]       memRequest_bits_data_hi_lo_16 = {_memRequest_bits_data_T_1991[8], _memRequest_bits_data_T_1798[8]};
  wire [1:0]       memRequest_bits_data_hi_hi_16 = {_memRequest_bits_data_T_2377[8], _memRequest_bits_data_T_2184[8]};
  wire [3:0]       memRequest_bits_data_hi_16 = {memRequest_bits_data_hi_hi_16, memRequest_bits_data_hi_lo_16};
  wire [1:0]       memRequest_bits_data_lo_lo_17 = {_memRequest_bits_data_T_1219[9], _memRequest_bits_data_T_1026[9]};
  wire [1:0]       memRequest_bits_data_lo_hi_17 = {_memRequest_bits_data_T_1605[9], _memRequest_bits_data_T_1412[9]};
  wire [3:0]       memRequest_bits_data_lo_17 = {memRequest_bits_data_lo_hi_17, memRequest_bits_data_lo_lo_17};
  wire [1:0]       memRequest_bits_data_hi_lo_17 = {_memRequest_bits_data_T_1991[9], _memRequest_bits_data_T_1798[9]};
  wire [1:0]       memRequest_bits_data_hi_hi_17 = {_memRequest_bits_data_T_2377[9], _memRequest_bits_data_T_2184[9]};
  wire [3:0]       memRequest_bits_data_hi_17 = {memRequest_bits_data_hi_hi_17, memRequest_bits_data_hi_lo_17};
  wire [1:0]       memRequest_bits_data_lo_lo_18 = {_memRequest_bits_data_T_1219[10], _memRequest_bits_data_T_1026[10]};
  wire [1:0]       memRequest_bits_data_lo_hi_18 = {_memRequest_bits_data_T_1605[10], _memRequest_bits_data_T_1412[10]};
  wire [3:0]       memRequest_bits_data_lo_18 = {memRequest_bits_data_lo_hi_18, memRequest_bits_data_lo_lo_18};
  wire [1:0]       memRequest_bits_data_hi_lo_18 = {_memRequest_bits_data_T_1991[10], _memRequest_bits_data_T_1798[10]};
  wire [1:0]       memRequest_bits_data_hi_hi_18 = {_memRequest_bits_data_T_2377[10], _memRequest_bits_data_T_2184[10]};
  wire [3:0]       memRequest_bits_data_hi_18 = {memRequest_bits_data_hi_hi_18, memRequest_bits_data_hi_lo_18};
  wire [1:0]       memRequest_bits_data_lo_lo_19 = {_memRequest_bits_data_T_1219[11], _memRequest_bits_data_T_1026[11]};
  wire [1:0]       memRequest_bits_data_lo_hi_19 = {_memRequest_bits_data_T_1605[11], _memRequest_bits_data_T_1412[11]};
  wire [3:0]       memRequest_bits_data_lo_19 = {memRequest_bits_data_lo_hi_19, memRequest_bits_data_lo_lo_19};
  wire [1:0]       memRequest_bits_data_hi_lo_19 = {_memRequest_bits_data_T_1991[11], _memRequest_bits_data_T_1798[11]};
  wire [1:0]       memRequest_bits_data_hi_hi_19 = {_memRequest_bits_data_T_2377[11], _memRequest_bits_data_T_2184[11]};
  wire [3:0]       memRequest_bits_data_hi_19 = {memRequest_bits_data_hi_hi_19, memRequest_bits_data_hi_lo_19};
  wire [1:0]       memRequest_bits_data_lo_lo_20 = {_memRequest_bits_data_T_1219[12], _memRequest_bits_data_T_1026[12]};
  wire [1:0]       memRequest_bits_data_lo_hi_20 = {_memRequest_bits_data_T_1605[12], _memRequest_bits_data_T_1412[12]};
  wire [3:0]       memRequest_bits_data_lo_20 = {memRequest_bits_data_lo_hi_20, memRequest_bits_data_lo_lo_20};
  wire [1:0]       memRequest_bits_data_hi_lo_20 = {_memRequest_bits_data_T_1991[12], _memRequest_bits_data_T_1798[12]};
  wire [1:0]       memRequest_bits_data_hi_hi_20 = {_memRequest_bits_data_T_2377[12], _memRequest_bits_data_T_2184[12]};
  wire [3:0]       memRequest_bits_data_hi_20 = {memRequest_bits_data_hi_hi_20, memRequest_bits_data_hi_lo_20};
  wire [1:0]       memRequest_bits_data_lo_lo_21 = {_memRequest_bits_data_T_1219[13], _memRequest_bits_data_T_1026[13]};
  wire [1:0]       memRequest_bits_data_lo_hi_21 = {_memRequest_bits_data_T_1605[13], _memRequest_bits_data_T_1412[13]};
  wire [3:0]       memRequest_bits_data_lo_21 = {memRequest_bits_data_lo_hi_21, memRequest_bits_data_lo_lo_21};
  wire [1:0]       memRequest_bits_data_hi_lo_21 = {_memRequest_bits_data_T_1991[13], _memRequest_bits_data_T_1798[13]};
  wire [1:0]       memRequest_bits_data_hi_hi_21 = {_memRequest_bits_data_T_2377[13], _memRequest_bits_data_T_2184[13]};
  wire [3:0]       memRequest_bits_data_hi_21 = {memRequest_bits_data_hi_hi_21, memRequest_bits_data_hi_lo_21};
  wire [1:0]       memRequest_bits_data_lo_lo_22 = {_memRequest_bits_data_T_1219[14], _memRequest_bits_data_T_1026[14]};
  wire [1:0]       memRequest_bits_data_lo_hi_22 = {_memRequest_bits_data_T_1605[14], _memRequest_bits_data_T_1412[14]};
  wire [3:0]       memRequest_bits_data_lo_22 = {memRequest_bits_data_lo_hi_22, memRequest_bits_data_lo_lo_22};
  wire [1:0]       memRequest_bits_data_hi_lo_22 = {_memRequest_bits_data_T_1991[14], _memRequest_bits_data_T_1798[14]};
  wire [1:0]       memRequest_bits_data_hi_hi_22 = {_memRequest_bits_data_T_2377[14], _memRequest_bits_data_T_2184[14]};
  wire [3:0]       memRequest_bits_data_hi_22 = {memRequest_bits_data_hi_hi_22, memRequest_bits_data_hi_lo_22};
  wire [1:0]       memRequest_bits_data_lo_lo_23 = {_memRequest_bits_data_T_1219[15], _memRequest_bits_data_T_1026[15]};
  wire [1:0]       memRequest_bits_data_lo_hi_23 = {_memRequest_bits_data_T_1605[15], _memRequest_bits_data_T_1412[15]};
  wire [3:0]       memRequest_bits_data_lo_23 = {memRequest_bits_data_lo_hi_23, memRequest_bits_data_lo_lo_23};
  wire [1:0]       memRequest_bits_data_hi_lo_23 = {_memRequest_bits_data_T_1991[15], _memRequest_bits_data_T_1798[15]};
  wire [1:0]       memRequest_bits_data_hi_hi_23 = {_memRequest_bits_data_T_2377[15], _memRequest_bits_data_T_2184[15]};
  wire [3:0]       memRequest_bits_data_hi_23 = {memRequest_bits_data_hi_hi_23, memRequest_bits_data_hi_lo_23};
  wire [1:0]       memRequest_bits_data_lo_lo_24 = {_memRequest_bits_data_T_1219[16], _memRequest_bits_data_T_1026[16]};
  wire [1:0]       memRequest_bits_data_lo_hi_24 = {_memRequest_bits_data_T_1605[16], _memRequest_bits_data_T_1412[16]};
  wire [3:0]       memRequest_bits_data_lo_24 = {memRequest_bits_data_lo_hi_24, memRequest_bits_data_lo_lo_24};
  wire [1:0]       memRequest_bits_data_hi_lo_24 = {_memRequest_bits_data_T_1991[16], _memRequest_bits_data_T_1798[16]};
  wire [1:0]       memRequest_bits_data_hi_hi_24 = {_memRequest_bits_data_T_2377[16], _memRequest_bits_data_T_2184[16]};
  wire [3:0]       memRequest_bits_data_hi_24 = {memRequest_bits_data_hi_hi_24, memRequest_bits_data_hi_lo_24};
  wire [1:0]       memRequest_bits_data_lo_lo_25 = {_memRequest_bits_data_T_1219[17], _memRequest_bits_data_T_1026[17]};
  wire [1:0]       memRequest_bits_data_lo_hi_25 = {_memRequest_bits_data_T_1605[17], _memRequest_bits_data_T_1412[17]};
  wire [3:0]       memRequest_bits_data_lo_25 = {memRequest_bits_data_lo_hi_25, memRequest_bits_data_lo_lo_25};
  wire [1:0]       memRequest_bits_data_hi_lo_25 = {_memRequest_bits_data_T_1991[17], _memRequest_bits_data_T_1798[17]};
  wire [1:0]       memRequest_bits_data_hi_hi_25 = {_memRequest_bits_data_T_2377[17], _memRequest_bits_data_T_2184[17]};
  wire [3:0]       memRequest_bits_data_hi_25 = {memRequest_bits_data_hi_hi_25, memRequest_bits_data_hi_lo_25};
  wire [1:0]       memRequest_bits_data_lo_lo_26 = {_memRequest_bits_data_T_1219[18], _memRequest_bits_data_T_1026[18]};
  wire [1:0]       memRequest_bits_data_lo_hi_26 = {_memRequest_bits_data_T_1605[18], _memRequest_bits_data_T_1412[18]};
  wire [3:0]       memRequest_bits_data_lo_26 = {memRequest_bits_data_lo_hi_26, memRequest_bits_data_lo_lo_26};
  wire [1:0]       memRequest_bits_data_hi_lo_26 = {_memRequest_bits_data_T_1991[18], _memRequest_bits_data_T_1798[18]};
  wire [1:0]       memRequest_bits_data_hi_hi_26 = {_memRequest_bits_data_T_2377[18], _memRequest_bits_data_T_2184[18]};
  wire [3:0]       memRequest_bits_data_hi_26 = {memRequest_bits_data_hi_hi_26, memRequest_bits_data_hi_lo_26};
  wire [1:0]       memRequest_bits_data_lo_lo_27 = {_memRequest_bits_data_T_1219[19], _memRequest_bits_data_T_1026[19]};
  wire [1:0]       memRequest_bits_data_lo_hi_27 = {_memRequest_bits_data_T_1605[19], _memRequest_bits_data_T_1412[19]};
  wire [3:0]       memRequest_bits_data_lo_27 = {memRequest_bits_data_lo_hi_27, memRequest_bits_data_lo_lo_27};
  wire [1:0]       memRequest_bits_data_hi_lo_27 = {_memRequest_bits_data_T_1991[19], _memRequest_bits_data_T_1798[19]};
  wire [1:0]       memRequest_bits_data_hi_hi_27 = {_memRequest_bits_data_T_2377[19], _memRequest_bits_data_T_2184[19]};
  wire [3:0]       memRequest_bits_data_hi_27 = {memRequest_bits_data_hi_hi_27, memRequest_bits_data_hi_lo_27};
  wire [1:0]       memRequest_bits_data_lo_lo_28 = {_memRequest_bits_data_T_1219[20], _memRequest_bits_data_T_1026[20]};
  wire [1:0]       memRequest_bits_data_lo_hi_28 = {_memRequest_bits_data_T_1605[20], _memRequest_bits_data_T_1412[20]};
  wire [3:0]       memRequest_bits_data_lo_28 = {memRequest_bits_data_lo_hi_28, memRequest_bits_data_lo_lo_28};
  wire [1:0]       memRequest_bits_data_hi_lo_28 = {_memRequest_bits_data_T_1991[20], _memRequest_bits_data_T_1798[20]};
  wire [1:0]       memRequest_bits_data_hi_hi_28 = {_memRequest_bits_data_T_2377[20], _memRequest_bits_data_T_2184[20]};
  wire [3:0]       memRequest_bits_data_hi_28 = {memRequest_bits_data_hi_hi_28, memRequest_bits_data_hi_lo_28};
  wire [1:0]       memRequest_bits_data_lo_lo_29 = {_memRequest_bits_data_T_1219[21], _memRequest_bits_data_T_1026[21]};
  wire [1:0]       memRequest_bits_data_lo_hi_29 = {_memRequest_bits_data_T_1605[21], _memRequest_bits_data_T_1412[21]};
  wire [3:0]       memRequest_bits_data_lo_29 = {memRequest_bits_data_lo_hi_29, memRequest_bits_data_lo_lo_29};
  wire [1:0]       memRequest_bits_data_hi_lo_29 = {_memRequest_bits_data_T_1991[21], _memRequest_bits_data_T_1798[21]};
  wire [1:0]       memRequest_bits_data_hi_hi_29 = {_memRequest_bits_data_T_2377[21], _memRequest_bits_data_T_2184[21]};
  wire [3:0]       memRequest_bits_data_hi_29 = {memRequest_bits_data_hi_hi_29, memRequest_bits_data_hi_lo_29};
  wire [1:0]       memRequest_bits_data_lo_lo_30 = {_memRequest_bits_data_T_1219[22], _memRequest_bits_data_T_1026[22]};
  wire [1:0]       memRequest_bits_data_lo_hi_30 = {_memRequest_bits_data_T_1605[22], _memRequest_bits_data_T_1412[22]};
  wire [3:0]       memRequest_bits_data_lo_30 = {memRequest_bits_data_lo_hi_30, memRequest_bits_data_lo_lo_30};
  wire [1:0]       memRequest_bits_data_hi_lo_30 = {_memRequest_bits_data_T_1991[22], _memRequest_bits_data_T_1798[22]};
  wire [1:0]       memRequest_bits_data_hi_hi_30 = {_memRequest_bits_data_T_2377[22], _memRequest_bits_data_T_2184[22]};
  wire [3:0]       memRequest_bits_data_hi_30 = {memRequest_bits_data_hi_hi_30, memRequest_bits_data_hi_lo_30};
  wire [1:0]       memRequest_bits_data_lo_lo_31 = {_memRequest_bits_data_T_1219[23], _memRequest_bits_data_T_1026[23]};
  wire [1:0]       memRequest_bits_data_lo_hi_31 = {_memRequest_bits_data_T_1605[23], _memRequest_bits_data_T_1412[23]};
  wire [3:0]       memRequest_bits_data_lo_31 = {memRequest_bits_data_lo_hi_31, memRequest_bits_data_lo_lo_31};
  wire [1:0]       memRequest_bits_data_hi_lo_31 = {_memRequest_bits_data_T_1991[23], _memRequest_bits_data_T_1798[23]};
  wire [1:0]       memRequest_bits_data_hi_hi_31 = {_memRequest_bits_data_T_2377[23], _memRequest_bits_data_T_2184[23]};
  wire [3:0]       memRequest_bits_data_hi_31 = {memRequest_bits_data_hi_hi_31, memRequest_bits_data_hi_lo_31};
  wire [1:0]       memRequest_bits_data_lo_lo_32 = {_memRequest_bits_data_T_1219[24], _memRequest_bits_data_T_1026[24]};
  wire [1:0]       memRequest_bits_data_lo_hi_32 = {_memRequest_bits_data_T_1605[24], _memRequest_bits_data_T_1412[24]};
  wire [3:0]       memRequest_bits_data_lo_32 = {memRequest_bits_data_lo_hi_32, memRequest_bits_data_lo_lo_32};
  wire [1:0]       memRequest_bits_data_hi_lo_32 = {_memRequest_bits_data_T_1991[24], _memRequest_bits_data_T_1798[24]};
  wire [1:0]       memRequest_bits_data_hi_hi_32 = {_memRequest_bits_data_T_2377[24], _memRequest_bits_data_T_2184[24]};
  wire [3:0]       memRequest_bits_data_hi_32 = {memRequest_bits_data_hi_hi_32, memRequest_bits_data_hi_lo_32};
  wire [1:0]       memRequest_bits_data_lo_lo_33 = {_memRequest_bits_data_T_1219[25], _memRequest_bits_data_T_1026[25]};
  wire [1:0]       memRequest_bits_data_lo_hi_33 = {_memRequest_bits_data_T_1605[25], _memRequest_bits_data_T_1412[25]};
  wire [3:0]       memRequest_bits_data_lo_33 = {memRequest_bits_data_lo_hi_33, memRequest_bits_data_lo_lo_33};
  wire [1:0]       memRequest_bits_data_hi_lo_33 = {_memRequest_bits_data_T_1991[25], _memRequest_bits_data_T_1798[25]};
  wire [1:0]       memRequest_bits_data_hi_hi_33 = {_memRequest_bits_data_T_2377[25], _memRequest_bits_data_T_2184[25]};
  wire [3:0]       memRequest_bits_data_hi_33 = {memRequest_bits_data_hi_hi_33, memRequest_bits_data_hi_lo_33};
  wire [1:0]       memRequest_bits_data_lo_lo_34 = {_memRequest_bits_data_T_1219[26], _memRequest_bits_data_T_1026[26]};
  wire [1:0]       memRequest_bits_data_lo_hi_34 = {_memRequest_bits_data_T_1605[26], _memRequest_bits_data_T_1412[26]};
  wire [3:0]       memRequest_bits_data_lo_34 = {memRequest_bits_data_lo_hi_34, memRequest_bits_data_lo_lo_34};
  wire [1:0]       memRequest_bits_data_hi_lo_34 = {_memRequest_bits_data_T_1991[26], _memRequest_bits_data_T_1798[26]};
  wire [1:0]       memRequest_bits_data_hi_hi_34 = {_memRequest_bits_data_T_2377[26], _memRequest_bits_data_T_2184[26]};
  wire [3:0]       memRequest_bits_data_hi_34 = {memRequest_bits_data_hi_hi_34, memRequest_bits_data_hi_lo_34};
  wire [1:0]       memRequest_bits_data_lo_lo_35 = {_memRequest_bits_data_T_1219[27], _memRequest_bits_data_T_1026[27]};
  wire [1:0]       memRequest_bits_data_lo_hi_35 = {_memRequest_bits_data_T_1605[27], _memRequest_bits_data_T_1412[27]};
  wire [3:0]       memRequest_bits_data_lo_35 = {memRequest_bits_data_lo_hi_35, memRequest_bits_data_lo_lo_35};
  wire [1:0]       memRequest_bits_data_hi_lo_35 = {_memRequest_bits_data_T_1991[27], _memRequest_bits_data_T_1798[27]};
  wire [1:0]       memRequest_bits_data_hi_hi_35 = {_memRequest_bits_data_T_2377[27], _memRequest_bits_data_T_2184[27]};
  wire [3:0]       memRequest_bits_data_hi_35 = {memRequest_bits_data_hi_hi_35, memRequest_bits_data_hi_lo_35};
  wire [1:0]       memRequest_bits_data_lo_lo_36 = {_memRequest_bits_data_T_1219[28], _memRequest_bits_data_T_1026[28]};
  wire [1:0]       memRequest_bits_data_lo_hi_36 = {_memRequest_bits_data_T_1605[28], _memRequest_bits_data_T_1412[28]};
  wire [3:0]       memRequest_bits_data_lo_36 = {memRequest_bits_data_lo_hi_36, memRequest_bits_data_lo_lo_36};
  wire [1:0]       memRequest_bits_data_hi_lo_36 = {_memRequest_bits_data_T_1991[28], _memRequest_bits_data_T_1798[28]};
  wire [1:0]       memRequest_bits_data_hi_hi_36 = {_memRequest_bits_data_T_2377[28], _memRequest_bits_data_T_2184[28]};
  wire [3:0]       memRequest_bits_data_hi_36 = {memRequest_bits_data_hi_hi_36, memRequest_bits_data_hi_lo_36};
  wire [1:0]       memRequest_bits_data_lo_lo_37 = {_memRequest_bits_data_T_1219[29], _memRequest_bits_data_T_1026[29]};
  wire [1:0]       memRequest_bits_data_lo_hi_37 = {_memRequest_bits_data_T_1605[29], _memRequest_bits_data_T_1412[29]};
  wire [3:0]       memRequest_bits_data_lo_37 = {memRequest_bits_data_lo_hi_37, memRequest_bits_data_lo_lo_37};
  wire [1:0]       memRequest_bits_data_hi_lo_37 = {_memRequest_bits_data_T_1991[29], _memRequest_bits_data_T_1798[29]};
  wire [1:0]       memRequest_bits_data_hi_hi_37 = {_memRequest_bits_data_T_2377[29], _memRequest_bits_data_T_2184[29]};
  wire [3:0]       memRequest_bits_data_hi_37 = {memRequest_bits_data_hi_hi_37, memRequest_bits_data_hi_lo_37};
  wire [1:0]       memRequest_bits_data_lo_lo_38 = {_memRequest_bits_data_T_1219[30], _memRequest_bits_data_T_1026[30]};
  wire [1:0]       memRequest_bits_data_lo_hi_38 = {_memRequest_bits_data_T_1605[30], _memRequest_bits_data_T_1412[30]};
  wire [3:0]       memRequest_bits_data_lo_38 = {memRequest_bits_data_lo_hi_38, memRequest_bits_data_lo_lo_38};
  wire [1:0]       memRequest_bits_data_hi_lo_38 = {_memRequest_bits_data_T_1991[30], _memRequest_bits_data_T_1798[30]};
  wire [1:0]       memRequest_bits_data_hi_hi_38 = {_memRequest_bits_data_T_2377[30], _memRequest_bits_data_T_2184[30]};
  wire [3:0]       memRequest_bits_data_hi_38 = {memRequest_bits_data_hi_hi_38, memRequest_bits_data_hi_lo_38};
  wire [1:0]       memRequest_bits_data_lo_lo_39 = {_memRequest_bits_data_T_1219[31], _memRequest_bits_data_T_1026[31]};
  wire [1:0]       memRequest_bits_data_lo_hi_39 = {_memRequest_bits_data_T_1605[31], _memRequest_bits_data_T_1412[31]};
  wire [3:0]       memRequest_bits_data_lo_39 = {memRequest_bits_data_lo_hi_39, memRequest_bits_data_lo_lo_39};
  wire [1:0]       memRequest_bits_data_hi_lo_39 = {_memRequest_bits_data_T_1991[31], _memRequest_bits_data_T_1798[31]};
  wire [1:0]       memRequest_bits_data_hi_hi_39 = {_memRequest_bits_data_T_2377[31], _memRequest_bits_data_T_2184[31]};
  wire [3:0]       memRequest_bits_data_hi_39 = {memRequest_bits_data_hi_hi_39, memRequest_bits_data_hi_lo_39};
  wire [1:0]       memRequest_bits_data_lo_lo_40 = {_memRequest_bits_data_T_1219[32], _memRequest_bits_data_T_1026[32]};
  wire [1:0]       memRequest_bits_data_lo_hi_40 = {_memRequest_bits_data_T_1605[32], _memRequest_bits_data_T_1412[32]};
  wire [3:0]       memRequest_bits_data_lo_40 = {memRequest_bits_data_lo_hi_40, memRequest_bits_data_lo_lo_40};
  wire [1:0]       memRequest_bits_data_hi_lo_40 = {_memRequest_bits_data_T_1991[32], _memRequest_bits_data_T_1798[32]};
  wire [1:0]       memRequest_bits_data_hi_hi_40 = {_memRequest_bits_data_T_2377[32], _memRequest_bits_data_T_2184[32]};
  wire [3:0]       memRequest_bits_data_hi_40 = {memRequest_bits_data_hi_hi_40, memRequest_bits_data_hi_lo_40};
  wire [1:0]       memRequest_bits_data_lo_lo_41 = {_memRequest_bits_data_T_1219[33], _memRequest_bits_data_T_1026[33]};
  wire [1:0]       memRequest_bits_data_lo_hi_41 = {_memRequest_bits_data_T_1605[33], _memRequest_bits_data_T_1412[33]};
  wire [3:0]       memRequest_bits_data_lo_41 = {memRequest_bits_data_lo_hi_41, memRequest_bits_data_lo_lo_41};
  wire [1:0]       memRequest_bits_data_hi_lo_41 = {_memRequest_bits_data_T_1991[33], _memRequest_bits_data_T_1798[33]};
  wire [1:0]       memRequest_bits_data_hi_hi_41 = {_memRequest_bits_data_T_2377[33], _memRequest_bits_data_T_2184[33]};
  wire [3:0]       memRequest_bits_data_hi_41 = {memRequest_bits_data_hi_hi_41, memRequest_bits_data_hi_lo_41};
  wire [1:0]       memRequest_bits_data_lo_lo_42 = {_memRequest_bits_data_T_1219[34], _memRequest_bits_data_T_1026[34]};
  wire [1:0]       memRequest_bits_data_lo_hi_42 = {_memRequest_bits_data_T_1605[34], _memRequest_bits_data_T_1412[34]};
  wire [3:0]       memRequest_bits_data_lo_42 = {memRequest_bits_data_lo_hi_42, memRequest_bits_data_lo_lo_42};
  wire [1:0]       memRequest_bits_data_hi_lo_42 = {_memRequest_bits_data_T_1991[34], _memRequest_bits_data_T_1798[34]};
  wire [1:0]       memRequest_bits_data_hi_hi_42 = {_memRequest_bits_data_T_2377[34], _memRequest_bits_data_T_2184[34]};
  wire [3:0]       memRequest_bits_data_hi_42 = {memRequest_bits_data_hi_hi_42, memRequest_bits_data_hi_lo_42};
  wire [1:0]       memRequest_bits_data_lo_lo_43 = {_memRequest_bits_data_T_1219[35], _memRequest_bits_data_T_1026[35]};
  wire [1:0]       memRequest_bits_data_lo_hi_43 = {_memRequest_bits_data_T_1605[35], _memRequest_bits_data_T_1412[35]};
  wire [3:0]       memRequest_bits_data_lo_43 = {memRequest_bits_data_lo_hi_43, memRequest_bits_data_lo_lo_43};
  wire [1:0]       memRequest_bits_data_hi_lo_43 = {_memRequest_bits_data_T_1991[35], _memRequest_bits_data_T_1798[35]};
  wire [1:0]       memRequest_bits_data_hi_hi_43 = {_memRequest_bits_data_T_2377[35], _memRequest_bits_data_T_2184[35]};
  wire [3:0]       memRequest_bits_data_hi_43 = {memRequest_bits_data_hi_hi_43, memRequest_bits_data_hi_lo_43};
  wire [1:0]       memRequest_bits_data_lo_lo_44 = {_memRequest_bits_data_T_1219[36], _memRequest_bits_data_T_1026[36]};
  wire [1:0]       memRequest_bits_data_lo_hi_44 = {_memRequest_bits_data_T_1605[36], _memRequest_bits_data_T_1412[36]};
  wire [3:0]       memRequest_bits_data_lo_44 = {memRequest_bits_data_lo_hi_44, memRequest_bits_data_lo_lo_44};
  wire [1:0]       memRequest_bits_data_hi_lo_44 = {_memRequest_bits_data_T_1991[36], _memRequest_bits_data_T_1798[36]};
  wire [1:0]       memRequest_bits_data_hi_hi_44 = {_memRequest_bits_data_T_2377[36], _memRequest_bits_data_T_2184[36]};
  wire [3:0]       memRequest_bits_data_hi_44 = {memRequest_bits_data_hi_hi_44, memRequest_bits_data_hi_lo_44};
  wire [1:0]       memRequest_bits_data_lo_lo_45 = {_memRequest_bits_data_T_1219[37], _memRequest_bits_data_T_1026[37]};
  wire [1:0]       memRequest_bits_data_lo_hi_45 = {_memRequest_bits_data_T_1605[37], _memRequest_bits_data_T_1412[37]};
  wire [3:0]       memRequest_bits_data_lo_45 = {memRequest_bits_data_lo_hi_45, memRequest_bits_data_lo_lo_45};
  wire [1:0]       memRequest_bits_data_hi_lo_45 = {_memRequest_bits_data_T_1991[37], _memRequest_bits_data_T_1798[37]};
  wire [1:0]       memRequest_bits_data_hi_hi_45 = {_memRequest_bits_data_T_2377[37], _memRequest_bits_data_T_2184[37]};
  wire [3:0]       memRequest_bits_data_hi_45 = {memRequest_bits_data_hi_hi_45, memRequest_bits_data_hi_lo_45};
  wire [1:0]       memRequest_bits_data_lo_lo_46 = {_memRequest_bits_data_T_1219[38], _memRequest_bits_data_T_1026[38]};
  wire [1:0]       memRequest_bits_data_lo_hi_46 = {_memRequest_bits_data_T_1605[38], _memRequest_bits_data_T_1412[38]};
  wire [3:0]       memRequest_bits_data_lo_46 = {memRequest_bits_data_lo_hi_46, memRequest_bits_data_lo_lo_46};
  wire [1:0]       memRequest_bits_data_hi_lo_46 = {_memRequest_bits_data_T_1991[38], _memRequest_bits_data_T_1798[38]};
  wire [1:0]       memRequest_bits_data_hi_hi_46 = {_memRequest_bits_data_T_2377[38], _memRequest_bits_data_T_2184[38]};
  wire [3:0]       memRequest_bits_data_hi_46 = {memRequest_bits_data_hi_hi_46, memRequest_bits_data_hi_lo_46};
  wire [1:0]       memRequest_bits_data_lo_lo_47 = {_memRequest_bits_data_T_1219[39], _memRequest_bits_data_T_1026[39]};
  wire [1:0]       memRequest_bits_data_lo_hi_47 = {_memRequest_bits_data_T_1605[39], _memRequest_bits_data_T_1412[39]};
  wire [3:0]       memRequest_bits_data_lo_47 = {memRequest_bits_data_lo_hi_47, memRequest_bits_data_lo_lo_47};
  wire [1:0]       memRequest_bits_data_hi_lo_47 = {_memRequest_bits_data_T_1991[39], _memRequest_bits_data_T_1798[39]};
  wire [1:0]       memRequest_bits_data_hi_hi_47 = {_memRequest_bits_data_T_2377[39], _memRequest_bits_data_T_2184[39]};
  wire [3:0]       memRequest_bits_data_hi_47 = {memRequest_bits_data_hi_hi_47, memRequest_bits_data_hi_lo_47};
  wire [1:0]       memRequest_bits_data_lo_lo_48 = {_memRequest_bits_data_T_1219[40], _memRequest_bits_data_T_1026[40]};
  wire [1:0]       memRequest_bits_data_lo_hi_48 = {_memRequest_bits_data_T_1605[40], _memRequest_bits_data_T_1412[40]};
  wire [3:0]       memRequest_bits_data_lo_48 = {memRequest_bits_data_lo_hi_48, memRequest_bits_data_lo_lo_48};
  wire [1:0]       memRequest_bits_data_hi_lo_48 = {_memRequest_bits_data_T_1991[40], _memRequest_bits_data_T_1798[40]};
  wire [1:0]       memRequest_bits_data_hi_hi_48 = {_memRequest_bits_data_T_2377[40], _memRequest_bits_data_T_2184[40]};
  wire [3:0]       memRequest_bits_data_hi_48 = {memRequest_bits_data_hi_hi_48, memRequest_bits_data_hi_lo_48};
  wire [1:0]       memRequest_bits_data_lo_lo_49 = {_memRequest_bits_data_T_1219[41], _memRequest_bits_data_T_1026[41]};
  wire [1:0]       memRequest_bits_data_lo_hi_49 = {_memRequest_bits_data_T_1605[41], _memRequest_bits_data_T_1412[41]};
  wire [3:0]       memRequest_bits_data_lo_49 = {memRequest_bits_data_lo_hi_49, memRequest_bits_data_lo_lo_49};
  wire [1:0]       memRequest_bits_data_hi_lo_49 = {_memRequest_bits_data_T_1991[41], _memRequest_bits_data_T_1798[41]};
  wire [1:0]       memRequest_bits_data_hi_hi_49 = {_memRequest_bits_data_T_2377[41], _memRequest_bits_data_T_2184[41]};
  wire [3:0]       memRequest_bits_data_hi_49 = {memRequest_bits_data_hi_hi_49, memRequest_bits_data_hi_lo_49};
  wire [1:0]       memRequest_bits_data_lo_lo_50 = {_memRequest_bits_data_T_1219[42], _memRequest_bits_data_T_1026[42]};
  wire [1:0]       memRequest_bits_data_lo_hi_50 = {_memRequest_bits_data_T_1605[42], _memRequest_bits_data_T_1412[42]};
  wire [3:0]       memRequest_bits_data_lo_50 = {memRequest_bits_data_lo_hi_50, memRequest_bits_data_lo_lo_50};
  wire [1:0]       memRequest_bits_data_hi_lo_50 = {_memRequest_bits_data_T_1991[42], _memRequest_bits_data_T_1798[42]};
  wire [1:0]       memRequest_bits_data_hi_hi_50 = {_memRequest_bits_data_T_2377[42], _memRequest_bits_data_T_2184[42]};
  wire [3:0]       memRequest_bits_data_hi_50 = {memRequest_bits_data_hi_hi_50, memRequest_bits_data_hi_lo_50};
  wire [1:0]       memRequest_bits_data_lo_lo_51 = {_memRequest_bits_data_T_1219[43], _memRequest_bits_data_T_1026[43]};
  wire [1:0]       memRequest_bits_data_lo_hi_51 = {_memRequest_bits_data_T_1605[43], _memRequest_bits_data_T_1412[43]};
  wire [3:0]       memRequest_bits_data_lo_51 = {memRequest_bits_data_lo_hi_51, memRequest_bits_data_lo_lo_51};
  wire [1:0]       memRequest_bits_data_hi_lo_51 = {_memRequest_bits_data_T_1991[43], _memRequest_bits_data_T_1798[43]};
  wire [1:0]       memRequest_bits_data_hi_hi_51 = {_memRequest_bits_data_T_2377[43], _memRequest_bits_data_T_2184[43]};
  wire [3:0]       memRequest_bits_data_hi_51 = {memRequest_bits_data_hi_hi_51, memRequest_bits_data_hi_lo_51};
  wire [1:0]       memRequest_bits_data_lo_lo_52 = {_memRequest_bits_data_T_1219[44], _memRequest_bits_data_T_1026[44]};
  wire [1:0]       memRequest_bits_data_lo_hi_52 = {_memRequest_bits_data_T_1605[44], _memRequest_bits_data_T_1412[44]};
  wire [3:0]       memRequest_bits_data_lo_52 = {memRequest_bits_data_lo_hi_52, memRequest_bits_data_lo_lo_52};
  wire [1:0]       memRequest_bits_data_hi_lo_52 = {_memRequest_bits_data_T_1991[44], _memRequest_bits_data_T_1798[44]};
  wire [1:0]       memRequest_bits_data_hi_hi_52 = {_memRequest_bits_data_T_2377[44], _memRequest_bits_data_T_2184[44]};
  wire [3:0]       memRequest_bits_data_hi_52 = {memRequest_bits_data_hi_hi_52, memRequest_bits_data_hi_lo_52};
  wire [1:0]       memRequest_bits_data_lo_lo_53 = {_memRequest_bits_data_T_1219[45], _memRequest_bits_data_T_1026[45]};
  wire [1:0]       memRequest_bits_data_lo_hi_53 = {_memRequest_bits_data_T_1605[45], _memRequest_bits_data_T_1412[45]};
  wire [3:0]       memRequest_bits_data_lo_53 = {memRequest_bits_data_lo_hi_53, memRequest_bits_data_lo_lo_53};
  wire [1:0]       memRequest_bits_data_hi_lo_53 = {_memRequest_bits_data_T_1991[45], _memRequest_bits_data_T_1798[45]};
  wire [1:0]       memRequest_bits_data_hi_hi_53 = {_memRequest_bits_data_T_2377[45], _memRequest_bits_data_T_2184[45]};
  wire [3:0]       memRequest_bits_data_hi_53 = {memRequest_bits_data_hi_hi_53, memRequest_bits_data_hi_lo_53};
  wire [1:0]       memRequest_bits_data_lo_lo_54 = {_memRequest_bits_data_T_1219[46], _memRequest_bits_data_T_1026[46]};
  wire [1:0]       memRequest_bits_data_lo_hi_54 = {_memRequest_bits_data_T_1605[46], _memRequest_bits_data_T_1412[46]};
  wire [3:0]       memRequest_bits_data_lo_54 = {memRequest_bits_data_lo_hi_54, memRequest_bits_data_lo_lo_54};
  wire [1:0]       memRequest_bits_data_hi_lo_54 = {_memRequest_bits_data_T_1991[46], _memRequest_bits_data_T_1798[46]};
  wire [1:0]       memRequest_bits_data_hi_hi_54 = {_memRequest_bits_data_T_2377[46], _memRequest_bits_data_T_2184[46]};
  wire [3:0]       memRequest_bits_data_hi_54 = {memRequest_bits_data_hi_hi_54, memRequest_bits_data_hi_lo_54};
  wire [1:0]       memRequest_bits_data_lo_lo_55 = {_memRequest_bits_data_T_1219[47], _memRequest_bits_data_T_1026[47]};
  wire [1:0]       memRequest_bits_data_lo_hi_55 = {_memRequest_bits_data_T_1605[47], _memRequest_bits_data_T_1412[47]};
  wire [3:0]       memRequest_bits_data_lo_55 = {memRequest_bits_data_lo_hi_55, memRequest_bits_data_lo_lo_55};
  wire [1:0]       memRequest_bits_data_hi_lo_55 = {_memRequest_bits_data_T_1991[47], _memRequest_bits_data_T_1798[47]};
  wire [1:0]       memRequest_bits_data_hi_hi_55 = {_memRequest_bits_data_T_2377[47], _memRequest_bits_data_T_2184[47]};
  wire [3:0]       memRequest_bits_data_hi_55 = {memRequest_bits_data_hi_hi_55, memRequest_bits_data_hi_lo_55};
  wire [1:0]       memRequest_bits_data_lo_lo_56 = {_memRequest_bits_data_T_1219[48], _memRequest_bits_data_T_1026[48]};
  wire [1:0]       memRequest_bits_data_lo_hi_56 = {_memRequest_bits_data_T_1605[48], _memRequest_bits_data_T_1412[48]};
  wire [3:0]       memRequest_bits_data_lo_56 = {memRequest_bits_data_lo_hi_56, memRequest_bits_data_lo_lo_56};
  wire [1:0]       memRequest_bits_data_hi_lo_56 = {_memRequest_bits_data_T_1991[48], _memRequest_bits_data_T_1798[48]};
  wire [1:0]       memRequest_bits_data_hi_hi_56 = {_memRequest_bits_data_T_2377[48], _memRequest_bits_data_T_2184[48]};
  wire [3:0]       memRequest_bits_data_hi_56 = {memRequest_bits_data_hi_hi_56, memRequest_bits_data_hi_lo_56};
  wire [1:0]       memRequest_bits_data_lo_lo_57 = {_memRequest_bits_data_T_1219[49], _memRequest_bits_data_T_1026[49]};
  wire [1:0]       memRequest_bits_data_lo_hi_57 = {_memRequest_bits_data_T_1605[49], _memRequest_bits_data_T_1412[49]};
  wire [3:0]       memRequest_bits_data_lo_57 = {memRequest_bits_data_lo_hi_57, memRequest_bits_data_lo_lo_57};
  wire [1:0]       memRequest_bits_data_hi_lo_57 = {_memRequest_bits_data_T_1991[49], _memRequest_bits_data_T_1798[49]};
  wire [1:0]       memRequest_bits_data_hi_hi_57 = {_memRequest_bits_data_T_2377[49], _memRequest_bits_data_T_2184[49]};
  wire [3:0]       memRequest_bits_data_hi_57 = {memRequest_bits_data_hi_hi_57, memRequest_bits_data_hi_lo_57};
  wire [1:0]       memRequest_bits_data_lo_lo_58 = {_memRequest_bits_data_T_1219[50], _memRequest_bits_data_T_1026[50]};
  wire [1:0]       memRequest_bits_data_lo_hi_58 = {_memRequest_bits_data_T_1605[50], _memRequest_bits_data_T_1412[50]};
  wire [3:0]       memRequest_bits_data_lo_58 = {memRequest_bits_data_lo_hi_58, memRequest_bits_data_lo_lo_58};
  wire [1:0]       memRequest_bits_data_hi_lo_58 = {_memRequest_bits_data_T_1991[50], _memRequest_bits_data_T_1798[50]};
  wire [1:0]       memRequest_bits_data_hi_hi_58 = {_memRequest_bits_data_T_2377[50], _memRequest_bits_data_T_2184[50]};
  wire [3:0]       memRequest_bits_data_hi_58 = {memRequest_bits_data_hi_hi_58, memRequest_bits_data_hi_lo_58};
  wire [1:0]       memRequest_bits_data_lo_lo_59 = {_memRequest_bits_data_T_1219[51], _memRequest_bits_data_T_1026[51]};
  wire [1:0]       memRequest_bits_data_lo_hi_59 = {_memRequest_bits_data_T_1605[51], _memRequest_bits_data_T_1412[51]};
  wire [3:0]       memRequest_bits_data_lo_59 = {memRequest_bits_data_lo_hi_59, memRequest_bits_data_lo_lo_59};
  wire [1:0]       memRequest_bits_data_hi_lo_59 = {_memRequest_bits_data_T_1991[51], _memRequest_bits_data_T_1798[51]};
  wire [1:0]       memRequest_bits_data_hi_hi_59 = {_memRequest_bits_data_T_2377[51], _memRequest_bits_data_T_2184[51]};
  wire [3:0]       memRequest_bits_data_hi_59 = {memRequest_bits_data_hi_hi_59, memRequest_bits_data_hi_lo_59};
  wire [1:0]       memRequest_bits_data_lo_lo_60 = {_memRequest_bits_data_T_1219[52], _memRequest_bits_data_T_1026[52]};
  wire [1:0]       memRequest_bits_data_lo_hi_60 = {_memRequest_bits_data_T_1605[52], _memRequest_bits_data_T_1412[52]};
  wire [3:0]       memRequest_bits_data_lo_60 = {memRequest_bits_data_lo_hi_60, memRequest_bits_data_lo_lo_60};
  wire [1:0]       memRequest_bits_data_hi_lo_60 = {_memRequest_bits_data_T_1991[52], _memRequest_bits_data_T_1798[52]};
  wire [1:0]       memRequest_bits_data_hi_hi_60 = {_memRequest_bits_data_T_2377[52], _memRequest_bits_data_T_2184[52]};
  wire [3:0]       memRequest_bits_data_hi_60 = {memRequest_bits_data_hi_hi_60, memRequest_bits_data_hi_lo_60};
  wire [1:0]       memRequest_bits_data_lo_lo_61 = {_memRequest_bits_data_T_1219[53], _memRequest_bits_data_T_1026[53]};
  wire [1:0]       memRequest_bits_data_lo_hi_61 = {_memRequest_bits_data_T_1605[53], _memRequest_bits_data_T_1412[53]};
  wire [3:0]       memRequest_bits_data_lo_61 = {memRequest_bits_data_lo_hi_61, memRequest_bits_data_lo_lo_61};
  wire [1:0]       memRequest_bits_data_hi_lo_61 = {_memRequest_bits_data_T_1991[53], _memRequest_bits_data_T_1798[53]};
  wire [1:0]       memRequest_bits_data_hi_hi_61 = {_memRequest_bits_data_T_2377[53], _memRequest_bits_data_T_2184[53]};
  wire [3:0]       memRequest_bits_data_hi_61 = {memRequest_bits_data_hi_hi_61, memRequest_bits_data_hi_lo_61};
  wire [1:0]       memRequest_bits_data_lo_lo_62 = {_memRequest_bits_data_T_1219[54], _memRequest_bits_data_T_1026[54]};
  wire [1:0]       memRequest_bits_data_lo_hi_62 = {_memRequest_bits_data_T_1605[54], _memRequest_bits_data_T_1412[54]};
  wire [3:0]       memRequest_bits_data_lo_62 = {memRequest_bits_data_lo_hi_62, memRequest_bits_data_lo_lo_62};
  wire [1:0]       memRequest_bits_data_hi_lo_62 = {_memRequest_bits_data_T_1991[54], _memRequest_bits_data_T_1798[54]};
  wire [1:0]       memRequest_bits_data_hi_hi_62 = {_memRequest_bits_data_T_2377[54], _memRequest_bits_data_T_2184[54]};
  wire [3:0]       memRequest_bits_data_hi_62 = {memRequest_bits_data_hi_hi_62, memRequest_bits_data_hi_lo_62};
  wire [1:0]       memRequest_bits_data_lo_lo_63 = {_memRequest_bits_data_T_1219[55], _memRequest_bits_data_T_1026[55]};
  wire [1:0]       memRequest_bits_data_lo_hi_63 = {_memRequest_bits_data_T_1605[55], _memRequest_bits_data_T_1412[55]};
  wire [3:0]       memRequest_bits_data_lo_63 = {memRequest_bits_data_lo_hi_63, memRequest_bits_data_lo_lo_63};
  wire [1:0]       memRequest_bits_data_hi_lo_63 = {_memRequest_bits_data_T_1991[55], _memRequest_bits_data_T_1798[55]};
  wire [1:0]       memRequest_bits_data_hi_hi_63 = {_memRequest_bits_data_T_2377[55], _memRequest_bits_data_T_2184[55]};
  wire [3:0]       memRequest_bits_data_hi_63 = {memRequest_bits_data_hi_hi_63, memRequest_bits_data_hi_lo_63};
  wire [1:0]       memRequest_bits_data_lo_lo_64 = {_memRequest_bits_data_T_1219[56], _memRequest_bits_data_T_1026[56]};
  wire [1:0]       memRequest_bits_data_lo_hi_64 = {_memRequest_bits_data_T_1605[56], _memRequest_bits_data_T_1412[56]};
  wire [3:0]       memRequest_bits_data_lo_64 = {memRequest_bits_data_lo_hi_64, memRequest_bits_data_lo_lo_64};
  wire [1:0]       memRequest_bits_data_hi_lo_64 = {_memRequest_bits_data_T_1991[56], _memRequest_bits_data_T_1798[56]};
  wire [1:0]       memRequest_bits_data_hi_hi_64 = {_memRequest_bits_data_T_2377[56], _memRequest_bits_data_T_2184[56]};
  wire [3:0]       memRequest_bits_data_hi_64 = {memRequest_bits_data_hi_hi_64, memRequest_bits_data_hi_lo_64};
  wire [1:0]       memRequest_bits_data_lo_lo_65 = {_memRequest_bits_data_T_1219[57], _memRequest_bits_data_T_1026[57]};
  wire [1:0]       memRequest_bits_data_lo_hi_65 = {_memRequest_bits_data_T_1605[57], _memRequest_bits_data_T_1412[57]};
  wire [3:0]       memRequest_bits_data_lo_65 = {memRequest_bits_data_lo_hi_65, memRequest_bits_data_lo_lo_65};
  wire [1:0]       memRequest_bits_data_hi_lo_65 = {_memRequest_bits_data_T_1991[57], _memRequest_bits_data_T_1798[57]};
  wire [1:0]       memRequest_bits_data_hi_hi_65 = {_memRequest_bits_data_T_2377[57], _memRequest_bits_data_T_2184[57]};
  wire [3:0]       memRequest_bits_data_hi_65 = {memRequest_bits_data_hi_hi_65, memRequest_bits_data_hi_lo_65};
  wire [1:0]       memRequest_bits_data_lo_lo_66 = {_memRequest_bits_data_T_1219[58], _memRequest_bits_data_T_1026[58]};
  wire [1:0]       memRequest_bits_data_lo_hi_66 = {_memRequest_bits_data_T_1605[58], _memRequest_bits_data_T_1412[58]};
  wire [3:0]       memRequest_bits_data_lo_66 = {memRequest_bits_data_lo_hi_66, memRequest_bits_data_lo_lo_66};
  wire [1:0]       memRequest_bits_data_hi_lo_66 = {_memRequest_bits_data_T_1991[58], _memRequest_bits_data_T_1798[58]};
  wire [1:0]       memRequest_bits_data_hi_hi_66 = {_memRequest_bits_data_T_2377[58], _memRequest_bits_data_T_2184[58]};
  wire [3:0]       memRequest_bits_data_hi_66 = {memRequest_bits_data_hi_hi_66, memRequest_bits_data_hi_lo_66};
  wire [1:0]       memRequest_bits_data_lo_lo_67 = {_memRequest_bits_data_T_1219[59], _memRequest_bits_data_T_1026[59]};
  wire [1:0]       memRequest_bits_data_lo_hi_67 = {_memRequest_bits_data_T_1605[59], _memRequest_bits_data_T_1412[59]};
  wire [3:0]       memRequest_bits_data_lo_67 = {memRequest_bits_data_lo_hi_67, memRequest_bits_data_lo_lo_67};
  wire [1:0]       memRequest_bits_data_hi_lo_67 = {_memRequest_bits_data_T_1991[59], _memRequest_bits_data_T_1798[59]};
  wire [1:0]       memRequest_bits_data_hi_hi_67 = {_memRequest_bits_data_T_2377[59], _memRequest_bits_data_T_2184[59]};
  wire [3:0]       memRequest_bits_data_hi_67 = {memRequest_bits_data_hi_hi_67, memRequest_bits_data_hi_lo_67};
  wire [1:0]       memRequest_bits_data_lo_lo_68 = {_memRequest_bits_data_T_1219[60], _memRequest_bits_data_T_1026[60]};
  wire [1:0]       memRequest_bits_data_lo_hi_68 = {_memRequest_bits_data_T_1605[60], _memRequest_bits_data_T_1412[60]};
  wire [3:0]       memRequest_bits_data_lo_68 = {memRequest_bits_data_lo_hi_68, memRequest_bits_data_lo_lo_68};
  wire [1:0]       memRequest_bits_data_hi_lo_68 = {_memRequest_bits_data_T_1991[60], _memRequest_bits_data_T_1798[60]};
  wire [1:0]       memRequest_bits_data_hi_hi_68 = {_memRequest_bits_data_T_2377[60], _memRequest_bits_data_T_2184[60]};
  wire [3:0]       memRequest_bits_data_hi_68 = {memRequest_bits_data_hi_hi_68, memRequest_bits_data_hi_lo_68};
  wire [1:0]       memRequest_bits_data_lo_lo_69 = {_memRequest_bits_data_T_1219[61], _memRequest_bits_data_T_1026[61]};
  wire [1:0]       memRequest_bits_data_lo_hi_69 = {_memRequest_bits_data_T_1605[61], _memRequest_bits_data_T_1412[61]};
  wire [3:0]       memRequest_bits_data_lo_69 = {memRequest_bits_data_lo_hi_69, memRequest_bits_data_lo_lo_69};
  wire [1:0]       memRequest_bits_data_hi_lo_69 = {_memRequest_bits_data_T_1991[61], _memRequest_bits_data_T_1798[61]};
  wire [1:0]       memRequest_bits_data_hi_hi_69 = {_memRequest_bits_data_T_2377[61], _memRequest_bits_data_T_2184[61]};
  wire [3:0]       memRequest_bits_data_hi_69 = {memRequest_bits_data_hi_hi_69, memRequest_bits_data_hi_lo_69};
  wire [1:0]       memRequest_bits_data_lo_lo_70 = {_memRequest_bits_data_T_1219[62], _memRequest_bits_data_T_1026[62]};
  wire [1:0]       memRequest_bits_data_lo_hi_70 = {_memRequest_bits_data_T_1605[62], _memRequest_bits_data_T_1412[62]};
  wire [3:0]       memRequest_bits_data_lo_70 = {memRequest_bits_data_lo_hi_70, memRequest_bits_data_lo_lo_70};
  wire [1:0]       memRequest_bits_data_hi_lo_70 = {_memRequest_bits_data_T_1991[62], _memRequest_bits_data_T_1798[62]};
  wire [1:0]       memRequest_bits_data_hi_hi_70 = {_memRequest_bits_data_T_2377[62], _memRequest_bits_data_T_2184[62]};
  wire [3:0]       memRequest_bits_data_hi_70 = {memRequest_bits_data_hi_hi_70, memRequest_bits_data_hi_lo_70};
  wire [1:0]       memRequest_bits_data_lo_lo_71 = {_memRequest_bits_data_T_1219[63], _memRequest_bits_data_T_1026[63]};
  wire [1:0]       memRequest_bits_data_lo_hi_71 = {_memRequest_bits_data_T_1605[63], _memRequest_bits_data_T_1412[63]};
  wire [3:0]       memRequest_bits_data_lo_71 = {memRequest_bits_data_lo_hi_71, memRequest_bits_data_lo_lo_71};
  wire [1:0]       memRequest_bits_data_hi_lo_71 = {_memRequest_bits_data_T_1991[63], _memRequest_bits_data_T_1798[63]};
  wire [1:0]       memRequest_bits_data_hi_hi_71 = {_memRequest_bits_data_T_2377[63], _memRequest_bits_data_T_2184[63]};
  wire [3:0]       memRequest_bits_data_hi_71 = {memRequest_bits_data_hi_hi_71, memRequest_bits_data_hi_lo_71};
  wire [1:0]       memRequest_bits_data_lo_lo_72 = {_memRequest_bits_data_T_1219[64], _memRequest_bits_data_T_1026[64]};
  wire [1:0]       memRequest_bits_data_lo_hi_72 = {_memRequest_bits_data_T_1605[64], _memRequest_bits_data_T_1412[64]};
  wire [3:0]       memRequest_bits_data_lo_72 = {memRequest_bits_data_lo_hi_72, memRequest_bits_data_lo_lo_72};
  wire [1:0]       memRequest_bits_data_hi_lo_72 = {_memRequest_bits_data_T_1991[64], _memRequest_bits_data_T_1798[64]};
  wire [1:0]       memRequest_bits_data_hi_hi_72 = {_memRequest_bits_data_T_2377[64], _memRequest_bits_data_T_2184[64]};
  wire [3:0]       memRequest_bits_data_hi_72 = {memRequest_bits_data_hi_hi_72, memRequest_bits_data_hi_lo_72};
  wire [1:0]       memRequest_bits_data_lo_lo_73 = {_memRequest_bits_data_T_1219[65], _memRequest_bits_data_T_1026[65]};
  wire [1:0]       memRequest_bits_data_lo_hi_73 = {_memRequest_bits_data_T_1605[65], _memRequest_bits_data_T_1412[65]};
  wire [3:0]       memRequest_bits_data_lo_73 = {memRequest_bits_data_lo_hi_73, memRequest_bits_data_lo_lo_73};
  wire [1:0]       memRequest_bits_data_hi_lo_73 = {_memRequest_bits_data_T_1991[65], _memRequest_bits_data_T_1798[65]};
  wire [1:0]       memRequest_bits_data_hi_hi_73 = {_memRequest_bits_data_T_2377[65], _memRequest_bits_data_T_2184[65]};
  wire [3:0]       memRequest_bits_data_hi_73 = {memRequest_bits_data_hi_hi_73, memRequest_bits_data_hi_lo_73};
  wire [1:0]       memRequest_bits_data_lo_lo_74 = {_memRequest_bits_data_T_1219[66], _memRequest_bits_data_T_1026[66]};
  wire [1:0]       memRequest_bits_data_lo_hi_74 = {_memRequest_bits_data_T_1605[66], _memRequest_bits_data_T_1412[66]};
  wire [3:0]       memRequest_bits_data_lo_74 = {memRequest_bits_data_lo_hi_74, memRequest_bits_data_lo_lo_74};
  wire [1:0]       memRequest_bits_data_hi_lo_74 = {_memRequest_bits_data_T_1991[66], _memRequest_bits_data_T_1798[66]};
  wire [1:0]       memRequest_bits_data_hi_hi_74 = {_memRequest_bits_data_T_2377[66], _memRequest_bits_data_T_2184[66]};
  wire [3:0]       memRequest_bits_data_hi_74 = {memRequest_bits_data_hi_hi_74, memRequest_bits_data_hi_lo_74};
  wire [1:0]       memRequest_bits_data_lo_lo_75 = {_memRequest_bits_data_T_1219[67], _memRequest_bits_data_T_1026[67]};
  wire [1:0]       memRequest_bits_data_lo_hi_75 = {_memRequest_bits_data_T_1605[67], _memRequest_bits_data_T_1412[67]};
  wire [3:0]       memRequest_bits_data_lo_75 = {memRequest_bits_data_lo_hi_75, memRequest_bits_data_lo_lo_75};
  wire [1:0]       memRequest_bits_data_hi_lo_75 = {_memRequest_bits_data_T_1991[67], _memRequest_bits_data_T_1798[67]};
  wire [1:0]       memRequest_bits_data_hi_hi_75 = {_memRequest_bits_data_T_2377[67], _memRequest_bits_data_T_2184[67]};
  wire [3:0]       memRequest_bits_data_hi_75 = {memRequest_bits_data_hi_hi_75, memRequest_bits_data_hi_lo_75};
  wire [1:0]       memRequest_bits_data_lo_lo_76 = {_memRequest_bits_data_T_1219[68], _memRequest_bits_data_T_1026[68]};
  wire [1:0]       memRequest_bits_data_lo_hi_76 = {_memRequest_bits_data_T_1605[68], _memRequest_bits_data_T_1412[68]};
  wire [3:0]       memRequest_bits_data_lo_76 = {memRequest_bits_data_lo_hi_76, memRequest_bits_data_lo_lo_76};
  wire [1:0]       memRequest_bits_data_hi_lo_76 = {_memRequest_bits_data_T_1991[68], _memRequest_bits_data_T_1798[68]};
  wire [1:0]       memRequest_bits_data_hi_hi_76 = {_memRequest_bits_data_T_2377[68], _memRequest_bits_data_T_2184[68]};
  wire [3:0]       memRequest_bits_data_hi_76 = {memRequest_bits_data_hi_hi_76, memRequest_bits_data_hi_lo_76};
  wire [1:0]       memRequest_bits_data_lo_lo_77 = {_memRequest_bits_data_T_1219[69], _memRequest_bits_data_T_1026[69]};
  wire [1:0]       memRequest_bits_data_lo_hi_77 = {_memRequest_bits_data_T_1605[69], _memRequest_bits_data_T_1412[69]};
  wire [3:0]       memRequest_bits_data_lo_77 = {memRequest_bits_data_lo_hi_77, memRequest_bits_data_lo_lo_77};
  wire [1:0]       memRequest_bits_data_hi_lo_77 = {_memRequest_bits_data_T_1991[69], _memRequest_bits_data_T_1798[69]};
  wire [1:0]       memRequest_bits_data_hi_hi_77 = {_memRequest_bits_data_T_2377[69], _memRequest_bits_data_T_2184[69]};
  wire [3:0]       memRequest_bits_data_hi_77 = {memRequest_bits_data_hi_hi_77, memRequest_bits_data_hi_lo_77};
  wire [1:0]       memRequest_bits_data_lo_lo_78 = {_memRequest_bits_data_T_1219[70], _memRequest_bits_data_T_1026[70]};
  wire [1:0]       memRequest_bits_data_lo_hi_78 = {_memRequest_bits_data_T_1605[70], _memRequest_bits_data_T_1412[70]};
  wire [3:0]       memRequest_bits_data_lo_78 = {memRequest_bits_data_lo_hi_78, memRequest_bits_data_lo_lo_78};
  wire [1:0]       memRequest_bits_data_hi_lo_78 = {_memRequest_bits_data_T_1991[70], _memRequest_bits_data_T_1798[70]};
  wire [1:0]       memRequest_bits_data_hi_hi_78 = {_memRequest_bits_data_T_2377[70], _memRequest_bits_data_T_2184[70]};
  wire [3:0]       memRequest_bits_data_hi_78 = {memRequest_bits_data_hi_hi_78, memRequest_bits_data_hi_lo_78};
  wire [1:0]       memRequest_bits_data_lo_lo_79 = {_memRequest_bits_data_T_1219[71], _memRequest_bits_data_T_1026[71]};
  wire [1:0]       memRequest_bits_data_lo_hi_79 = {_memRequest_bits_data_T_1605[71], _memRequest_bits_data_T_1412[71]};
  wire [3:0]       memRequest_bits_data_lo_79 = {memRequest_bits_data_lo_hi_79, memRequest_bits_data_lo_lo_79};
  wire [1:0]       memRequest_bits_data_hi_lo_79 = {_memRequest_bits_data_T_1991[71], _memRequest_bits_data_T_1798[71]};
  wire [1:0]       memRequest_bits_data_hi_hi_79 = {_memRequest_bits_data_T_2377[71], _memRequest_bits_data_T_2184[71]};
  wire [3:0]       memRequest_bits_data_hi_79 = {memRequest_bits_data_hi_hi_79, memRequest_bits_data_hi_lo_79};
  wire [1:0]       memRequest_bits_data_lo_lo_80 = {_memRequest_bits_data_T_1219[72], _memRequest_bits_data_T_1026[72]};
  wire [1:0]       memRequest_bits_data_lo_hi_80 = {_memRequest_bits_data_T_1605[72], _memRequest_bits_data_T_1412[72]};
  wire [3:0]       memRequest_bits_data_lo_80 = {memRequest_bits_data_lo_hi_80, memRequest_bits_data_lo_lo_80};
  wire [1:0]       memRequest_bits_data_hi_lo_80 = {_memRequest_bits_data_T_1991[72], _memRequest_bits_data_T_1798[72]};
  wire [1:0]       memRequest_bits_data_hi_hi_80 = {_memRequest_bits_data_T_2377[72], _memRequest_bits_data_T_2184[72]};
  wire [3:0]       memRequest_bits_data_hi_80 = {memRequest_bits_data_hi_hi_80, memRequest_bits_data_hi_lo_80};
  wire [1:0]       memRequest_bits_data_lo_lo_81 = {_memRequest_bits_data_T_1219[73], _memRequest_bits_data_T_1026[73]};
  wire [1:0]       memRequest_bits_data_lo_hi_81 = {_memRequest_bits_data_T_1605[73], _memRequest_bits_data_T_1412[73]};
  wire [3:0]       memRequest_bits_data_lo_81 = {memRequest_bits_data_lo_hi_81, memRequest_bits_data_lo_lo_81};
  wire [1:0]       memRequest_bits_data_hi_lo_81 = {_memRequest_bits_data_T_1991[73], _memRequest_bits_data_T_1798[73]};
  wire [1:0]       memRequest_bits_data_hi_hi_81 = {_memRequest_bits_data_T_2377[73], _memRequest_bits_data_T_2184[73]};
  wire [3:0]       memRequest_bits_data_hi_81 = {memRequest_bits_data_hi_hi_81, memRequest_bits_data_hi_lo_81};
  wire [1:0]       memRequest_bits_data_lo_lo_82 = {_memRequest_bits_data_T_1219[74], _memRequest_bits_data_T_1026[74]};
  wire [1:0]       memRequest_bits_data_lo_hi_82 = {_memRequest_bits_data_T_1605[74], _memRequest_bits_data_T_1412[74]};
  wire [3:0]       memRequest_bits_data_lo_82 = {memRequest_bits_data_lo_hi_82, memRequest_bits_data_lo_lo_82};
  wire [1:0]       memRequest_bits_data_hi_lo_82 = {_memRequest_bits_data_T_1991[74], _memRequest_bits_data_T_1798[74]};
  wire [1:0]       memRequest_bits_data_hi_hi_82 = {_memRequest_bits_data_T_2377[74], _memRequest_bits_data_T_2184[74]};
  wire [3:0]       memRequest_bits_data_hi_82 = {memRequest_bits_data_hi_hi_82, memRequest_bits_data_hi_lo_82};
  wire [1:0]       memRequest_bits_data_lo_lo_83 = {_memRequest_bits_data_T_1219[75], _memRequest_bits_data_T_1026[75]};
  wire [1:0]       memRequest_bits_data_lo_hi_83 = {_memRequest_bits_data_T_1605[75], _memRequest_bits_data_T_1412[75]};
  wire [3:0]       memRequest_bits_data_lo_83 = {memRequest_bits_data_lo_hi_83, memRequest_bits_data_lo_lo_83};
  wire [1:0]       memRequest_bits_data_hi_lo_83 = {_memRequest_bits_data_T_1991[75], _memRequest_bits_data_T_1798[75]};
  wire [1:0]       memRequest_bits_data_hi_hi_83 = {_memRequest_bits_data_T_2377[75], _memRequest_bits_data_T_2184[75]};
  wire [3:0]       memRequest_bits_data_hi_83 = {memRequest_bits_data_hi_hi_83, memRequest_bits_data_hi_lo_83};
  wire [1:0]       memRequest_bits_data_lo_lo_84 = {_memRequest_bits_data_T_1219[76], _memRequest_bits_data_T_1026[76]};
  wire [1:0]       memRequest_bits_data_lo_hi_84 = {_memRequest_bits_data_T_1605[76], _memRequest_bits_data_T_1412[76]};
  wire [3:0]       memRequest_bits_data_lo_84 = {memRequest_bits_data_lo_hi_84, memRequest_bits_data_lo_lo_84};
  wire [1:0]       memRequest_bits_data_hi_lo_84 = {_memRequest_bits_data_T_1991[76], _memRequest_bits_data_T_1798[76]};
  wire [1:0]       memRequest_bits_data_hi_hi_84 = {_memRequest_bits_data_T_2377[76], _memRequest_bits_data_T_2184[76]};
  wire [3:0]       memRequest_bits_data_hi_84 = {memRequest_bits_data_hi_hi_84, memRequest_bits_data_hi_lo_84};
  wire [1:0]       memRequest_bits_data_lo_lo_85 = {_memRequest_bits_data_T_1219[77], _memRequest_bits_data_T_1026[77]};
  wire [1:0]       memRequest_bits_data_lo_hi_85 = {_memRequest_bits_data_T_1605[77], _memRequest_bits_data_T_1412[77]};
  wire [3:0]       memRequest_bits_data_lo_85 = {memRequest_bits_data_lo_hi_85, memRequest_bits_data_lo_lo_85};
  wire [1:0]       memRequest_bits_data_hi_lo_85 = {_memRequest_bits_data_T_1991[77], _memRequest_bits_data_T_1798[77]};
  wire [1:0]       memRequest_bits_data_hi_hi_85 = {_memRequest_bits_data_T_2377[77], _memRequest_bits_data_T_2184[77]};
  wire [3:0]       memRequest_bits_data_hi_85 = {memRequest_bits_data_hi_hi_85, memRequest_bits_data_hi_lo_85};
  wire [1:0]       memRequest_bits_data_lo_lo_86 = {_memRequest_bits_data_T_1219[78], _memRequest_bits_data_T_1026[78]};
  wire [1:0]       memRequest_bits_data_lo_hi_86 = {_memRequest_bits_data_T_1605[78], _memRequest_bits_data_T_1412[78]};
  wire [3:0]       memRequest_bits_data_lo_86 = {memRequest_bits_data_lo_hi_86, memRequest_bits_data_lo_lo_86};
  wire [1:0]       memRequest_bits_data_hi_lo_86 = {_memRequest_bits_data_T_1991[78], _memRequest_bits_data_T_1798[78]};
  wire [1:0]       memRequest_bits_data_hi_hi_86 = {_memRequest_bits_data_T_2377[78], _memRequest_bits_data_T_2184[78]};
  wire [3:0]       memRequest_bits_data_hi_86 = {memRequest_bits_data_hi_hi_86, memRequest_bits_data_hi_lo_86};
  wire [1:0]       memRequest_bits_data_lo_lo_87 = {_memRequest_bits_data_T_1219[79], _memRequest_bits_data_T_1026[79]};
  wire [1:0]       memRequest_bits_data_lo_hi_87 = {_memRequest_bits_data_T_1605[79], _memRequest_bits_data_T_1412[79]};
  wire [3:0]       memRequest_bits_data_lo_87 = {memRequest_bits_data_lo_hi_87, memRequest_bits_data_lo_lo_87};
  wire [1:0]       memRequest_bits_data_hi_lo_87 = {_memRequest_bits_data_T_1991[79], _memRequest_bits_data_T_1798[79]};
  wire [1:0]       memRequest_bits_data_hi_hi_87 = {_memRequest_bits_data_T_2377[79], _memRequest_bits_data_T_2184[79]};
  wire [3:0]       memRequest_bits_data_hi_87 = {memRequest_bits_data_hi_hi_87, memRequest_bits_data_hi_lo_87};
  wire [1:0]       memRequest_bits_data_lo_lo_88 = {_memRequest_bits_data_T_1219[80], _memRequest_bits_data_T_1026[80]};
  wire [1:0]       memRequest_bits_data_lo_hi_88 = {_memRequest_bits_data_T_1605[80], _memRequest_bits_data_T_1412[80]};
  wire [3:0]       memRequest_bits_data_lo_88 = {memRequest_bits_data_lo_hi_88, memRequest_bits_data_lo_lo_88};
  wire [1:0]       memRequest_bits_data_hi_lo_88 = {_memRequest_bits_data_T_1991[80], _memRequest_bits_data_T_1798[80]};
  wire [1:0]       memRequest_bits_data_hi_hi_88 = {_memRequest_bits_data_T_2377[80], _memRequest_bits_data_T_2184[80]};
  wire [3:0]       memRequest_bits_data_hi_88 = {memRequest_bits_data_hi_hi_88, memRequest_bits_data_hi_lo_88};
  wire [1:0]       memRequest_bits_data_lo_lo_89 = {_memRequest_bits_data_T_1219[81], _memRequest_bits_data_T_1026[81]};
  wire [1:0]       memRequest_bits_data_lo_hi_89 = {_memRequest_bits_data_T_1605[81], _memRequest_bits_data_T_1412[81]};
  wire [3:0]       memRequest_bits_data_lo_89 = {memRequest_bits_data_lo_hi_89, memRequest_bits_data_lo_lo_89};
  wire [1:0]       memRequest_bits_data_hi_lo_89 = {_memRequest_bits_data_T_1991[81], _memRequest_bits_data_T_1798[81]};
  wire [1:0]       memRequest_bits_data_hi_hi_89 = {_memRequest_bits_data_T_2377[81], _memRequest_bits_data_T_2184[81]};
  wire [3:0]       memRequest_bits_data_hi_89 = {memRequest_bits_data_hi_hi_89, memRequest_bits_data_hi_lo_89};
  wire [1:0]       memRequest_bits_data_lo_lo_90 = {_memRequest_bits_data_T_1219[82], _memRequest_bits_data_T_1026[82]};
  wire [1:0]       memRequest_bits_data_lo_hi_90 = {_memRequest_bits_data_T_1605[82], _memRequest_bits_data_T_1412[82]};
  wire [3:0]       memRequest_bits_data_lo_90 = {memRequest_bits_data_lo_hi_90, memRequest_bits_data_lo_lo_90};
  wire [1:0]       memRequest_bits_data_hi_lo_90 = {_memRequest_bits_data_T_1991[82], _memRequest_bits_data_T_1798[82]};
  wire [1:0]       memRequest_bits_data_hi_hi_90 = {_memRequest_bits_data_T_2377[82], _memRequest_bits_data_T_2184[82]};
  wire [3:0]       memRequest_bits_data_hi_90 = {memRequest_bits_data_hi_hi_90, memRequest_bits_data_hi_lo_90};
  wire [1:0]       memRequest_bits_data_lo_lo_91 = {_memRequest_bits_data_T_1219[83], _memRequest_bits_data_T_1026[83]};
  wire [1:0]       memRequest_bits_data_lo_hi_91 = {_memRequest_bits_data_T_1605[83], _memRequest_bits_data_T_1412[83]};
  wire [3:0]       memRequest_bits_data_lo_91 = {memRequest_bits_data_lo_hi_91, memRequest_bits_data_lo_lo_91};
  wire [1:0]       memRequest_bits_data_hi_lo_91 = {_memRequest_bits_data_T_1991[83], _memRequest_bits_data_T_1798[83]};
  wire [1:0]       memRequest_bits_data_hi_hi_91 = {_memRequest_bits_data_T_2377[83], _memRequest_bits_data_T_2184[83]};
  wire [3:0]       memRequest_bits_data_hi_91 = {memRequest_bits_data_hi_hi_91, memRequest_bits_data_hi_lo_91};
  wire [1:0]       memRequest_bits_data_lo_lo_92 = {_memRequest_bits_data_T_1219[84], _memRequest_bits_data_T_1026[84]};
  wire [1:0]       memRequest_bits_data_lo_hi_92 = {_memRequest_bits_data_T_1605[84], _memRequest_bits_data_T_1412[84]};
  wire [3:0]       memRequest_bits_data_lo_92 = {memRequest_bits_data_lo_hi_92, memRequest_bits_data_lo_lo_92};
  wire [1:0]       memRequest_bits_data_hi_lo_92 = {_memRequest_bits_data_T_1991[84], _memRequest_bits_data_T_1798[84]};
  wire [1:0]       memRequest_bits_data_hi_hi_92 = {_memRequest_bits_data_T_2377[84], _memRequest_bits_data_T_2184[84]};
  wire [3:0]       memRequest_bits_data_hi_92 = {memRequest_bits_data_hi_hi_92, memRequest_bits_data_hi_lo_92};
  wire [1:0]       memRequest_bits_data_lo_lo_93 = {_memRequest_bits_data_T_1219[85], _memRequest_bits_data_T_1026[85]};
  wire [1:0]       memRequest_bits_data_lo_hi_93 = {_memRequest_bits_data_T_1605[85], _memRequest_bits_data_T_1412[85]};
  wire [3:0]       memRequest_bits_data_lo_93 = {memRequest_bits_data_lo_hi_93, memRequest_bits_data_lo_lo_93};
  wire [1:0]       memRequest_bits_data_hi_lo_93 = {_memRequest_bits_data_T_1991[85], _memRequest_bits_data_T_1798[85]};
  wire [1:0]       memRequest_bits_data_hi_hi_93 = {_memRequest_bits_data_T_2377[85], _memRequest_bits_data_T_2184[85]};
  wire [3:0]       memRequest_bits_data_hi_93 = {memRequest_bits_data_hi_hi_93, memRequest_bits_data_hi_lo_93};
  wire [1:0]       memRequest_bits_data_lo_lo_94 = {_memRequest_bits_data_T_1219[86], _memRequest_bits_data_T_1026[86]};
  wire [1:0]       memRequest_bits_data_lo_hi_94 = {_memRequest_bits_data_T_1605[86], _memRequest_bits_data_T_1412[86]};
  wire [3:0]       memRequest_bits_data_lo_94 = {memRequest_bits_data_lo_hi_94, memRequest_bits_data_lo_lo_94};
  wire [1:0]       memRequest_bits_data_hi_lo_94 = {_memRequest_bits_data_T_1991[86], _memRequest_bits_data_T_1798[86]};
  wire [1:0]       memRequest_bits_data_hi_hi_94 = {_memRequest_bits_data_T_2377[86], _memRequest_bits_data_T_2184[86]};
  wire [3:0]       memRequest_bits_data_hi_94 = {memRequest_bits_data_hi_hi_94, memRequest_bits_data_hi_lo_94};
  wire [1:0]       memRequest_bits_data_lo_lo_95 = {_memRequest_bits_data_T_1219[87], _memRequest_bits_data_T_1026[87]};
  wire [1:0]       memRequest_bits_data_lo_hi_95 = {_memRequest_bits_data_T_1605[87], _memRequest_bits_data_T_1412[87]};
  wire [3:0]       memRequest_bits_data_lo_95 = {memRequest_bits_data_lo_hi_95, memRequest_bits_data_lo_lo_95};
  wire [1:0]       memRequest_bits_data_hi_lo_95 = {_memRequest_bits_data_T_1991[87], _memRequest_bits_data_T_1798[87]};
  wire [1:0]       memRequest_bits_data_hi_hi_95 = {_memRequest_bits_data_T_2377[87], _memRequest_bits_data_T_2184[87]};
  wire [3:0]       memRequest_bits_data_hi_95 = {memRequest_bits_data_hi_hi_95, memRequest_bits_data_hi_lo_95};
  wire [1:0]       memRequest_bits_data_lo_lo_96 = {_memRequest_bits_data_T_1219[88], _memRequest_bits_data_T_1026[88]};
  wire [1:0]       memRequest_bits_data_lo_hi_96 = {_memRequest_bits_data_T_1605[88], _memRequest_bits_data_T_1412[88]};
  wire [3:0]       memRequest_bits_data_lo_96 = {memRequest_bits_data_lo_hi_96, memRequest_bits_data_lo_lo_96};
  wire [1:0]       memRequest_bits_data_hi_lo_96 = {_memRequest_bits_data_T_1991[88], _memRequest_bits_data_T_1798[88]};
  wire [1:0]       memRequest_bits_data_hi_hi_96 = {_memRequest_bits_data_T_2377[88], _memRequest_bits_data_T_2184[88]};
  wire [3:0]       memRequest_bits_data_hi_96 = {memRequest_bits_data_hi_hi_96, memRequest_bits_data_hi_lo_96};
  wire [1:0]       memRequest_bits_data_lo_lo_97 = {_memRequest_bits_data_T_1219[89], _memRequest_bits_data_T_1026[89]};
  wire [1:0]       memRequest_bits_data_lo_hi_97 = {_memRequest_bits_data_T_1605[89], _memRequest_bits_data_T_1412[89]};
  wire [3:0]       memRequest_bits_data_lo_97 = {memRequest_bits_data_lo_hi_97, memRequest_bits_data_lo_lo_97};
  wire [1:0]       memRequest_bits_data_hi_lo_97 = {_memRequest_bits_data_T_1991[89], _memRequest_bits_data_T_1798[89]};
  wire [1:0]       memRequest_bits_data_hi_hi_97 = {_memRequest_bits_data_T_2377[89], _memRequest_bits_data_T_2184[89]};
  wire [3:0]       memRequest_bits_data_hi_97 = {memRequest_bits_data_hi_hi_97, memRequest_bits_data_hi_lo_97};
  wire [1:0]       memRequest_bits_data_lo_lo_98 = {_memRequest_bits_data_T_1219[90], _memRequest_bits_data_T_1026[90]};
  wire [1:0]       memRequest_bits_data_lo_hi_98 = {_memRequest_bits_data_T_1605[90], _memRequest_bits_data_T_1412[90]};
  wire [3:0]       memRequest_bits_data_lo_98 = {memRequest_bits_data_lo_hi_98, memRequest_bits_data_lo_lo_98};
  wire [1:0]       memRequest_bits_data_hi_lo_98 = {_memRequest_bits_data_T_1991[90], _memRequest_bits_data_T_1798[90]};
  wire [1:0]       memRequest_bits_data_hi_hi_98 = {_memRequest_bits_data_T_2377[90], _memRequest_bits_data_T_2184[90]};
  wire [3:0]       memRequest_bits_data_hi_98 = {memRequest_bits_data_hi_hi_98, memRequest_bits_data_hi_lo_98};
  wire [1:0]       memRequest_bits_data_lo_lo_99 = {_memRequest_bits_data_T_1219[91], _memRequest_bits_data_T_1026[91]};
  wire [1:0]       memRequest_bits_data_lo_hi_99 = {_memRequest_bits_data_T_1605[91], _memRequest_bits_data_T_1412[91]};
  wire [3:0]       memRequest_bits_data_lo_99 = {memRequest_bits_data_lo_hi_99, memRequest_bits_data_lo_lo_99};
  wire [1:0]       memRequest_bits_data_hi_lo_99 = {_memRequest_bits_data_T_1991[91], _memRequest_bits_data_T_1798[91]};
  wire [1:0]       memRequest_bits_data_hi_hi_99 = {_memRequest_bits_data_T_2377[91], _memRequest_bits_data_T_2184[91]};
  wire [3:0]       memRequest_bits_data_hi_99 = {memRequest_bits_data_hi_hi_99, memRequest_bits_data_hi_lo_99};
  wire [1:0]       memRequest_bits_data_lo_lo_100 = {_memRequest_bits_data_T_1219[92], _memRequest_bits_data_T_1026[92]};
  wire [1:0]       memRequest_bits_data_lo_hi_100 = {_memRequest_bits_data_T_1605[92], _memRequest_bits_data_T_1412[92]};
  wire [3:0]       memRequest_bits_data_lo_100 = {memRequest_bits_data_lo_hi_100, memRequest_bits_data_lo_lo_100};
  wire [1:0]       memRequest_bits_data_hi_lo_100 = {_memRequest_bits_data_T_1991[92], _memRequest_bits_data_T_1798[92]};
  wire [1:0]       memRequest_bits_data_hi_hi_100 = {_memRequest_bits_data_T_2377[92], _memRequest_bits_data_T_2184[92]};
  wire [3:0]       memRequest_bits_data_hi_100 = {memRequest_bits_data_hi_hi_100, memRequest_bits_data_hi_lo_100};
  wire [1:0]       memRequest_bits_data_lo_lo_101 = {_memRequest_bits_data_T_1219[93], _memRequest_bits_data_T_1026[93]};
  wire [1:0]       memRequest_bits_data_lo_hi_101 = {_memRequest_bits_data_T_1605[93], _memRequest_bits_data_T_1412[93]};
  wire [3:0]       memRequest_bits_data_lo_101 = {memRequest_bits_data_lo_hi_101, memRequest_bits_data_lo_lo_101};
  wire [1:0]       memRequest_bits_data_hi_lo_101 = {_memRequest_bits_data_T_1991[93], _memRequest_bits_data_T_1798[93]};
  wire [1:0]       memRequest_bits_data_hi_hi_101 = {_memRequest_bits_data_T_2377[93], _memRequest_bits_data_T_2184[93]};
  wire [3:0]       memRequest_bits_data_hi_101 = {memRequest_bits_data_hi_hi_101, memRequest_bits_data_hi_lo_101};
  wire [1:0]       memRequest_bits_data_lo_lo_102 = {_memRequest_bits_data_T_1219[94], _memRequest_bits_data_T_1026[94]};
  wire [1:0]       memRequest_bits_data_lo_hi_102 = {_memRequest_bits_data_T_1605[94], _memRequest_bits_data_T_1412[94]};
  wire [3:0]       memRequest_bits_data_lo_102 = {memRequest_bits_data_lo_hi_102, memRequest_bits_data_lo_lo_102};
  wire [1:0]       memRequest_bits_data_hi_lo_102 = {_memRequest_bits_data_T_1991[94], _memRequest_bits_data_T_1798[94]};
  wire [1:0]       memRequest_bits_data_hi_hi_102 = {_memRequest_bits_data_T_2377[94], _memRequest_bits_data_T_2184[94]};
  wire [3:0]       memRequest_bits_data_hi_102 = {memRequest_bits_data_hi_hi_102, memRequest_bits_data_hi_lo_102};
  wire [1:0]       memRequest_bits_data_lo_lo_103 = {_memRequest_bits_data_T_1219[95], _memRequest_bits_data_T_1026[95]};
  wire [1:0]       memRequest_bits_data_lo_hi_103 = {_memRequest_bits_data_T_1605[95], _memRequest_bits_data_T_1412[95]};
  wire [3:0]       memRequest_bits_data_lo_103 = {memRequest_bits_data_lo_hi_103, memRequest_bits_data_lo_lo_103};
  wire [1:0]       memRequest_bits_data_hi_lo_103 = {_memRequest_bits_data_T_1991[95], _memRequest_bits_data_T_1798[95]};
  wire [1:0]       memRequest_bits_data_hi_hi_103 = {_memRequest_bits_data_T_2377[95], _memRequest_bits_data_T_2184[95]};
  wire [3:0]       memRequest_bits_data_hi_103 = {memRequest_bits_data_hi_hi_103, memRequest_bits_data_hi_lo_103};
  wire [1:0]       memRequest_bits_data_lo_lo_104 = {_memRequest_bits_data_T_1219[96], _memRequest_bits_data_T_1026[96]};
  wire [1:0]       memRequest_bits_data_lo_hi_104 = {_memRequest_bits_data_T_1605[96], _memRequest_bits_data_T_1412[96]};
  wire [3:0]       memRequest_bits_data_lo_104 = {memRequest_bits_data_lo_hi_104, memRequest_bits_data_lo_lo_104};
  wire [1:0]       memRequest_bits_data_hi_lo_104 = {_memRequest_bits_data_T_1991[96], _memRequest_bits_data_T_1798[96]};
  wire [1:0]       memRequest_bits_data_hi_hi_104 = {_memRequest_bits_data_T_2377[96], _memRequest_bits_data_T_2184[96]};
  wire [3:0]       memRequest_bits_data_hi_104 = {memRequest_bits_data_hi_hi_104, memRequest_bits_data_hi_lo_104};
  wire [1:0]       memRequest_bits_data_lo_lo_105 = {_memRequest_bits_data_T_1219[97], _memRequest_bits_data_T_1026[97]};
  wire [1:0]       memRequest_bits_data_lo_hi_105 = {_memRequest_bits_data_T_1605[97], _memRequest_bits_data_T_1412[97]};
  wire [3:0]       memRequest_bits_data_lo_105 = {memRequest_bits_data_lo_hi_105, memRequest_bits_data_lo_lo_105};
  wire [1:0]       memRequest_bits_data_hi_lo_105 = {_memRequest_bits_data_T_1991[97], _memRequest_bits_data_T_1798[97]};
  wire [1:0]       memRequest_bits_data_hi_hi_105 = {_memRequest_bits_data_T_2377[97], _memRequest_bits_data_T_2184[97]};
  wire [3:0]       memRequest_bits_data_hi_105 = {memRequest_bits_data_hi_hi_105, memRequest_bits_data_hi_lo_105};
  wire [1:0]       memRequest_bits_data_lo_lo_106 = {_memRequest_bits_data_T_1219[98], _memRequest_bits_data_T_1026[98]};
  wire [1:0]       memRequest_bits_data_lo_hi_106 = {_memRequest_bits_data_T_1605[98], _memRequest_bits_data_T_1412[98]};
  wire [3:0]       memRequest_bits_data_lo_106 = {memRequest_bits_data_lo_hi_106, memRequest_bits_data_lo_lo_106};
  wire [1:0]       memRequest_bits_data_hi_lo_106 = {_memRequest_bits_data_T_1991[98], _memRequest_bits_data_T_1798[98]};
  wire [1:0]       memRequest_bits_data_hi_hi_106 = {_memRequest_bits_data_T_2377[98], _memRequest_bits_data_T_2184[98]};
  wire [3:0]       memRequest_bits_data_hi_106 = {memRequest_bits_data_hi_hi_106, memRequest_bits_data_hi_lo_106};
  wire [1:0]       memRequest_bits_data_lo_lo_107 = {_memRequest_bits_data_T_1219[99], _memRequest_bits_data_T_1026[99]};
  wire [1:0]       memRequest_bits_data_lo_hi_107 = {_memRequest_bits_data_T_1605[99], _memRequest_bits_data_T_1412[99]};
  wire [3:0]       memRequest_bits_data_lo_107 = {memRequest_bits_data_lo_hi_107, memRequest_bits_data_lo_lo_107};
  wire [1:0]       memRequest_bits_data_hi_lo_107 = {_memRequest_bits_data_T_1991[99], _memRequest_bits_data_T_1798[99]};
  wire [1:0]       memRequest_bits_data_hi_hi_107 = {_memRequest_bits_data_T_2377[99], _memRequest_bits_data_T_2184[99]};
  wire [3:0]       memRequest_bits_data_hi_107 = {memRequest_bits_data_hi_hi_107, memRequest_bits_data_hi_lo_107};
  wire [1:0]       memRequest_bits_data_lo_lo_108 = {_memRequest_bits_data_T_1219[100], _memRequest_bits_data_T_1026[100]};
  wire [1:0]       memRequest_bits_data_lo_hi_108 = {_memRequest_bits_data_T_1605[100], _memRequest_bits_data_T_1412[100]};
  wire [3:0]       memRequest_bits_data_lo_108 = {memRequest_bits_data_lo_hi_108, memRequest_bits_data_lo_lo_108};
  wire [1:0]       memRequest_bits_data_hi_lo_108 = {_memRequest_bits_data_T_1991[100], _memRequest_bits_data_T_1798[100]};
  wire [1:0]       memRequest_bits_data_hi_hi_108 = {_memRequest_bits_data_T_2377[100], _memRequest_bits_data_T_2184[100]};
  wire [3:0]       memRequest_bits_data_hi_108 = {memRequest_bits_data_hi_hi_108, memRequest_bits_data_hi_lo_108};
  wire [1:0]       memRequest_bits_data_lo_lo_109 = {_memRequest_bits_data_T_1219[101], _memRequest_bits_data_T_1026[101]};
  wire [1:0]       memRequest_bits_data_lo_hi_109 = {_memRequest_bits_data_T_1605[101], _memRequest_bits_data_T_1412[101]};
  wire [3:0]       memRequest_bits_data_lo_109 = {memRequest_bits_data_lo_hi_109, memRequest_bits_data_lo_lo_109};
  wire [1:0]       memRequest_bits_data_hi_lo_109 = {_memRequest_bits_data_T_1991[101], _memRequest_bits_data_T_1798[101]};
  wire [1:0]       memRequest_bits_data_hi_hi_109 = {_memRequest_bits_data_T_2377[101], _memRequest_bits_data_T_2184[101]};
  wire [3:0]       memRequest_bits_data_hi_109 = {memRequest_bits_data_hi_hi_109, memRequest_bits_data_hi_lo_109};
  wire [1:0]       memRequest_bits_data_lo_lo_110 = {_memRequest_bits_data_T_1219[102], _memRequest_bits_data_T_1026[102]};
  wire [1:0]       memRequest_bits_data_lo_hi_110 = {_memRequest_bits_data_T_1605[102], _memRequest_bits_data_T_1412[102]};
  wire [3:0]       memRequest_bits_data_lo_110 = {memRequest_bits_data_lo_hi_110, memRequest_bits_data_lo_lo_110};
  wire [1:0]       memRequest_bits_data_hi_lo_110 = {_memRequest_bits_data_T_1991[102], _memRequest_bits_data_T_1798[102]};
  wire [1:0]       memRequest_bits_data_hi_hi_110 = {_memRequest_bits_data_T_2377[102], _memRequest_bits_data_T_2184[102]};
  wire [3:0]       memRequest_bits_data_hi_110 = {memRequest_bits_data_hi_hi_110, memRequest_bits_data_hi_lo_110};
  wire [1:0]       memRequest_bits_data_lo_lo_111 = {_memRequest_bits_data_T_1219[103], _memRequest_bits_data_T_1026[103]};
  wire [1:0]       memRequest_bits_data_lo_hi_111 = {_memRequest_bits_data_T_1605[103], _memRequest_bits_data_T_1412[103]};
  wire [3:0]       memRequest_bits_data_lo_111 = {memRequest_bits_data_lo_hi_111, memRequest_bits_data_lo_lo_111};
  wire [1:0]       memRequest_bits_data_hi_lo_111 = {_memRequest_bits_data_T_1991[103], _memRequest_bits_data_T_1798[103]};
  wire [1:0]       memRequest_bits_data_hi_hi_111 = {_memRequest_bits_data_T_2377[103], _memRequest_bits_data_T_2184[103]};
  wire [3:0]       memRequest_bits_data_hi_111 = {memRequest_bits_data_hi_hi_111, memRequest_bits_data_hi_lo_111};
  wire [1:0]       memRequest_bits_data_lo_lo_112 = {_memRequest_bits_data_T_1219[104], _memRequest_bits_data_T_1026[104]};
  wire [1:0]       memRequest_bits_data_lo_hi_112 = {_memRequest_bits_data_T_1605[104], _memRequest_bits_data_T_1412[104]};
  wire [3:0]       memRequest_bits_data_lo_112 = {memRequest_bits_data_lo_hi_112, memRequest_bits_data_lo_lo_112};
  wire [1:0]       memRequest_bits_data_hi_lo_112 = {_memRequest_bits_data_T_1991[104], _memRequest_bits_data_T_1798[104]};
  wire [1:0]       memRequest_bits_data_hi_hi_112 = {_memRequest_bits_data_T_2377[104], _memRequest_bits_data_T_2184[104]};
  wire [3:0]       memRequest_bits_data_hi_112 = {memRequest_bits_data_hi_hi_112, memRequest_bits_data_hi_lo_112};
  wire [1:0]       memRequest_bits_data_lo_lo_113 = {_memRequest_bits_data_T_1219[105], _memRequest_bits_data_T_1026[105]};
  wire [1:0]       memRequest_bits_data_lo_hi_113 = {_memRequest_bits_data_T_1605[105], _memRequest_bits_data_T_1412[105]};
  wire [3:0]       memRequest_bits_data_lo_113 = {memRequest_bits_data_lo_hi_113, memRequest_bits_data_lo_lo_113};
  wire [1:0]       memRequest_bits_data_hi_lo_113 = {_memRequest_bits_data_T_1991[105], _memRequest_bits_data_T_1798[105]};
  wire [1:0]       memRequest_bits_data_hi_hi_113 = {_memRequest_bits_data_T_2377[105], _memRequest_bits_data_T_2184[105]};
  wire [3:0]       memRequest_bits_data_hi_113 = {memRequest_bits_data_hi_hi_113, memRequest_bits_data_hi_lo_113};
  wire [1:0]       memRequest_bits_data_lo_lo_114 = {_memRequest_bits_data_T_1219[106], _memRequest_bits_data_T_1026[106]};
  wire [1:0]       memRequest_bits_data_lo_hi_114 = {_memRequest_bits_data_T_1605[106], _memRequest_bits_data_T_1412[106]};
  wire [3:0]       memRequest_bits_data_lo_114 = {memRequest_bits_data_lo_hi_114, memRequest_bits_data_lo_lo_114};
  wire [1:0]       memRequest_bits_data_hi_lo_114 = {_memRequest_bits_data_T_1991[106], _memRequest_bits_data_T_1798[106]};
  wire [1:0]       memRequest_bits_data_hi_hi_114 = {_memRequest_bits_data_T_2377[106], _memRequest_bits_data_T_2184[106]};
  wire [3:0]       memRequest_bits_data_hi_114 = {memRequest_bits_data_hi_hi_114, memRequest_bits_data_hi_lo_114};
  wire [1:0]       memRequest_bits_data_lo_lo_115 = {_memRequest_bits_data_T_1219[107], _memRequest_bits_data_T_1026[107]};
  wire [1:0]       memRequest_bits_data_lo_hi_115 = {_memRequest_bits_data_T_1605[107], _memRequest_bits_data_T_1412[107]};
  wire [3:0]       memRequest_bits_data_lo_115 = {memRequest_bits_data_lo_hi_115, memRequest_bits_data_lo_lo_115};
  wire [1:0]       memRequest_bits_data_hi_lo_115 = {_memRequest_bits_data_T_1991[107], _memRequest_bits_data_T_1798[107]};
  wire [1:0]       memRequest_bits_data_hi_hi_115 = {_memRequest_bits_data_T_2377[107], _memRequest_bits_data_T_2184[107]};
  wire [3:0]       memRequest_bits_data_hi_115 = {memRequest_bits_data_hi_hi_115, memRequest_bits_data_hi_lo_115};
  wire [1:0]       memRequest_bits_data_lo_lo_116 = {_memRequest_bits_data_T_1219[108], _memRequest_bits_data_T_1026[108]};
  wire [1:0]       memRequest_bits_data_lo_hi_116 = {_memRequest_bits_data_T_1605[108], _memRequest_bits_data_T_1412[108]};
  wire [3:0]       memRequest_bits_data_lo_116 = {memRequest_bits_data_lo_hi_116, memRequest_bits_data_lo_lo_116};
  wire [1:0]       memRequest_bits_data_hi_lo_116 = {_memRequest_bits_data_T_1991[108], _memRequest_bits_data_T_1798[108]};
  wire [1:0]       memRequest_bits_data_hi_hi_116 = {_memRequest_bits_data_T_2377[108], _memRequest_bits_data_T_2184[108]};
  wire [3:0]       memRequest_bits_data_hi_116 = {memRequest_bits_data_hi_hi_116, memRequest_bits_data_hi_lo_116};
  wire [1:0]       memRequest_bits_data_lo_lo_117 = {_memRequest_bits_data_T_1219[109], _memRequest_bits_data_T_1026[109]};
  wire [1:0]       memRequest_bits_data_lo_hi_117 = {_memRequest_bits_data_T_1605[109], _memRequest_bits_data_T_1412[109]};
  wire [3:0]       memRequest_bits_data_lo_117 = {memRequest_bits_data_lo_hi_117, memRequest_bits_data_lo_lo_117};
  wire [1:0]       memRequest_bits_data_hi_lo_117 = {_memRequest_bits_data_T_1991[109], _memRequest_bits_data_T_1798[109]};
  wire [1:0]       memRequest_bits_data_hi_hi_117 = {_memRequest_bits_data_T_2377[109], _memRequest_bits_data_T_2184[109]};
  wire [3:0]       memRequest_bits_data_hi_117 = {memRequest_bits_data_hi_hi_117, memRequest_bits_data_hi_lo_117};
  wire [1:0]       memRequest_bits_data_lo_lo_118 = {_memRequest_bits_data_T_1219[110], _memRequest_bits_data_T_1026[110]};
  wire [1:0]       memRequest_bits_data_lo_hi_118 = {_memRequest_bits_data_T_1605[110], _memRequest_bits_data_T_1412[110]};
  wire [3:0]       memRequest_bits_data_lo_118 = {memRequest_bits_data_lo_hi_118, memRequest_bits_data_lo_lo_118};
  wire [1:0]       memRequest_bits_data_hi_lo_118 = {_memRequest_bits_data_T_1991[110], _memRequest_bits_data_T_1798[110]};
  wire [1:0]       memRequest_bits_data_hi_hi_118 = {_memRequest_bits_data_T_2377[110], _memRequest_bits_data_T_2184[110]};
  wire [3:0]       memRequest_bits_data_hi_118 = {memRequest_bits_data_hi_hi_118, memRequest_bits_data_hi_lo_118};
  wire [1:0]       memRequest_bits_data_lo_lo_119 = {_memRequest_bits_data_T_1219[111], _memRequest_bits_data_T_1026[111]};
  wire [1:0]       memRequest_bits_data_lo_hi_119 = {_memRequest_bits_data_T_1605[111], _memRequest_bits_data_T_1412[111]};
  wire [3:0]       memRequest_bits_data_lo_119 = {memRequest_bits_data_lo_hi_119, memRequest_bits_data_lo_lo_119};
  wire [1:0]       memRequest_bits_data_hi_lo_119 = {_memRequest_bits_data_T_1991[111], _memRequest_bits_data_T_1798[111]};
  wire [1:0]       memRequest_bits_data_hi_hi_119 = {_memRequest_bits_data_T_2377[111], _memRequest_bits_data_T_2184[111]};
  wire [3:0]       memRequest_bits_data_hi_119 = {memRequest_bits_data_hi_hi_119, memRequest_bits_data_hi_lo_119};
  wire [1:0]       memRequest_bits_data_lo_lo_120 = {_memRequest_bits_data_T_1219[112], _memRequest_bits_data_T_1026[112]};
  wire [1:0]       memRequest_bits_data_lo_hi_120 = {_memRequest_bits_data_T_1605[112], _memRequest_bits_data_T_1412[112]};
  wire [3:0]       memRequest_bits_data_lo_120 = {memRequest_bits_data_lo_hi_120, memRequest_bits_data_lo_lo_120};
  wire [1:0]       memRequest_bits_data_hi_lo_120 = {_memRequest_bits_data_T_1991[112], _memRequest_bits_data_T_1798[112]};
  wire [1:0]       memRequest_bits_data_hi_hi_120 = {_memRequest_bits_data_T_2377[112], _memRequest_bits_data_T_2184[112]};
  wire [3:0]       memRequest_bits_data_hi_120 = {memRequest_bits_data_hi_hi_120, memRequest_bits_data_hi_lo_120};
  wire [1:0]       memRequest_bits_data_lo_lo_121 = {_memRequest_bits_data_T_1219[113], _memRequest_bits_data_T_1026[113]};
  wire [1:0]       memRequest_bits_data_lo_hi_121 = {_memRequest_bits_data_T_1605[113], _memRequest_bits_data_T_1412[113]};
  wire [3:0]       memRequest_bits_data_lo_121 = {memRequest_bits_data_lo_hi_121, memRequest_bits_data_lo_lo_121};
  wire [1:0]       memRequest_bits_data_hi_lo_121 = {_memRequest_bits_data_T_1991[113], _memRequest_bits_data_T_1798[113]};
  wire [1:0]       memRequest_bits_data_hi_hi_121 = {_memRequest_bits_data_T_2377[113], _memRequest_bits_data_T_2184[113]};
  wire [3:0]       memRequest_bits_data_hi_121 = {memRequest_bits_data_hi_hi_121, memRequest_bits_data_hi_lo_121};
  wire [1:0]       memRequest_bits_data_lo_lo_122 = {_memRequest_bits_data_T_1219[114], _memRequest_bits_data_T_1026[114]};
  wire [1:0]       memRequest_bits_data_lo_hi_122 = {_memRequest_bits_data_T_1605[114], _memRequest_bits_data_T_1412[114]};
  wire [3:0]       memRequest_bits_data_lo_122 = {memRequest_bits_data_lo_hi_122, memRequest_bits_data_lo_lo_122};
  wire [1:0]       memRequest_bits_data_hi_lo_122 = {_memRequest_bits_data_T_1991[114], _memRequest_bits_data_T_1798[114]};
  wire [1:0]       memRequest_bits_data_hi_hi_122 = {_memRequest_bits_data_T_2377[114], _memRequest_bits_data_T_2184[114]};
  wire [3:0]       memRequest_bits_data_hi_122 = {memRequest_bits_data_hi_hi_122, memRequest_bits_data_hi_lo_122};
  wire [1:0]       memRequest_bits_data_lo_lo_123 = {_memRequest_bits_data_T_1219[115], _memRequest_bits_data_T_1026[115]};
  wire [1:0]       memRequest_bits_data_lo_hi_123 = {_memRequest_bits_data_T_1605[115], _memRequest_bits_data_T_1412[115]};
  wire [3:0]       memRequest_bits_data_lo_123 = {memRequest_bits_data_lo_hi_123, memRequest_bits_data_lo_lo_123};
  wire [1:0]       memRequest_bits_data_hi_lo_123 = {_memRequest_bits_data_T_1991[115], _memRequest_bits_data_T_1798[115]};
  wire [1:0]       memRequest_bits_data_hi_hi_123 = {_memRequest_bits_data_T_2377[115], _memRequest_bits_data_T_2184[115]};
  wire [3:0]       memRequest_bits_data_hi_123 = {memRequest_bits_data_hi_hi_123, memRequest_bits_data_hi_lo_123};
  wire [1:0]       memRequest_bits_data_lo_lo_124 = {_memRequest_bits_data_T_1219[116], _memRequest_bits_data_T_1026[116]};
  wire [1:0]       memRequest_bits_data_lo_hi_124 = {_memRequest_bits_data_T_1605[116], _memRequest_bits_data_T_1412[116]};
  wire [3:0]       memRequest_bits_data_lo_124 = {memRequest_bits_data_lo_hi_124, memRequest_bits_data_lo_lo_124};
  wire [1:0]       memRequest_bits_data_hi_lo_124 = {_memRequest_bits_data_T_1991[116], _memRequest_bits_data_T_1798[116]};
  wire [1:0]       memRequest_bits_data_hi_hi_124 = {_memRequest_bits_data_T_2377[116], _memRequest_bits_data_T_2184[116]};
  wire [3:0]       memRequest_bits_data_hi_124 = {memRequest_bits_data_hi_hi_124, memRequest_bits_data_hi_lo_124};
  wire [1:0]       memRequest_bits_data_lo_lo_125 = {_memRequest_bits_data_T_1219[117], _memRequest_bits_data_T_1026[117]};
  wire [1:0]       memRequest_bits_data_lo_hi_125 = {_memRequest_bits_data_T_1605[117], _memRequest_bits_data_T_1412[117]};
  wire [3:0]       memRequest_bits_data_lo_125 = {memRequest_bits_data_lo_hi_125, memRequest_bits_data_lo_lo_125};
  wire [1:0]       memRequest_bits_data_hi_lo_125 = {_memRequest_bits_data_T_1991[117], _memRequest_bits_data_T_1798[117]};
  wire [1:0]       memRequest_bits_data_hi_hi_125 = {_memRequest_bits_data_T_2377[117], _memRequest_bits_data_T_2184[117]};
  wire [3:0]       memRequest_bits_data_hi_125 = {memRequest_bits_data_hi_hi_125, memRequest_bits_data_hi_lo_125};
  wire [1:0]       memRequest_bits_data_lo_lo_126 = {_memRequest_bits_data_T_1219[118], _memRequest_bits_data_T_1026[118]};
  wire [1:0]       memRequest_bits_data_lo_hi_126 = {_memRequest_bits_data_T_1605[118], _memRequest_bits_data_T_1412[118]};
  wire [3:0]       memRequest_bits_data_lo_126 = {memRequest_bits_data_lo_hi_126, memRequest_bits_data_lo_lo_126};
  wire [1:0]       memRequest_bits_data_hi_lo_126 = {_memRequest_bits_data_T_1991[118], _memRequest_bits_data_T_1798[118]};
  wire [1:0]       memRequest_bits_data_hi_hi_126 = {_memRequest_bits_data_T_2377[118], _memRequest_bits_data_T_2184[118]};
  wire [3:0]       memRequest_bits_data_hi_126 = {memRequest_bits_data_hi_hi_126, memRequest_bits_data_hi_lo_126};
  wire [1:0]       memRequest_bits_data_lo_lo_127 = {_memRequest_bits_data_T_1219[119], _memRequest_bits_data_T_1026[119]};
  wire [1:0]       memRequest_bits_data_lo_hi_127 = {_memRequest_bits_data_T_1605[119], _memRequest_bits_data_T_1412[119]};
  wire [3:0]       memRequest_bits_data_lo_127 = {memRequest_bits_data_lo_hi_127, memRequest_bits_data_lo_lo_127};
  wire [1:0]       memRequest_bits_data_hi_lo_127 = {_memRequest_bits_data_T_1991[119], _memRequest_bits_data_T_1798[119]};
  wire [1:0]       memRequest_bits_data_hi_hi_127 = {_memRequest_bits_data_T_2377[119], _memRequest_bits_data_T_2184[119]};
  wire [3:0]       memRequest_bits_data_hi_127 = {memRequest_bits_data_hi_hi_127, memRequest_bits_data_hi_lo_127};
  wire [1:0]       memRequest_bits_data_lo_lo_128 = {_memRequest_bits_data_T_1219[120], _memRequest_bits_data_T_1026[120]};
  wire [1:0]       memRequest_bits_data_lo_hi_128 = {_memRequest_bits_data_T_1605[120], _memRequest_bits_data_T_1412[120]};
  wire [3:0]       memRequest_bits_data_lo_128 = {memRequest_bits_data_lo_hi_128, memRequest_bits_data_lo_lo_128};
  wire [1:0]       memRequest_bits_data_hi_lo_128 = {_memRequest_bits_data_T_1991[120], _memRequest_bits_data_T_1798[120]};
  wire [1:0]       memRequest_bits_data_hi_hi_128 = {_memRequest_bits_data_T_2377[120], _memRequest_bits_data_T_2184[120]};
  wire [3:0]       memRequest_bits_data_hi_128 = {memRequest_bits_data_hi_hi_128, memRequest_bits_data_hi_lo_128};
  wire [1:0]       memRequest_bits_data_lo_lo_129 = {_memRequest_bits_data_T_1219[121], _memRequest_bits_data_T_1026[121]};
  wire [1:0]       memRequest_bits_data_lo_hi_129 = {_memRequest_bits_data_T_1605[121], _memRequest_bits_data_T_1412[121]};
  wire [3:0]       memRequest_bits_data_lo_129 = {memRequest_bits_data_lo_hi_129, memRequest_bits_data_lo_lo_129};
  wire [1:0]       memRequest_bits_data_hi_lo_129 = {_memRequest_bits_data_T_1991[121], _memRequest_bits_data_T_1798[121]};
  wire [1:0]       memRequest_bits_data_hi_hi_129 = {_memRequest_bits_data_T_2377[121], _memRequest_bits_data_T_2184[121]};
  wire [3:0]       memRequest_bits_data_hi_129 = {memRequest_bits_data_hi_hi_129, memRequest_bits_data_hi_lo_129};
  wire [1:0]       memRequest_bits_data_lo_lo_130 = {_memRequest_bits_data_T_1219[122], _memRequest_bits_data_T_1026[122]};
  wire [1:0]       memRequest_bits_data_lo_hi_130 = {_memRequest_bits_data_T_1605[122], _memRequest_bits_data_T_1412[122]};
  wire [3:0]       memRequest_bits_data_lo_130 = {memRequest_bits_data_lo_hi_130, memRequest_bits_data_lo_lo_130};
  wire [1:0]       memRequest_bits_data_hi_lo_130 = {_memRequest_bits_data_T_1991[122], _memRequest_bits_data_T_1798[122]};
  wire [1:0]       memRequest_bits_data_hi_hi_130 = {_memRequest_bits_data_T_2377[122], _memRequest_bits_data_T_2184[122]};
  wire [3:0]       memRequest_bits_data_hi_130 = {memRequest_bits_data_hi_hi_130, memRequest_bits_data_hi_lo_130};
  wire [1:0]       memRequest_bits_data_lo_lo_131 = {_memRequest_bits_data_T_1219[123], _memRequest_bits_data_T_1026[123]};
  wire [1:0]       memRequest_bits_data_lo_hi_131 = {_memRequest_bits_data_T_1605[123], _memRequest_bits_data_T_1412[123]};
  wire [3:0]       memRequest_bits_data_lo_131 = {memRequest_bits_data_lo_hi_131, memRequest_bits_data_lo_lo_131};
  wire [1:0]       memRequest_bits_data_hi_lo_131 = {_memRequest_bits_data_T_1991[123], _memRequest_bits_data_T_1798[123]};
  wire [1:0]       memRequest_bits_data_hi_hi_131 = {_memRequest_bits_data_T_2377[123], _memRequest_bits_data_T_2184[123]};
  wire [3:0]       memRequest_bits_data_hi_131 = {memRequest_bits_data_hi_hi_131, memRequest_bits_data_hi_lo_131};
  wire [1:0]       memRequest_bits_data_lo_lo_132 = {_memRequest_bits_data_T_1219[124], _memRequest_bits_data_T_1026[124]};
  wire [1:0]       memRequest_bits_data_lo_hi_132 = {_memRequest_bits_data_T_1605[124], _memRequest_bits_data_T_1412[124]};
  wire [3:0]       memRequest_bits_data_lo_132 = {memRequest_bits_data_lo_hi_132, memRequest_bits_data_lo_lo_132};
  wire [1:0]       memRequest_bits_data_hi_lo_132 = {_memRequest_bits_data_T_1991[124], _memRequest_bits_data_T_1798[124]};
  wire [1:0]       memRequest_bits_data_hi_hi_132 = {_memRequest_bits_data_T_2377[124], _memRequest_bits_data_T_2184[124]};
  wire [3:0]       memRequest_bits_data_hi_132 = {memRequest_bits_data_hi_hi_132, memRequest_bits_data_hi_lo_132};
  wire [1:0]       memRequest_bits_data_lo_lo_133 = {_memRequest_bits_data_T_1219[125], _memRequest_bits_data_T_1026[125]};
  wire [1:0]       memRequest_bits_data_lo_hi_133 = {_memRequest_bits_data_T_1605[125], _memRequest_bits_data_T_1412[125]};
  wire [3:0]       memRequest_bits_data_lo_133 = {memRequest_bits_data_lo_hi_133, memRequest_bits_data_lo_lo_133};
  wire [1:0]       memRequest_bits_data_hi_lo_133 = {_memRequest_bits_data_T_1991[125], _memRequest_bits_data_T_1798[125]};
  wire [1:0]       memRequest_bits_data_hi_hi_133 = {_memRequest_bits_data_T_2377[125], _memRequest_bits_data_T_2184[125]};
  wire [3:0]       memRequest_bits_data_hi_133 = {memRequest_bits_data_hi_hi_133, memRequest_bits_data_hi_lo_133};
  wire [1:0]       memRequest_bits_data_lo_lo_134 = {_memRequest_bits_data_T_1219[126], _memRequest_bits_data_T_1026[126]};
  wire [1:0]       memRequest_bits_data_lo_hi_134 = {_memRequest_bits_data_T_1605[126], _memRequest_bits_data_T_1412[126]};
  wire [3:0]       memRequest_bits_data_lo_134 = {memRequest_bits_data_lo_hi_134, memRequest_bits_data_lo_lo_134};
  wire [1:0]       memRequest_bits_data_hi_lo_134 = {_memRequest_bits_data_T_1991[126], _memRequest_bits_data_T_1798[126]};
  wire [1:0]       memRequest_bits_data_hi_hi_134 = {_memRequest_bits_data_T_2377[126], _memRequest_bits_data_T_2184[126]};
  wire [3:0]       memRequest_bits_data_hi_134 = {memRequest_bits_data_hi_hi_134, memRequest_bits_data_hi_lo_134};
  wire [1:0]       memRequest_bits_data_lo_lo_135 = {_memRequest_bits_data_T_1219[127], _memRequest_bits_data_T_1026[127]};
  wire [1:0]       memRequest_bits_data_lo_hi_135 = {_memRequest_bits_data_T_1605[127], _memRequest_bits_data_T_1412[127]};
  wire [3:0]       memRequest_bits_data_lo_135 = {memRequest_bits_data_lo_hi_135, memRequest_bits_data_lo_lo_135};
  wire [1:0]       memRequest_bits_data_hi_lo_135 = {_memRequest_bits_data_T_1991[127], _memRequest_bits_data_T_1798[127]};
  wire [1:0]       memRequest_bits_data_hi_hi_135 = {_memRequest_bits_data_T_2377[127], _memRequest_bits_data_T_2184[127]};
  wire [3:0]       memRequest_bits_data_hi_135 = {memRequest_bits_data_hi_hi_135, memRequest_bits_data_hi_lo_135};
  wire [1:0]       memRequest_bits_data_lo_lo_136 = {_memRequest_bits_data_T_1219[128], _memRequest_bits_data_T_1026[128]};
  wire [1:0]       memRequest_bits_data_lo_hi_136 = {_memRequest_bits_data_T_1605[128], _memRequest_bits_data_T_1412[128]};
  wire [3:0]       memRequest_bits_data_lo_136 = {memRequest_bits_data_lo_hi_136, memRequest_bits_data_lo_lo_136};
  wire [1:0]       memRequest_bits_data_hi_lo_136 = {_memRequest_bits_data_T_1991[128], _memRequest_bits_data_T_1798[128]};
  wire [1:0]       memRequest_bits_data_hi_hi_136 = {_memRequest_bits_data_T_2377[128], _memRequest_bits_data_T_2184[128]};
  wire [3:0]       memRequest_bits_data_hi_136 = {memRequest_bits_data_hi_hi_136, memRequest_bits_data_hi_lo_136};
  wire [1:0]       memRequest_bits_data_lo_lo_137 = {_memRequest_bits_data_T_1219[129], _memRequest_bits_data_T_1026[129]};
  wire [1:0]       memRequest_bits_data_lo_hi_137 = {_memRequest_bits_data_T_1605[129], _memRequest_bits_data_T_1412[129]};
  wire [3:0]       memRequest_bits_data_lo_137 = {memRequest_bits_data_lo_hi_137, memRequest_bits_data_lo_lo_137};
  wire [1:0]       memRequest_bits_data_hi_lo_137 = {_memRequest_bits_data_T_1991[129], _memRequest_bits_data_T_1798[129]};
  wire [1:0]       memRequest_bits_data_hi_hi_137 = {_memRequest_bits_data_T_2377[129], _memRequest_bits_data_T_2184[129]};
  wire [3:0]       memRequest_bits_data_hi_137 = {memRequest_bits_data_hi_hi_137, memRequest_bits_data_hi_lo_137};
  wire [1:0]       memRequest_bits_data_lo_lo_138 = {_memRequest_bits_data_T_1219[130], _memRequest_bits_data_T_1026[130]};
  wire [1:0]       memRequest_bits_data_lo_hi_138 = {_memRequest_bits_data_T_1605[130], _memRequest_bits_data_T_1412[130]};
  wire [3:0]       memRequest_bits_data_lo_138 = {memRequest_bits_data_lo_hi_138, memRequest_bits_data_lo_lo_138};
  wire [1:0]       memRequest_bits_data_hi_lo_138 = {_memRequest_bits_data_T_1991[130], _memRequest_bits_data_T_1798[130]};
  wire [1:0]       memRequest_bits_data_hi_hi_138 = {_memRequest_bits_data_T_2377[130], _memRequest_bits_data_T_2184[130]};
  wire [3:0]       memRequest_bits_data_hi_138 = {memRequest_bits_data_hi_hi_138, memRequest_bits_data_hi_lo_138};
  wire [1:0]       memRequest_bits_data_lo_lo_139 = {_memRequest_bits_data_T_1219[131], _memRequest_bits_data_T_1026[131]};
  wire [1:0]       memRequest_bits_data_lo_hi_139 = {_memRequest_bits_data_T_1605[131], _memRequest_bits_data_T_1412[131]};
  wire [3:0]       memRequest_bits_data_lo_139 = {memRequest_bits_data_lo_hi_139, memRequest_bits_data_lo_lo_139};
  wire [1:0]       memRequest_bits_data_hi_lo_139 = {_memRequest_bits_data_T_1991[131], _memRequest_bits_data_T_1798[131]};
  wire [1:0]       memRequest_bits_data_hi_hi_139 = {_memRequest_bits_data_T_2377[131], _memRequest_bits_data_T_2184[131]};
  wire [3:0]       memRequest_bits_data_hi_139 = {memRequest_bits_data_hi_hi_139, memRequest_bits_data_hi_lo_139};
  wire [1:0]       memRequest_bits_data_lo_lo_140 = {_memRequest_bits_data_T_1219[132], _memRequest_bits_data_T_1026[132]};
  wire [1:0]       memRequest_bits_data_lo_hi_140 = {_memRequest_bits_data_T_1605[132], _memRequest_bits_data_T_1412[132]};
  wire [3:0]       memRequest_bits_data_lo_140 = {memRequest_bits_data_lo_hi_140, memRequest_bits_data_lo_lo_140};
  wire [1:0]       memRequest_bits_data_hi_lo_140 = {_memRequest_bits_data_T_1991[132], _memRequest_bits_data_T_1798[132]};
  wire [1:0]       memRequest_bits_data_hi_hi_140 = {_memRequest_bits_data_T_2377[132], _memRequest_bits_data_T_2184[132]};
  wire [3:0]       memRequest_bits_data_hi_140 = {memRequest_bits_data_hi_hi_140, memRequest_bits_data_hi_lo_140};
  wire [1:0]       memRequest_bits_data_lo_lo_141 = {_memRequest_bits_data_T_1219[133], _memRequest_bits_data_T_1026[133]};
  wire [1:0]       memRequest_bits_data_lo_hi_141 = {_memRequest_bits_data_T_1605[133], _memRequest_bits_data_T_1412[133]};
  wire [3:0]       memRequest_bits_data_lo_141 = {memRequest_bits_data_lo_hi_141, memRequest_bits_data_lo_lo_141};
  wire [1:0]       memRequest_bits_data_hi_lo_141 = {_memRequest_bits_data_T_1991[133], _memRequest_bits_data_T_1798[133]};
  wire [1:0]       memRequest_bits_data_hi_hi_141 = {_memRequest_bits_data_T_2377[133], _memRequest_bits_data_T_2184[133]};
  wire [3:0]       memRequest_bits_data_hi_141 = {memRequest_bits_data_hi_hi_141, memRequest_bits_data_hi_lo_141};
  wire [1:0]       memRequest_bits_data_lo_lo_142 = {_memRequest_bits_data_T_1219[134], _memRequest_bits_data_T_1026[134]};
  wire [1:0]       memRequest_bits_data_lo_hi_142 = {_memRequest_bits_data_T_1605[134], _memRequest_bits_data_T_1412[134]};
  wire [3:0]       memRequest_bits_data_lo_142 = {memRequest_bits_data_lo_hi_142, memRequest_bits_data_lo_lo_142};
  wire [1:0]       memRequest_bits_data_hi_lo_142 = {_memRequest_bits_data_T_1991[134], _memRequest_bits_data_T_1798[134]};
  wire [1:0]       memRequest_bits_data_hi_hi_142 = {_memRequest_bits_data_T_2377[134], _memRequest_bits_data_T_2184[134]};
  wire [3:0]       memRequest_bits_data_hi_142 = {memRequest_bits_data_hi_hi_142, memRequest_bits_data_hi_lo_142};
  wire [1:0]       memRequest_bits_data_lo_lo_143 = {_memRequest_bits_data_T_1219[135], _memRequest_bits_data_T_1026[135]};
  wire [1:0]       memRequest_bits_data_lo_hi_143 = {_memRequest_bits_data_T_1605[135], _memRequest_bits_data_T_1412[135]};
  wire [3:0]       memRequest_bits_data_lo_143 = {memRequest_bits_data_lo_hi_143, memRequest_bits_data_lo_lo_143};
  wire [1:0]       memRequest_bits_data_hi_lo_143 = {_memRequest_bits_data_T_1991[135], _memRequest_bits_data_T_1798[135]};
  wire [1:0]       memRequest_bits_data_hi_hi_143 = {_memRequest_bits_data_T_2377[135], _memRequest_bits_data_T_2184[135]};
  wire [3:0]       memRequest_bits_data_hi_143 = {memRequest_bits_data_hi_hi_143, memRequest_bits_data_hi_lo_143};
  wire [1:0]       memRequest_bits_data_lo_lo_144 = {_memRequest_bits_data_T_1219[136], _memRequest_bits_data_T_1026[136]};
  wire [1:0]       memRequest_bits_data_lo_hi_144 = {_memRequest_bits_data_T_1605[136], _memRequest_bits_data_T_1412[136]};
  wire [3:0]       memRequest_bits_data_lo_144 = {memRequest_bits_data_lo_hi_144, memRequest_bits_data_lo_lo_144};
  wire [1:0]       memRequest_bits_data_hi_lo_144 = {_memRequest_bits_data_T_1991[136], _memRequest_bits_data_T_1798[136]};
  wire [1:0]       memRequest_bits_data_hi_hi_144 = {_memRequest_bits_data_T_2377[136], _memRequest_bits_data_T_2184[136]};
  wire [3:0]       memRequest_bits_data_hi_144 = {memRequest_bits_data_hi_hi_144, memRequest_bits_data_hi_lo_144};
  wire [1:0]       memRequest_bits_data_lo_lo_145 = {_memRequest_bits_data_T_1219[137], _memRequest_bits_data_T_1026[137]};
  wire [1:0]       memRequest_bits_data_lo_hi_145 = {_memRequest_bits_data_T_1605[137], _memRequest_bits_data_T_1412[137]};
  wire [3:0]       memRequest_bits_data_lo_145 = {memRequest_bits_data_lo_hi_145, memRequest_bits_data_lo_lo_145};
  wire [1:0]       memRequest_bits_data_hi_lo_145 = {_memRequest_bits_data_T_1991[137], _memRequest_bits_data_T_1798[137]};
  wire [1:0]       memRequest_bits_data_hi_hi_145 = {_memRequest_bits_data_T_2377[137], _memRequest_bits_data_T_2184[137]};
  wire [3:0]       memRequest_bits_data_hi_145 = {memRequest_bits_data_hi_hi_145, memRequest_bits_data_hi_lo_145};
  wire [1:0]       memRequest_bits_data_lo_lo_146 = {_memRequest_bits_data_T_1219[138], _memRequest_bits_data_T_1026[138]};
  wire [1:0]       memRequest_bits_data_lo_hi_146 = {_memRequest_bits_data_T_1605[138], _memRequest_bits_data_T_1412[138]};
  wire [3:0]       memRequest_bits_data_lo_146 = {memRequest_bits_data_lo_hi_146, memRequest_bits_data_lo_lo_146};
  wire [1:0]       memRequest_bits_data_hi_lo_146 = {_memRequest_bits_data_T_1991[138], _memRequest_bits_data_T_1798[138]};
  wire [1:0]       memRequest_bits_data_hi_hi_146 = {_memRequest_bits_data_T_2377[138], _memRequest_bits_data_T_2184[138]};
  wire [3:0]       memRequest_bits_data_hi_146 = {memRequest_bits_data_hi_hi_146, memRequest_bits_data_hi_lo_146};
  wire [1:0]       memRequest_bits_data_lo_lo_147 = {_memRequest_bits_data_T_1219[139], _memRequest_bits_data_T_1026[139]};
  wire [1:0]       memRequest_bits_data_lo_hi_147 = {_memRequest_bits_data_T_1605[139], _memRequest_bits_data_T_1412[139]};
  wire [3:0]       memRequest_bits_data_lo_147 = {memRequest_bits_data_lo_hi_147, memRequest_bits_data_lo_lo_147};
  wire [1:0]       memRequest_bits_data_hi_lo_147 = {_memRequest_bits_data_T_1991[139], _memRequest_bits_data_T_1798[139]};
  wire [1:0]       memRequest_bits_data_hi_hi_147 = {_memRequest_bits_data_T_2377[139], _memRequest_bits_data_T_2184[139]};
  wire [3:0]       memRequest_bits_data_hi_147 = {memRequest_bits_data_hi_hi_147, memRequest_bits_data_hi_lo_147};
  wire [1:0]       memRequest_bits_data_lo_lo_148 = {_memRequest_bits_data_T_1219[140], _memRequest_bits_data_T_1026[140]};
  wire [1:0]       memRequest_bits_data_lo_hi_148 = {_memRequest_bits_data_T_1605[140], _memRequest_bits_data_T_1412[140]};
  wire [3:0]       memRequest_bits_data_lo_148 = {memRequest_bits_data_lo_hi_148, memRequest_bits_data_lo_lo_148};
  wire [1:0]       memRequest_bits_data_hi_lo_148 = {_memRequest_bits_data_T_1991[140], _memRequest_bits_data_T_1798[140]};
  wire [1:0]       memRequest_bits_data_hi_hi_148 = {_memRequest_bits_data_T_2377[140], _memRequest_bits_data_T_2184[140]};
  wire [3:0]       memRequest_bits_data_hi_148 = {memRequest_bits_data_hi_hi_148, memRequest_bits_data_hi_lo_148};
  wire [1:0]       memRequest_bits_data_lo_lo_149 = {_memRequest_bits_data_T_1219[141], _memRequest_bits_data_T_1026[141]};
  wire [1:0]       memRequest_bits_data_lo_hi_149 = {_memRequest_bits_data_T_1605[141], _memRequest_bits_data_T_1412[141]};
  wire [3:0]       memRequest_bits_data_lo_149 = {memRequest_bits_data_lo_hi_149, memRequest_bits_data_lo_lo_149};
  wire [1:0]       memRequest_bits_data_hi_lo_149 = {_memRequest_bits_data_T_1991[141], _memRequest_bits_data_T_1798[141]};
  wire [1:0]       memRequest_bits_data_hi_hi_149 = {_memRequest_bits_data_T_2377[141], _memRequest_bits_data_T_2184[141]};
  wire [3:0]       memRequest_bits_data_hi_149 = {memRequest_bits_data_hi_hi_149, memRequest_bits_data_hi_lo_149};
  wire [1:0]       memRequest_bits_data_lo_lo_150 = {_memRequest_bits_data_T_1219[142], _memRequest_bits_data_T_1026[142]};
  wire [1:0]       memRequest_bits_data_lo_hi_150 = {_memRequest_bits_data_T_1605[142], _memRequest_bits_data_T_1412[142]};
  wire [3:0]       memRequest_bits_data_lo_150 = {memRequest_bits_data_lo_hi_150, memRequest_bits_data_lo_lo_150};
  wire [1:0]       memRequest_bits_data_hi_lo_150 = {_memRequest_bits_data_T_1991[142], _memRequest_bits_data_T_1798[142]};
  wire [1:0]       memRequest_bits_data_hi_hi_150 = {_memRequest_bits_data_T_2377[142], _memRequest_bits_data_T_2184[142]};
  wire [3:0]       memRequest_bits_data_hi_150 = {memRequest_bits_data_hi_hi_150, memRequest_bits_data_hi_lo_150};
  wire [1:0]       memRequest_bits_data_lo_lo_151 = {_memRequest_bits_data_T_1219[143], _memRequest_bits_data_T_1026[143]};
  wire [1:0]       memRequest_bits_data_lo_hi_151 = {_memRequest_bits_data_T_1605[143], _memRequest_bits_data_T_1412[143]};
  wire [3:0]       memRequest_bits_data_lo_151 = {memRequest_bits_data_lo_hi_151, memRequest_bits_data_lo_lo_151};
  wire [1:0]       memRequest_bits_data_hi_lo_151 = {_memRequest_bits_data_T_1991[143], _memRequest_bits_data_T_1798[143]};
  wire [1:0]       memRequest_bits_data_hi_hi_151 = {_memRequest_bits_data_T_2377[143], _memRequest_bits_data_T_2184[143]};
  wire [3:0]       memRequest_bits_data_hi_151 = {memRequest_bits_data_hi_hi_151, memRequest_bits_data_hi_lo_151};
  wire [1:0]       memRequest_bits_data_lo_lo_152 = {_memRequest_bits_data_T_1219[144], _memRequest_bits_data_T_1026[144]};
  wire [1:0]       memRequest_bits_data_lo_hi_152 = {_memRequest_bits_data_T_1605[144], _memRequest_bits_data_T_1412[144]};
  wire [3:0]       memRequest_bits_data_lo_152 = {memRequest_bits_data_lo_hi_152, memRequest_bits_data_lo_lo_152};
  wire [1:0]       memRequest_bits_data_hi_lo_152 = {_memRequest_bits_data_T_1991[144], _memRequest_bits_data_T_1798[144]};
  wire [1:0]       memRequest_bits_data_hi_hi_152 = {_memRequest_bits_data_T_2377[144], _memRequest_bits_data_T_2184[144]};
  wire [3:0]       memRequest_bits_data_hi_152 = {memRequest_bits_data_hi_hi_152, memRequest_bits_data_hi_lo_152};
  wire [1:0]       memRequest_bits_data_lo_lo_153 = {_memRequest_bits_data_T_1219[145], _memRequest_bits_data_T_1026[145]};
  wire [1:0]       memRequest_bits_data_lo_hi_153 = {_memRequest_bits_data_T_1605[145], _memRequest_bits_data_T_1412[145]};
  wire [3:0]       memRequest_bits_data_lo_153 = {memRequest_bits_data_lo_hi_153, memRequest_bits_data_lo_lo_153};
  wire [1:0]       memRequest_bits_data_hi_lo_153 = {_memRequest_bits_data_T_1991[145], _memRequest_bits_data_T_1798[145]};
  wire [1:0]       memRequest_bits_data_hi_hi_153 = {_memRequest_bits_data_T_2377[145], _memRequest_bits_data_T_2184[145]};
  wire [3:0]       memRequest_bits_data_hi_153 = {memRequest_bits_data_hi_hi_153, memRequest_bits_data_hi_lo_153};
  wire [1:0]       memRequest_bits_data_lo_lo_154 = {_memRequest_bits_data_T_1219[146], _memRequest_bits_data_T_1026[146]};
  wire [1:0]       memRequest_bits_data_lo_hi_154 = {_memRequest_bits_data_T_1605[146], _memRequest_bits_data_T_1412[146]};
  wire [3:0]       memRequest_bits_data_lo_154 = {memRequest_bits_data_lo_hi_154, memRequest_bits_data_lo_lo_154};
  wire [1:0]       memRequest_bits_data_hi_lo_154 = {_memRequest_bits_data_T_1991[146], _memRequest_bits_data_T_1798[146]};
  wire [1:0]       memRequest_bits_data_hi_hi_154 = {_memRequest_bits_data_T_2377[146], _memRequest_bits_data_T_2184[146]};
  wire [3:0]       memRequest_bits_data_hi_154 = {memRequest_bits_data_hi_hi_154, memRequest_bits_data_hi_lo_154};
  wire [1:0]       memRequest_bits_data_lo_lo_155 = {_memRequest_bits_data_T_1219[147], _memRequest_bits_data_T_1026[147]};
  wire [1:0]       memRequest_bits_data_lo_hi_155 = {_memRequest_bits_data_T_1605[147], _memRequest_bits_data_T_1412[147]};
  wire [3:0]       memRequest_bits_data_lo_155 = {memRequest_bits_data_lo_hi_155, memRequest_bits_data_lo_lo_155};
  wire [1:0]       memRequest_bits_data_hi_lo_155 = {_memRequest_bits_data_T_1991[147], _memRequest_bits_data_T_1798[147]};
  wire [1:0]       memRequest_bits_data_hi_hi_155 = {_memRequest_bits_data_T_2377[147], _memRequest_bits_data_T_2184[147]};
  wire [3:0]       memRequest_bits_data_hi_155 = {memRequest_bits_data_hi_hi_155, memRequest_bits_data_hi_lo_155};
  wire [1:0]       memRequest_bits_data_lo_lo_156 = {_memRequest_bits_data_T_1219[148], _memRequest_bits_data_T_1026[148]};
  wire [1:0]       memRequest_bits_data_lo_hi_156 = {_memRequest_bits_data_T_1605[148], _memRequest_bits_data_T_1412[148]};
  wire [3:0]       memRequest_bits_data_lo_156 = {memRequest_bits_data_lo_hi_156, memRequest_bits_data_lo_lo_156};
  wire [1:0]       memRequest_bits_data_hi_lo_156 = {_memRequest_bits_data_T_1991[148], _memRequest_bits_data_T_1798[148]};
  wire [1:0]       memRequest_bits_data_hi_hi_156 = {_memRequest_bits_data_T_2377[148], _memRequest_bits_data_T_2184[148]};
  wire [3:0]       memRequest_bits_data_hi_156 = {memRequest_bits_data_hi_hi_156, memRequest_bits_data_hi_lo_156};
  wire [1:0]       memRequest_bits_data_lo_lo_157 = {_memRequest_bits_data_T_1219[149], _memRequest_bits_data_T_1026[149]};
  wire [1:0]       memRequest_bits_data_lo_hi_157 = {_memRequest_bits_data_T_1605[149], _memRequest_bits_data_T_1412[149]};
  wire [3:0]       memRequest_bits_data_lo_157 = {memRequest_bits_data_lo_hi_157, memRequest_bits_data_lo_lo_157};
  wire [1:0]       memRequest_bits_data_hi_lo_157 = {_memRequest_bits_data_T_1991[149], _memRequest_bits_data_T_1798[149]};
  wire [1:0]       memRequest_bits_data_hi_hi_157 = {_memRequest_bits_data_T_2377[149], _memRequest_bits_data_T_2184[149]};
  wire [3:0]       memRequest_bits_data_hi_157 = {memRequest_bits_data_hi_hi_157, memRequest_bits_data_hi_lo_157};
  wire [1:0]       memRequest_bits_data_lo_lo_158 = {_memRequest_bits_data_T_1219[150], _memRequest_bits_data_T_1026[150]};
  wire [1:0]       memRequest_bits_data_lo_hi_158 = {_memRequest_bits_data_T_1605[150], _memRequest_bits_data_T_1412[150]};
  wire [3:0]       memRequest_bits_data_lo_158 = {memRequest_bits_data_lo_hi_158, memRequest_bits_data_lo_lo_158};
  wire [1:0]       memRequest_bits_data_hi_lo_158 = {_memRequest_bits_data_T_1991[150], _memRequest_bits_data_T_1798[150]};
  wire [1:0]       memRequest_bits_data_hi_hi_158 = {_memRequest_bits_data_T_2377[150], _memRequest_bits_data_T_2184[150]};
  wire [3:0]       memRequest_bits_data_hi_158 = {memRequest_bits_data_hi_hi_158, memRequest_bits_data_hi_lo_158};
  wire [1:0]       memRequest_bits_data_lo_lo_159 = {_memRequest_bits_data_T_1219[151], _memRequest_bits_data_T_1026[151]};
  wire [1:0]       memRequest_bits_data_lo_hi_159 = {_memRequest_bits_data_T_1605[151], _memRequest_bits_data_T_1412[151]};
  wire [3:0]       memRequest_bits_data_lo_159 = {memRequest_bits_data_lo_hi_159, memRequest_bits_data_lo_lo_159};
  wire [1:0]       memRequest_bits_data_hi_lo_159 = {_memRequest_bits_data_T_1991[151], _memRequest_bits_data_T_1798[151]};
  wire [1:0]       memRequest_bits_data_hi_hi_159 = {_memRequest_bits_data_T_2377[151], _memRequest_bits_data_T_2184[151]};
  wire [3:0]       memRequest_bits_data_hi_159 = {memRequest_bits_data_hi_hi_159, memRequest_bits_data_hi_lo_159};
  wire [1:0]       memRequest_bits_data_lo_lo_160 = {_memRequest_bits_data_T_1219[152], _memRequest_bits_data_T_1026[152]};
  wire [1:0]       memRequest_bits_data_lo_hi_160 = {_memRequest_bits_data_T_1605[152], _memRequest_bits_data_T_1412[152]};
  wire [3:0]       memRequest_bits_data_lo_160 = {memRequest_bits_data_lo_hi_160, memRequest_bits_data_lo_lo_160};
  wire [1:0]       memRequest_bits_data_hi_lo_160 = {_memRequest_bits_data_T_1991[152], _memRequest_bits_data_T_1798[152]};
  wire [1:0]       memRequest_bits_data_hi_hi_160 = {_memRequest_bits_data_T_2377[152], _memRequest_bits_data_T_2184[152]};
  wire [3:0]       memRequest_bits_data_hi_160 = {memRequest_bits_data_hi_hi_160, memRequest_bits_data_hi_lo_160};
  wire [1:0]       memRequest_bits_data_lo_lo_161 = {_memRequest_bits_data_T_1219[153], _memRequest_bits_data_T_1026[153]};
  wire [1:0]       memRequest_bits_data_lo_hi_161 = {_memRequest_bits_data_T_1605[153], _memRequest_bits_data_T_1412[153]};
  wire [3:0]       memRequest_bits_data_lo_161 = {memRequest_bits_data_lo_hi_161, memRequest_bits_data_lo_lo_161};
  wire [1:0]       memRequest_bits_data_hi_lo_161 = {_memRequest_bits_data_T_1991[153], _memRequest_bits_data_T_1798[153]};
  wire [1:0]       memRequest_bits_data_hi_hi_161 = {_memRequest_bits_data_T_2377[153], _memRequest_bits_data_T_2184[153]};
  wire [3:0]       memRequest_bits_data_hi_161 = {memRequest_bits_data_hi_hi_161, memRequest_bits_data_hi_lo_161};
  wire [1:0]       memRequest_bits_data_lo_lo_162 = {_memRequest_bits_data_T_1219[154], _memRequest_bits_data_T_1026[154]};
  wire [1:0]       memRequest_bits_data_lo_hi_162 = {_memRequest_bits_data_T_1605[154], _memRequest_bits_data_T_1412[154]};
  wire [3:0]       memRequest_bits_data_lo_162 = {memRequest_bits_data_lo_hi_162, memRequest_bits_data_lo_lo_162};
  wire [1:0]       memRequest_bits_data_hi_lo_162 = {_memRequest_bits_data_T_1991[154], _memRequest_bits_data_T_1798[154]};
  wire [1:0]       memRequest_bits_data_hi_hi_162 = {_memRequest_bits_data_T_2377[154], _memRequest_bits_data_T_2184[154]};
  wire [3:0]       memRequest_bits_data_hi_162 = {memRequest_bits_data_hi_hi_162, memRequest_bits_data_hi_lo_162};
  wire [1:0]       memRequest_bits_data_lo_lo_163 = {_memRequest_bits_data_T_1219[155], _memRequest_bits_data_T_1026[155]};
  wire [1:0]       memRequest_bits_data_lo_hi_163 = {_memRequest_bits_data_T_1605[155], _memRequest_bits_data_T_1412[155]};
  wire [3:0]       memRequest_bits_data_lo_163 = {memRequest_bits_data_lo_hi_163, memRequest_bits_data_lo_lo_163};
  wire [1:0]       memRequest_bits_data_hi_lo_163 = {_memRequest_bits_data_T_1991[155], _memRequest_bits_data_T_1798[155]};
  wire [1:0]       memRequest_bits_data_hi_hi_163 = {_memRequest_bits_data_T_2377[155], _memRequest_bits_data_T_2184[155]};
  wire [3:0]       memRequest_bits_data_hi_163 = {memRequest_bits_data_hi_hi_163, memRequest_bits_data_hi_lo_163};
  wire [1:0]       memRequest_bits_data_lo_lo_164 = {_memRequest_bits_data_T_1219[156], _memRequest_bits_data_T_1026[156]};
  wire [1:0]       memRequest_bits_data_lo_hi_164 = {_memRequest_bits_data_T_1605[156], _memRequest_bits_data_T_1412[156]};
  wire [3:0]       memRequest_bits_data_lo_164 = {memRequest_bits_data_lo_hi_164, memRequest_bits_data_lo_lo_164};
  wire [1:0]       memRequest_bits_data_hi_lo_164 = {_memRequest_bits_data_T_1991[156], _memRequest_bits_data_T_1798[156]};
  wire [1:0]       memRequest_bits_data_hi_hi_164 = {_memRequest_bits_data_T_2377[156], _memRequest_bits_data_T_2184[156]};
  wire [3:0]       memRequest_bits_data_hi_164 = {memRequest_bits_data_hi_hi_164, memRequest_bits_data_hi_lo_164};
  wire [1:0]       memRequest_bits_data_lo_lo_165 = {_memRequest_bits_data_T_1219[157], _memRequest_bits_data_T_1026[157]};
  wire [1:0]       memRequest_bits_data_lo_hi_165 = {_memRequest_bits_data_T_1605[157], _memRequest_bits_data_T_1412[157]};
  wire [3:0]       memRequest_bits_data_lo_165 = {memRequest_bits_data_lo_hi_165, memRequest_bits_data_lo_lo_165};
  wire [1:0]       memRequest_bits_data_hi_lo_165 = {_memRequest_bits_data_T_1991[157], _memRequest_bits_data_T_1798[157]};
  wire [1:0]       memRequest_bits_data_hi_hi_165 = {_memRequest_bits_data_T_2377[157], _memRequest_bits_data_T_2184[157]};
  wire [3:0]       memRequest_bits_data_hi_165 = {memRequest_bits_data_hi_hi_165, memRequest_bits_data_hi_lo_165};
  wire [1:0]       memRequest_bits_data_lo_lo_166 = {_memRequest_bits_data_T_1219[158], _memRequest_bits_data_T_1026[158]};
  wire [1:0]       memRequest_bits_data_lo_hi_166 = {_memRequest_bits_data_T_1605[158], _memRequest_bits_data_T_1412[158]};
  wire [3:0]       memRequest_bits_data_lo_166 = {memRequest_bits_data_lo_hi_166, memRequest_bits_data_lo_lo_166};
  wire [1:0]       memRequest_bits_data_hi_lo_166 = {_memRequest_bits_data_T_1991[158], _memRequest_bits_data_T_1798[158]};
  wire [1:0]       memRequest_bits_data_hi_hi_166 = {_memRequest_bits_data_T_2377[158], _memRequest_bits_data_T_2184[158]};
  wire [3:0]       memRequest_bits_data_hi_166 = {memRequest_bits_data_hi_hi_166, memRequest_bits_data_hi_lo_166};
  wire [1:0]       memRequest_bits_data_lo_lo_167 = {_memRequest_bits_data_T_1219[159], _memRequest_bits_data_T_1026[159]};
  wire [1:0]       memRequest_bits_data_lo_hi_167 = {_memRequest_bits_data_T_1605[159], _memRequest_bits_data_T_1412[159]};
  wire [3:0]       memRequest_bits_data_lo_167 = {memRequest_bits_data_lo_hi_167, memRequest_bits_data_lo_lo_167};
  wire [1:0]       memRequest_bits_data_hi_lo_167 = {_memRequest_bits_data_T_1991[159], _memRequest_bits_data_T_1798[159]};
  wire [1:0]       memRequest_bits_data_hi_hi_167 = {_memRequest_bits_data_T_2377[159], _memRequest_bits_data_T_2184[159]};
  wire [3:0]       memRequest_bits_data_hi_167 = {memRequest_bits_data_hi_hi_167, memRequest_bits_data_hi_lo_167};
  wire [1:0]       memRequest_bits_data_lo_lo_168 = {_memRequest_bits_data_T_1219[160], _memRequest_bits_data_T_1026[160]};
  wire [1:0]       memRequest_bits_data_lo_hi_168 = {_memRequest_bits_data_T_1605[160], _memRequest_bits_data_T_1412[160]};
  wire [3:0]       memRequest_bits_data_lo_168 = {memRequest_bits_data_lo_hi_168, memRequest_bits_data_lo_lo_168};
  wire [1:0]       memRequest_bits_data_hi_lo_168 = {_memRequest_bits_data_T_1991[160], _memRequest_bits_data_T_1798[160]};
  wire [1:0]       memRequest_bits_data_hi_hi_168 = {_memRequest_bits_data_T_2377[160], _memRequest_bits_data_T_2184[160]};
  wire [3:0]       memRequest_bits_data_hi_168 = {memRequest_bits_data_hi_hi_168, memRequest_bits_data_hi_lo_168};
  wire [1:0]       memRequest_bits_data_lo_lo_169 = {_memRequest_bits_data_T_1219[161], _memRequest_bits_data_T_1026[161]};
  wire [1:0]       memRequest_bits_data_lo_hi_169 = {_memRequest_bits_data_T_1605[161], _memRequest_bits_data_T_1412[161]};
  wire [3:0]       memRequest_bits_data_lo_169 = {memRequest_bits_data_lo_hi_169, memRequest_bits_data_lo_lo_169};
  wire [1:0]       memRequest_bits_data_hi_lo_169 = {_memRequest_bits_data_T_1991[161], _memRequest_bits_data_T_1798[161]};
  wire [1:0]       memRequest_bits_data_hi_hi_169 = {_memRequest_bits_data_T_2377[161], _memRequest_bits_data_T_2184[161]};
  wire [3:0]       memRequest_bits_data_hi_169 = {memRequest_bits_data_hi_hi_169, memRequest_bits_data_hi_lo_169};
  wire [1:0]       memRequest_bits_data_lo_lo_170 = {_memRequest_bits_data_T_1219[162], _memRequest_bits_data_T_1026[162]};
  wire [1:0]       memRequest_bits_data_lo_hi_170 = {_memRequest_bits_data_T_1605[162], _memRequest_bits_data_T_1412[162]};
  wire [3:0]       memRequest_bits_data_lo_170 = {memRequest_bits_data_lo_hi_170, memRequest_bits_data_lo_lo_170};
  wire [1:0]       memRequest_bits_data_hi_lo_170 = {_memRequest_bits_data_T_1991[162], _memRequest_bits_data_T_1798[162]};
  wire [1:0]       memRequest_bits_data_hi_hi_170 = {_memRequest_bits_data_T_2377[162], _memRequest_bits_data_T_2184[162]};
  wire [3:0]       memRequest_bits_data_hi_170 = {memRequest_bits_data_hi_hi_170, memRequest_bits_data_hi_lo_170};
  wire [1:0]       memRequest_bits_data_lo_lo_171 = {_memRequest_bits_data_T_1219[163], _memRequest_bits_data_T_1026[163]};
  wire [1:0]       memRequest_bits_data_lo_hi_171 = {_memRequest_bits_data_T_1605[163], _memRequest_bits_data_T_1412[163]};
  wire [3:0]       memRequest_bits_data_lo_171 = {memRequest_bits_data_lo_hi_171, memRequest_bits_data_lo_lo_171};
  wire [1:0]       memRequest_bits_data_hi_lo_171 = {_memRequest_bits_data_T_1991[163], _memRequest_bits_data_T_1798[163]};
  wire [1:0]       memRequest_bits_data_hi_hi_171 = {_memRequest_bits_data_T_2377[163], _memRequest_bits_data_T_2184[163]};
  wire [3:0]       memRequest_bits_data_hi_171 = {memRequest_bits_data_hi_hi_171, memRequest_bits_data_hi_lo_171};
  wire [1:0]       memRequest_bits_data_lo_lo_172 = {_memRequest_bits_data_T_1219[164], _memRequest_bits_data_T_1026[164]};
  wire [1:0]       memRequest_bits_data_lo_hi_172 = {_memRequest_bits_data_T_1605[164], _memRequest_bits_data_T_1412[164]};
  wire [3:0]       memRequest_bits_data_lo_172 = {memRequest_bits_data_lo_hi_172, memRequest_bits_data_lo_lo_172};
  wire [1:0]       memRequest_bits_data_hi_lo_172 = {_memRequest_bits_data_T_1991[164], _memRequest_bits_data_T_1798[164]};
  wire [1:0]       memRequest_bits_data_hi_hi_172 = {_memRequest_bits_data_T_2377[164], _memRequest_bits_data_T_2184[164]};
  wire [3:0]       memRequest_bits_data_hi_172 = {memRequest_bits_data_hi_hi_172, memRequest_bits_data_hi_lo_172};
  wire [1:0]       memRequest_bits_data_lo_lo_173 = {_memRequest_bits_data_T_1219[165], _memRequest_bits_data_T_1026[165]};
  wire [1:0]       memRequest_bits_data_lo_hi_173 = {_memRequest_bits_data_T_1605[165], _memRequest_bits_data_T_1412[165]};
  wire [3:0]       memRequest_bits_data_lo_173 = {memRequest_bits_data_lo_hi_173, memRequest_bits_data_lo_lo_173};
  wire [1:0]       memRequest_bits_data_hi_lo_173 = {_memRequest_bits_data_T_1991[165], _memRequest_bits_data_T_1798[165]};
  wire [1:0]       memRequest_bits_data_hi_hi_173 = {_memRequest_bits_data_T_2377[165], _memRequest_bits_data_T_2184[165]};
  wire [3:0]       memRequest_bits_data_hi_173 = {memRequest_bits_data_hi_hi_173, memRequest_bits_data_hi_lo_173};
  wire [1:0]       memRequest_bits_data_lo_lo_174 = {_memRequest_bits_data_T_1219[166], _memRequest_bits_data_T_1026[166]};
  wire [1:0]       memRequest_bits_data_lo_hi_174 = {_memRequest_bits_data_T_1605[166], _memRequest_bits_data_T_1412[166]};
  wire [3:0]       memRequest_bits_data_lo_174 = {memRequest_bits_data_lo_hi_174, memRequest_bits_data_lo_lo_174};
  wire [1:0]       memRequest_bits_data_hi_lo_174 = {_memRequest_bits_data_T_1991[166], _memRequest_bits_data_T_1798[166]};
  wire [1:0]       memRequest_bits_data_hi_hi_174 = {_memRequest_bits_data_T_2377[166], _memRequest_bits_data_T_2184[166]};
  wire [3:0]       memRequest_bits_data_hi_174 = {memRequest_bits_data_hi_hi_174, memRequest_bits_data_hi_lo_174};
  wire [1:0]       memRequest_bits_data_lo_lo_175 = {_memRequest_bits_data_T_1219[167], _memRequest_bits_data_T_1026[167]};
  wire [1:0]       memRequest_bits_data_lo_hi_175 = {_memRequest_bits_data_T_1605[167], _memRequest_bits_data_T_1412[167]};
  wire [3:0]       memRequest_bits_data_lo_175 = {memRequest_bits_data_lo_hi_175, memRequest_bits_data_lo_lo_175};
  wire [1:0]       memRequest_bits_data_hi_lo_175 = {_memRequest_bits_data_T_1991[167], _memRequest_bits_data_T_1798[167]};
  wire [1:0]       memRequest_bits_data_hi_hi_175 = {_memRequest_bits_data_T_2377[167], _memRequest_bits_data_T_2184[167]};
  wire [3:0]       memRequest_bits_data_hi_175 = {memRequest_bits_data_hi_hi_175, memRequest_bits_data_hi_lo_175};
  wire [1:0]       memRequest_bits_data_lo_lo_176 = {_memRequest_bits_data_T_1219[168], _memRequest_bits_data_T_1026[168]};
  wire [1:0]       memRequest_bits_data_lo_hi_176 = {_memRequest_bits_data_T_1605[168], _memRequest_bits_data_T_1412[168]};
  wire [3:0]       memRequest_bits_data_lo_176 = {memRequest_bits_data_lo_hi_176, memRequest_bits_data_lo_lo_176};
  wire [1:0]       memRequest_bits_data_hi_lo_176 = {_memRequest_bits_data_T_1991[168], _memRequest_bits_data_T_1798[168]};
  wire [1:0]       memRequest_bits_data_hi_hi_176 = {_memRequest_bits_data_T_2377[168], _memRequest_bits_data_T_2184[168]};
  wire [3:0]       memRequest_bits_data_hi_176 = {memRequest_bits_data_hi_hi_176, memRequest_bits_data_hi_lo_176};
  wire [1:0]       memRequest_bits_data_lo_lo_177 = {_memRequest_bits_data_T_1219[169], _memRequest_bits_data_T_1026[169]};
  wire [1:0]       memRequest_bits_data_lo_hi_177 = {_memRequest_bits_data_T_1605[169], _memRequest_bits_data_T_1412[169]};
  wire [3:0]       memRequest_bits_data_lo_177 = {memRequest_bits_data_lo_hi_177, memRequest_bits_data_lo_lo_177};
  wire [1:0]       memRequest_bits_data_hi_lo_177 = {_memRequest_bits_data_T_1991[169], _memRequest_bits_data_T_1798[169]};
  wire [1:0]       memRequest_bits_data_hi_hi_177 = {_memRequest_bits_data_T_2377[169], _memRequest_bits_data_T_2184[169]};
  wire [3:0]       memRequest_bits_data_hi_177 = {memRequest_bits_data_hi_hi_177, memRequest_bits_data_hi_lo_177};
  wire [1:0]       memRequest_bits_data_lo_lo_178 = {_memRequest_bits_data_T_1219[170], _memRequest_bits_data_T_1026[170]};
  wire [1:0]       memRequest_bits_data_lo_hi_178 = {_memRequest_bits_data_T_1605[170], _memRequest_bits_data_T_1412[170]};
  wire [3:0]       memRequest_bits_data_lo_178 = {memRequest_bits_data_lo_hi_178, memRequest_bits_data_lo_lo_178};
  wire [1:0]       memRequest_bits_data_hi_lo_178 = {_memRequest_bits_data_T_1991[170], _memRequest_bits_data_T_1798[170]};
  wire [1:0]       memRequest_bits_data_hi_hi_178 = {_memRequest_bits_data_T_2377[170], _memRequest_bits_data_T_2184[170]};
  wire [3:0]       memRequest_bits_data_hi_178 = {memRequest_bits_data_hi_hi_178, memRequest_bits_data_hi_lo_178};
  wire [1:0]       memRequest_bits_data_lo_lo_179 = {_memRequest_bits_data_T_1219[171], _memRequest_bits_data_T_1026[171]};
  wire [1:0]       memRequest_bits_data_lo_hi_179 = {_memRequest_bits_data_T_1605[171], _memRequest_bits_data_T_1412[171]};
  wire [3:0]       memRequest_bits_data_lo_179 = {memRequest_bits_data_lo_hi_179, memRequest_bits_data_lo_lo_179};
  wire [1:0]       memRequest_bits_data_hi_lo_179 = {_memRequest_bits_data_T_1991[171], _memRequest_bits_data_T_1798[171]};
  wire [1:0]       memRequest_bits_data_hi_hi_179 = {_memRequest_bits_data_T_2377[171], _memRequest_bits_data_T_2184[171]};
  wire [3:0]       memRequest_bits_data_hi_179 = {memRequest_bits_data_hi_hi_179, memRequest_bits_data_hi_lo_179};
  wire [1:0]       memRequest_bits_data_lo_lo_180 = {_memRequest_bits_data_T_1219[172], _memRequest_bits_data_T_1026[172]};
  wire [1:0]       memRequest_bits_data_lo_hi_180 = {_memRequest_bits_data_T_1605[172], _memRequest_bits_data_T_1412[172]};
  wire [3:0]       memRequest_bits_data_lo_180 = {memRequest_bits_data_lo_hi_180, memRequest_bits_data_lo_lo_180};
  wire [1:0]       memRequest_bits_data_hi_lo_180 = {_memRequest_bits_data_T_1991[172], _memRequest_bits_data_T_1798[172]};
  wire [1:0]       memRequest_bits_data_hi_hi_180 = {_memRequest_bits_data_T_2377[172], _memRequest_bits_data_T_2184[172]};
  wire [3:0]       memRequest_bits_data_hi_180 = {memRequest_bits_data_hi_hi_180, memRequest_bits_data_hi_lo_180};
  wire [1:0]       memRequest_bits_data_lo_lo_181 = {_memRequest_bits_data_T_1219[173], _memRequest_bits_data_T_1026[173]};
  wire [1:0]       memRequest_bits_data_lo_hi_181 = {_memRequest_bits_data_T_1605[173], _memRequest_bits_data_T_1412[173]};
  wire [3:0]       memRequest_bits_data_lo_181 = {memRequest_bits_data_lo_hi_181, memRequest_bits_data_lo_lo_181};
  wire [1:0]       memRequest_bits_data_hi_lo_181 = {_memRequest_bits_data_T_1991[173], _memRequest_bits_data_T_1798[173]};
  wire [1:0]       memRequest_bits_data_hi_hi_181 = {_memRequest_bits_data_T_2377[173], _memRequest_bits_data_T_2184[173]};
  wire [3:0]       memRequest_bits_data_hi_181 = {memRequest_bits_data_hi_hi_181, memRequest_bits_data_hi_lo_181};
  wire [1:0]       memRequest_bits_data_lo_lo_182 = {_memRequest_bits_data_T_1219[174], _memRequest_bits_data_T_1026[174]};
  wire [1:0]       memRequest_bits_data_lo_hi_182 = {_memRequest_bits_data_T_1605[174], _memRequest_bits_data_T_1412[174]};
  wire [3:0]       memRequest_bits_data_lo_182 = {memRequest_bits_data_lo_hi_182, memRequest_bits_data_lo_lo_182};
  wire [1:0]       memRequest_bits_data_hi_lo_182 = {_memRequest_bits_data_T_1991[174], _memRequest_bits_data_T_1798[174]};
  wire [1:0]       memRequest_bits_data_hi_hi_182 = {_memRequest_bits_data_T_2377[174], _memRequest_bits_data_T_2184[174]};
  wire [3:0]       memRequest_bits_data_hi_182 = {memRequest_bits_data_hi_hi_182, memRequest_bits_data_hi_lo_182};
  wire [1:0]       memRequest_bits_data_lo_lo_183 = {_memRequest_bits_data_T_1219[175], _memRequest_bits_data_T_1026[175]};
  wire [1:0]       memRequest_bits_data_lo_hi_183 = {_memRequest_bits_data_T_1605[175], _memRequest_bits_data_T_1412[175]};
  wire [3:0]       memRequest_bits_data_lo_183 = {memRequest_bits_data_lo_hi_183, memRequest_bits_data_lo_lo_183};
  wire [1:0]       memRequest_bits_data_hi_lo_183 = {_memRequest_bits_data_T_1991[175], _memRequest_bits_data_T_1798[175]};
  wire [1:0]       memRequest_bits_data_hi_hi_183 = {_memRequest_bits_data_T_2377[175], _memRequest_bits_data_T_2184[175]};
  wire [3:0]       memRequest_bits_data_hi_183 = {memRequest_bits_data_hi_hi_183, memRequest_bits_data_hi_lo_183};
  wire [1:0]       memRequest_bits_data_lo_lo_184 = {_memRequest_bits_data_T_1219[176], _memRequest_bits_data_T_1026[176]};
  wire [1:0]       memRequest_bits_data_lo_hi_184 = {_memRequest_bits_data_T_1605[176], _memRequest_bits_data_T_1412[176]};
  wire [3:0]       memRequest_bits_data_lo_184 = {memRequest_bits_data_lo_hi_184, memRequest_bits_data_lo_lo_184};
  wire [1:0]       memRequest_bits_data_hi_lo_184 = {_memRequest_bits_data_T_1991[176], _memRequest_bits_data_T_1798[176]};
  wire [1:0]       memRequest_bits_data_hi_hi_184 = {_memRequest_bits_data_T_2377[176], _memRequest_bits_data_T_2184[176]};
  wire [3:0]       memRequest_bits_data_hi_184 = {memRequest_bits_data_hi_hi_184, memRequest_bits_data_hi_lo_184};
  wire [1:0]       memRequest_bits_data_lo_lo_185 = {_memRequest_bits_data_T_1219[177], _memRequest_bits_data_T_1026[177]};
  wire [1:0]       memRequest_bits_data_lo_hi_185 = {_memRequest_bits_data_T_1605[177], _memRequest_bits_data_T_1412[177]};
  wire [3:0]       memRequest_bits_data_lo_185 = {memRequest_bits_data_lo_hi_185, memRequest_bits_data_lo_lo_185};
  wire [1:0]       memRequest_bits_data_hi_lo_185 = {_memRequest_bits_data_T_1991[177], _memRequest_bits_data_T_1798[177]};
  wire [1:0]       memRequest_bits_data_hi_hi_185 = {_memRequest_bits_data_T_2377[177], _memRequest_bits_data_T_2184[177]};
  wire [3:0]       memRequest_bits_data_hi_185 = {memRequest_bits_data_hi_hi_185, memRequest_bits_data_hi_lo_185};
  wire [1:0]       memRequest_bits_data_lo_lo_186 = {_memRequest_bits_data_T_1219[178], _memRequest_bits_data_T_1026[178]};
  wire [1:0]       memRequest_bits_data_lo_hi_186 = {_memRequest_bits_data_T_1605[178], _memRequest_bits_data_T_1412[178]};
  wire [3:0]       memRequest_bits_data_lo_186 = {memRequest_bits_data_lo_hi_186, memRequest_bits_data_lo_lo_186};
  wire [1:0]       memRequest_bits_data_hi_lo_186 = {_memRequest_bits_data_T_1991[178], _memRequest_bits_data_T_1798[178]};
  wire [1:0]       memRequest_bits_data_hi_hi_186 = {_memRequest_bits_data_T_2377[178], _memRequest_bits_data_T_2184[178]};
  wire [3:0]       memRequest_bits_data_hi_186 = {memRequest_bits_data_hi_hi_186, memRequest_bits_data_hi_lo_186};
  wire [1:0]       memRequest_bits_data_lo_lo_187 = {_memRequest_bits_data_T_1219[179], _memRequest_bits_data_T_1026[179]};
  wire [1:0]       memRequest_bits_data_lo_hi_187 = {_memRequest_bits_data_T_1605[179], _memRequest_bits_data_T_1412[179]};
  wire [3:0]       memRequest_bits_data_lo_187 = {memRequest_bits_data_lo_hi_187, memRequest_bits_data_lo_lo_187};
  wire [1:0]       memRequest_bits_data_hi_lo_187 = {_memRequest_bits_data_T_1991[179], _memRequest_bits_data_T_1798[179]};
  wire [1:0]       memRequest_bits_data_hi_hi_187 = {_memRequest_bits_data_T_2377[179], _memRequest_bits_data_T_2184[179]};
  wire [3:0]       memRequest_bits_data_hi_187 = {memRequest_bits_data_hi_hi_187, memRequest_bits_data_hi_lo_187};
  wire [1:0]       memRequest_bits_data_lo_lo_188 = {_memRequest_bits_data_T_1219[180], _memRequest_bits_data_T_1026[180]};
  wire [1:0]       memRequest_bits_data_lo_hi_188 = {_memRequest_bits_data_T_1605[180], _memRequest_bits_data_T_1412[180]};
  wire [3:0]       memRequest_bits_data_lo_188 = {memRequest_bits_data_lo_hi_188, memRequest_bits_data_lo_lo_188};
  wire [1:0]       memRequest_bits_data_hi_lo_188 = {_memRequest_bits_data_T_1991[180], _memRequest_bits_data_T_1798[180]};
  wire [1:0]       memRequest_bits_data_hi_hi_188 = {_memRequest_bits_data_T_2377[180], _memRequest_bits_data_T_2184[180]};
  wire [3:0]       memRequest_bits_data_hi_188 = {memRequest_bits_data_hi_hi_188, memRequest_bits_data_hi_lo_188};
  wire [1:0]       memRequest_bits_data_lo_lo_189 = {_memRequest_bits_data_T_1219[181], _memRequest_bits_data_T_1026[181]};
  wire [1:0]       memRequest_bits_data_lo_hi_189 = {_memRequest_bits_data_T_1605[181], _memRequest_bits_data_T_1412[181]};
  wire [3:0]       memRequest_bits_data_lo_189 = {memRequest_bits_data_lo_hi_189, memRequest_bits_data_lo_lo_189};
  wire [1:0]       memRequest_bits_data_hi_lo_189 = {_memRequest_bits_data_T_1991[181], _memRequest_bits_data_T_1798[181]};
  wire [1:0]       memRequest_bits_data_hi_hi_189 = {_memRequest_bits_data_T_2377[181], _memRequest_bits_data_T_2184[181]};
  wire [3:0]       memRequest_bits_data_hi_189 = {memRequest_bits_data_hi_hi_189, memRequest_bits_data_hi_lo_189};
  wire [1:0]       memRequest_bits_data_lo_lo_190 = {_memRequest_bits_data_T_1219[182], _memRequest_bits_data_T_1026[182]};
  wire [1:0]       memRequest_bits_data_lo_hi_190 = {_memRequest_bits_data_T_1605[182], _memRequest_bits_data_T_1412[182]};
  wire [3:0]       memRequest_bits_data_lo_190 = {memRequest_bits_data_lo_hi_190, memRequest_bits_data_lo_lo_190};
  wire [1:0]       memRequest_bits_data_hi_lo_190 = {_memRequest_bits_data_T_1991[182], _memRequest_bits_data_T_1798[182]};
  wire [1:0]       memRequest_bits_data_hi_hi_190 = {_memRequest_bits_data_T_2377[182], _memRequest_bits_data_T_2184[182]};
  wire [3:0]       memRequest_bits_data_hi_190 = {memRequest_bits_data_hi_hi_190, memRequest_bits_data_hi_lo_190};
  wire [1:0]       memRequest_bits_data_lo_lo_191 = {_memRequest_bits_data_T_1219[183], _memRequest_bits_data_T_1026[183]};
  wire [1:0]       memRequest_bits_data_lo_hi_191 = {_memRequest_bits_data_T_1605[183], _memRequest_bits_data_T_1412[183]};
  wire [3:0]       memRequest_bits_data_lo_191 = {memRequest_bits_data_lo_hi_191, memRequest_bits_data_lo_lo_191};
  wire [1:0]       memRequest_bits_data_hi_lo_191 = {_memRequest_bits_data_T_1991[183], _memRequest_bits_data_T_1798[183]};
  wire [1:0]       memRequest_bits_data_hi_hi_191 = {_memRequest_bits_data_T_2377[183], _memRequest_bits_data_T_2184[183]};
  wire [3:0]       memRequest_bits_data_hi_191 = {memRequest_bits_data_hi_hi_191, memRequest_bits_data_hi_lo_191};
  wire [1:0]       memRequest_bits_data_lo_lo_192 = {_memRequest_bits_data_T_1219[184], _memRequest_bits_data_T_1026[184]};
  wire [1:0]       memRequest_bits_data_lo_hi_192 = {_memRequest_bits_data_T_1605[184], _memRequest_bits_data_T_1412[184]};
  wire [3:0]       memRequest_bits_data_lo_192 = {memRequest_bits_data_lo_hi_192, memRequest_bits_data_lo_lo_192};
  wire [1:0]       memRequest_bits_data_hi_lo_192 = {_memRequest_bits_data_T_1991[184], _memRequest_bits_data_T_1798[184]};
  wire [1:0]       memRequest_bits_data_hi_hi_192 = {_memRequest_bits_data_T_2377[184], _memRequest_bits_data_T_2184[184]};
  wire [3:0]       memRequest_bits_data_hi_192 = {memRequest_bits_data_hi_hi_192, memRequest_bits_data_hi_lo_192};
  wire [1:0]       memRequest_bits_data_lo_lo_193 = {_memRequest_bits_data_T_1219[185], _memRequest_bits_data_T_1026[185]};
  wire [1:0]       memRequest_bits_data_lo_hi_193 = {_memRequest_bits_data_T_1605[185], _memRequest_bits_data_T_1412[185]};
  wire [3:0]       memRequest_bits_data_lo_193 = {memRequest_bits_data_lo_hi_193, memRequest_bits_data_lo_lo_193};
  wire [1:0]       memRequest_bits_data_hi_lo_193 = {_memRequest_bits_data_T_1991[185], _memRequest_bits_data_T_1798[185]};
  wire [1:0]       memRequest_bits_data_hi_hi_193 = {_memRequest_bits_data_T_2377[185], _memRequest_bits_data_T_2184[185]};
  wire [3:0]       memRequest_bits_data_hi_193 = {memRequest_bits_data_hi_hi_193, memRequest_bits_data_hi_lo_193};
  wire [1:0]       memRequest_bits_data_lo_lo_194 = {_memRequest_bits_data_T_1219[186], _memRequest_bits_data_T_1026[186]};
  wire [1:0]       memRequest_bits_data_lo_hi_194 = {_memRequest_bits_data_T_1605[186], _memRequest_bits_data_T_1412[186]};
  wire [3:0]       memRequest_bits_data_lo_194 = {memRequest_bits_data_lo_hi_194, memRequest_bits_data_lo_lo_194};
  wire [1:0]       memRequest_bits_data_hi_lo_194 = {_memRequest_bits_data_T_1991[186], _memRequest_bits_data_T_1798[186]};
  wire [1:0]       memRequest_bits_data_hi_hi_194 = {_memRequest_bits_data_T_2377[186], _memRequest_bits_data_T_2184[186]};
  wire [3:0]       memRequest_bits_data_hi_194 = {memRequest_bits_data_hi_hi_194, memRequest_bits_data_hi_lo_194};
  wire [1:0]       memRequest_bits_data_lo_lo_195 = {_memRequest_bits_data_T_1219[187], _memRequest_bits_data_T_1026[187]};
  wire [1:0]       memRequest_bits_data_lo_hi_195 = {_memRequest_bits_data_T_1605[187], _memRequest_bits_data_T_1412[187]};
  wire [3:0]       memRequest_bits_data_lo_195 = {memRequest_bits_data_lo_hi_195, memRequest_bits_data_lo_lo_195};
  wire [1:0]       memRequest_bits_data_hi_lo_195 = {_memRequest_bits_data_T_1991[187], _memRequest_bits_data_T_1798[187]};
  wire [1:0]       memRequest_bits_data_hi_hi_195 = {_memRequest_bits_data_T_2377[187], _memRequest_bits_data_T_2184[187]};
  wire [3:0]       memRequest_bits_data_hi_195 = {memRequest_bits_data_hi_hi_195, memRequest_bits_data_hi_lo_195};
  wire [1:0]       memRequest_bits_data_lo_lo_196 = {_memRequest_bits_data_T_1219[188], _memRequest_bits_data_T_1026[188]};
  wire [1:0]       memRequest_bits_data_lo_hi_196 = {_memRequest_bits_data_T_1605[188], _memRequest_bits_data_T_1412[188]};
  wire [3:0]       memRequest_bits_data_lo_196 = {memRequest_bits_data_lo_hi_196, memRequest_bits_data_lo_lo_196};
  wire [1:0]       memRequest_bits_data_hi_lo_196 = {_memRequest_bits_data_T_1991[188], _memRequest_bits_data_T_1798[188]};
  wire [1:0]       memRequest_bits_data_hi_hi_196 = {_memRequest_bits_data_T_2377[188], _memRequest_bits_data_T_2184[188]};
  wire [3:0]       memRequest_bits_data_hi_196 = {memRequest_bits_data_hi_hi_196, memRequest_bits_data_hi_lo_196};
  wire [1:0]       memRequest_bits_data_lo_lo_197 = {_memRequest_bits_data_T_1219[189], _memRequest_bits_data_T_1026[189]};
  wire [1:0]       memRequest_bits_data_lo_hi_197 = {_memRequest_bits_data_T_1605[189], _memRequest_bits_data_T_1412[189]};
  wire [3:0]       memRequest_bits_data_lo_197 = {memRequest_bits_data_lo_hi_197, memRequest_bits_data_lo_lo_197};
  wire [1:0]       memRequest_bits_data_hi_lo_197 = {_memRequest_bits_data_T_1991[189], _memRequest_bits_data_T_1798[189]};
  wire [1:0]       memRequest_bits_data_hi_hi_197 = {_memRequest_bits_data_T_2377[189], _memRequest_bits_data_T_2184[189]};
  wire [3:0]       memRequest_bits_data_hi_197 = {memRequest_bits_data_hi_hi_197, memRequest_bits_data_hi_lo_197};
  wire [1:0]       memRequest_bits_data_lo_lo_198 = {_memRequest_bits_data_T_1219[190], _memRequest_bits_data_T_1026[190]};
  wire [1:0]       memRequest_bits_data_lo_hi_198 = {_memRequest_bits_data_T_1605[190], _memRequest_bits_data_T_1412[190]};
  wire [3:0]       memRequest_bits_data_lo_198 = {memRequest_bits_data_lo_hi_198, memRequest_bits_data_lo_lo_198};
  wire [1:0]       memRequest_bits_data_hi_lo_198 = {_memRequest_bits_data_T_1991[190], _memRequest_bits_data_T_1798[190]};
  wire [1:0]       memRequest_bits_data_hi_hi_198 = {_memRequest_bits_data_T_2377[190], _memRequest_bits_data_T_2184[190]};
  wire [3:0]       memRequest_bits_data_hi_198 = {memRequest_bits_data_hi_hi_198, memRequest_bits_data_hi_lo_198};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_9, memRequest_bits_data_lo_9, memRequest_bits_data_hi_8, memRequest_bits_data_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_12, memRequest_bits_data_lo_12, memRequest_bits_data_hi_11, memRequest_bits_data_lo_11};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_10, memRequest_bits_data_lo_10};
  wire [39:0]      memRequest_bits_data_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_15, memRequest_bits_data_lo_15, memRequest_bits_data_hi_14, memRequest_bits_data_lo_14};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_13, memRequest_bits_data_lo_13};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_18, memRequest_bits_data_lo_18, memRequest_bits_data_hi_17, memRequest_bits_data_lo_17};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_16, memRequest_bits_data_lo_16};
  wire [47:0]      memRequest_bits_data_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_lo_hi_lo_8};
  wire [87:0]      memRequest_bits_data_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_21, memRequest_bits_data_lo_21, memRequest_bits_data_hi_20, memRequest_bits_data_lo_20};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_19, memRequest_bits_data_lo_19};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_24, memRequest_bits_data_lo_24, memRequest_bits_data_hi_23, memRequest_bits_data_lo_23};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_22, memRequest_bits_data_lo_22};
  wire [47:0]      memRequest_bits_data_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_27, memRequest_bits_data_lo_27, memRequest_bits_data_hi_26, memRequest_bits_data_lo_26};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_25, memRequest_bits_data_lo_25};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_30, memRequest_bits_data_lo_30, memRequest_bits_data_hi_29, memRequest_bits_data_lo_29};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_28, memRequest_bits_data_lo_28};
  wire [47:0]      memRequest_bits_data_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_8};
  wire [183:0]     memRequest_bits_data_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_33, memRequest_bits_data_lo_33, memRequest_bits_data_hi_32, memRequest_bits_data_lo_32};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_31, memRequest_bits_data_lo_31};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_36, memRequest_bits_data_lo_36, memRequest_bits_data_hi_35, memRequest_bits_data_lo_35};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_34, memRequest_bits_data_lo_34};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_39, memRequest_bits_data_lo_39, memRequest_bits_data_hi_38, memRequest_bits_data_lo_38};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_37, memRequest_bits_data_lo_37};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_42, memRequest_bits_data_lo_42, memRequest_bits_data_hi_41, memRequest_bits_data_lo_41};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_40, memRequest_bits_data_lo_40};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_45, memRequest_bits_data_lo_45, memRequest_bits_data_hi_44, memRequest_bits_data_lo_44};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_43, memRequest_bits_data_lo_43};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_48, memRequest_bits_data_lo_48, memRequest_bits_data_hi_47, memRequest_bits_data_lo_47};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_46, memRequest_bits_data_lo_46};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_51, memRequest_bits_data_lo_51, memRequest_bits_data_hi_50, memRequest_bits_data_lo_50};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_49, memRequest_bits_data_lo_49};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_54, memRequest_bits_data_lo_54, memRequest_bits_data_hi_53, memRequest_bits_data_lo_53};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_52, memRequest_bits_data_lo_52};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_8};
  wire [375:0]     memRequest_bits_data_lo_lo_199 = {memRequest_bits_data_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_57, memRequest_bits_data_lo_57, memRequest_bits_data_hi_56, memRequest_bits_data_lo_56};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_55, memRequest_bits_data_lo_55};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_60, memRequest_bits_data_lo_60, memRequest_bits_data_hi_59, memRequest_bits_data_lo_59};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_58, memRequest_bits_data_lo_58};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_63, memRequest_bits_data_lo_63, memRequest_bits_data_hi_62, memRequest_bits_data_lo_62};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_61, memRequest_bits_data_lo_61};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_66, memRequest_bits_data_lo_66, memRequest_bits_data_hi_65, memRequest_bits_data_lo_65};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_64, memRequest_bits_data_lo_64};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_69, memRequest_bits_data_lo_69, memRequest_bits_data_hi_68, memRequest_bits_data_lo_68};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_67, memRequest_bits_data_lo_67};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_72, memRequest_bits_data_lo_72, memRequest_bits_data_hi_71, memRequest_bits_data_lo_71};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_70, memRequest_bits_data_lo_70};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_75, memRequest_bits_data_lo_75, memRequest_bits_data_hi_74, memRequest_bits_data_lo_74};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_73, memRequest_bits_data_lo_73};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_78, memRequest_bits_data_lo_78, memRequest_bits_data_hi_77, memRequest_bits_data_lo_77};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_76, memRequest_bits_data_lo_76};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_8};
  wire [191:0]     memRequest_bits_data_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_81, memRequest_bits_data_lo_81, memRequest_bits_data_hi_80, memRequest_bits_data_lo_80};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_79, memRequest_bits_data_lo_79};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_84, memRequest_bits_data_lo_84, memRequest_bits_data_hi_83, memRequest_bits_data_lo_83};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_82, memRequest_bits_data_lo_82};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_87, memRequest_bits_data_lo_87, memRequest_bits_data_hi_86, memRequest_bits_data_lo_86};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_85, memRequest_bits_data_lo_85};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_90, memRequest_bits_data_lo_90, memRequest_bits_data_hi_89, memRequest_bits_data_lo_89};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_88, memRequest_bits_data_lo_88};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_93, memRequest_bits_data_lo_93, memRequest_bits_data_hi_92, memRequest_bits_data_lo_92};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_91, memRequest_bits_data_lo_91};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_96, memRequest_bits_data_lo_96, memRequest_bits_data_hi_95, memRequest_bits_data_lo_95};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_94, memRequest_bits_data_lo_94};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_99, memRequest_bits_data_lo_99, memRequest_bits_data_hi_98, memRequest_bits_data_lo_98};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_97, memRequest_bits_data_lo_97};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_102, memRequest_bits_data_lo_102, memRequest_bits_data_hi_101, memRequest_bits_data_lo_101};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_100, memRequest_bits_data_lo_100};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_8};
  wire [383:0]     memRequest_bits_data_lo_hi_199 = {memRequest_bits_data_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_8};
  wire [759:0]     memRequest_bits_data_lo_199 = {memRequest_bits_data_lo_hi_199, memRequest_bits_data_lo_lo_199};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_105, memRequest_bits_data_lo_105, memRequest_bits_data_hi_104, memRequest_bits_data_lo_104};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi, memRequest_bits_data_hi_103, memRequest_bits_data_lo_103};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_108, memRequest_bits_data_lo_108, memRequest_bits_data_hi_107, memRequest_bits_data_lo_107};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_106, memRequest_bits_data_lo_106};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_111, memRequest_bits_data_lo_111, memRequest_bits_data_hi_110, memRequest_bits_data_lo_110};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_109, memRequest_bits_data_lo_109};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_114, memRequest_bits_data_lo_114, memRequest_bits_data_hi_113, memRequest_bits_data_lo_113};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_112, memRequest_bits_data_lo_112};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_117, memRequest_bits_data_lo_117, memRequest_bits_data_hi_116, memRequest_bits_data_lo_116};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_115, memRequest_bits_data_lo_115};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_120, memRequest_bits_data_lo_120, memRequest_bits_data_hi_119, memRequest_bits_data_lo_119};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_118, memRequest_bits_data_lo_118};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_123, memRequest_bits_data_lo_123, memRequest_bits_data_hi_122, memRequest_bits_data_lo_122};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_121, memRequest_bits_data_lo_121};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_126, memRequest_bits_data_lo_126, memRequest_bits_data_hi_125, memRequest_bits_data_lo_125};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_124, memRequest_bits_data_lo_124};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_129, memRequest_bits_data_lo_129, memRequest_bits_data_hi_128, memRequest_bits_data_lo_128};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_127, memRequest_bits_data_lo_127};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_132, memRequest_bits_data_lo_132, memRequest_bits_data_hi_131, memRequest_bits_data_lo_131};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_130, memRequest_bits_data_lo_130};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_135, memRequest_bits_data_lo_135, memRequest_bits_data_hi_134, memRequest_bits_data_lo_134};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_133, memRequest_bits_data_lo_133};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_138, memRequest_bits_data_lo_138, memRequest_bits_data_hi_137, memRequest_bits_data_lo_137};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_136, memRequest_bits_data_lo_136};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_141, memRequest_bits_data_lo_141, memRequest_bits_data_hi_140, memRequest_bits_data_lo_140};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_139, memRequest_bits_data_lo_139};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_144, memRequest_bits_data_lo_144, memRequest_bits_data_hi_143, memRequest_bits_data_lo_143};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_142, memRequest_bits_data_lo_142};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_147, memRequest_bits_data_lo_147, memRequest_bits_data_hi_146, memRequest_bits_data_lo_146};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_145, memRequest_bits_data_lo_145};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_150, memRequest_bits_data_lo_150, memRequest_bits_data_hi_149, memRequest_bits_data_lo_149};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_148, memRequest_bits_data_lo_148};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_8};
  wire [383:0]     memRequest_bits_data_hi_lo_199 = {memRequest_bits_data_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_153, memRequest_bits_data_lo_153, memRequest_bits_data_hi_152, memRequest_bits_data_lo_152};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_151, memRequest_bits_data_lo_151};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_156, memRequest_bits_data_lo_156, memRequest_bits_data_hi_155, memRequest_bits_data_lo_155};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_154, memRequest_bits_data_lo_154};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_159, memRequest_bits_data_lo_159, memRequest_bits_data_hi_158, memRequest_bits_data_lo_158};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_157, memRequest_bits_data_lo_157};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_162, memRequest_bits_data_lo_162, memRequest_bits_data_hi_161, memRequest_bits_data_lo_161};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_160, memRequest_bits_data_lo_160};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_165, memRequest_bits_data_lo_165, memRequest_bits_data_hi_164, memRequest_bits_data_lo_164};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_163, memRequest_bits_data_lo_163};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_168, memRequest_bits_data_lo_168, memRequest_bits_data_hi_167, memRequest_bits_data_lo_167};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_166, memRequest_bits_data_lo_166};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_171, memRequest_bits_data_lo_171, memRequest_bits_data_hi_170, memRequest_bits_data_lo_170};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_169, memRequest_bits_data_lo_169};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_174, memRequest_bits_data_lo_174, memRequest_bits_data_hi_173, memRequest_bits_data_lo_173};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_172, memRequest_bits_data_lo_172};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_177, memRequest_bits_data_lo_177, memRequest_bits_data_hi_176, memRequest_bits_data_lo_176};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_175, memRequest_bits_data_lo_175};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_180, memRequest_bits_data_lo_180, memRequest_bits_data_hi_179, memRequest_bits_data_lo_179};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_178, memRequest_bits_data_lo_178};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_183, memRequest_bits_data_lo_183, memRequest_bits_data_hi_182, memRequest_bits_data_lo_182};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_181, memRequest_bits_data_lo_181};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_186, memRequest_bits_data_lo_186, memRequest_bits_data_hi_185, memRequest_bits_data_lo_185};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_184, memRequest_bits_data_lo_184};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_189, memRequest_bits_data_lo_189, memRequest_bits_data_hi_188, memRequest_bits_data_lo_188};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_187, memRequest_bits_data_lo_187};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_192, memRequest_bits_data_lo_192, memRequest_bits_data_hi_191, memRequest_bits_data_lo_191};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_190, memRequest_bits_data_lo_190};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_195, memRequest_bits_data_lo_195, memRequest_bits_data_hi_194, memRequest_bits_data_lo_194};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_193, memRequest_bits_data_lo_193};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_198, memRequest_bits_data_lo_198, memRequest_bits_data_hi_197, memRequest_bits_data_lo_197};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_196, memRequest_bits_data_lo_196};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_8};
  wire [383:0]     memRequest_bits_data_hi_hi_199 = {memRequest_bits_data_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_8};
  wire [767:0]     memRequest_bits_data_hi_199 = {memRequest_bits_data_hi_hi_199, memRequest_bits_data_hi_lo_199};
  wire [511:0]     memRequest_bits_data_0 = {memRequest_bits_data_hi_199[263:0], memRequest_bits_data_lo_199[759:512]};
  wire [63:0]      selectMaskForTail = bufferValid ? _GEN_568 : 64'h0;
  wire [190:0]     _memRequest_bits_mask_T_1 = {63'h0, selectMaskForTail, maskTemp} << _GEN_569;
  wire [63:0]      memRequest_bits_mask_0 = _memRequest_bits_mask_T_1[127:64];
  assign alignedDequeueAddress = {lsuRequestReg_rs1Data[31:6] + {20'h0, bufferBaseCacheLineIndex}, 6'h0};
  wire [31:0]      memRequest_bits_address_0 = alignedDequeueAddress;
  wire [31:0]      addressQueue_enq_bits = alignedDequeueAddress;
  assign addressQueueFree = addressQueue_enq_ready;
  wire             addressQueue_deq_valid;
  assign addressQueue_deq_valid = ~_addressQueue_fifo_empty;
  assign addressQueue_enq_ready = ~_addressQueue_fifo_full;
  wire             _status_idle_output = ~bufferValid & ~readStageValid & readQueueClear & ~bufferFull & ~addressQueue_deq_valid;
  reg              idleNext;
  wire [31:0]      addressQueue_deq_bits;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 12'h0;
      csrInterfaceReg_vStart <= 12'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 64'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 63'h0;
      maskGroupCounter <= 5'h0;
      maskCounterInGroup <= 2'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 512'h0;
      accessData_1 <= 512'h0;
      accessData_2 <= 512'h0;
      accessData_3 <= 512'h0;
      accessData_4 <= 512'h0;
      accessData_5 <= 512'h0;
      accessData_6 <= 512'h0;
      accessData_7 <= 512'h0;
      accessPtr <= 3'h0;
      dataGroup <= 5'h0;
      dataBuffer_0 <= 512'h0;
      dataBuffer_1 <= 512'h0;
      dataBuffer_2 <= 512'h0;
      dataBuffer_3 <= 512'h0;
      dataBuffer_4 <= 512'h0;
      dataBuffer_5 <= 512'h0;
      dataBuffer_6 <= 512'h0;
      dataBuffer_7 <= 512'h0;
      bufferBaseCacheLineIndex <= 6'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 13'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 13'h0;
      lastDataGroupReg <= 9'h0;
      hazardCheck <= 1'h0;
      readStageValid_segPtr <= 3'h0;
      readStageValid_readCount <= 5'h0;
      readStageValid_stageValid <= 1'h0;
      readStageValid_readCounter <= 4'h0;
      readStageValid_segPtr_1 <= 3'h0;
      readStageValid_readCount_1 <= 5'h0;
      readStageValid_stageValid_1 <= 1'h0;
      readStageValid_readCounter_1 <= 4'h0;
      readStageValid_segPtr_2 <= 3'h0;
      readStageValid_readCount_2 <= 5'h0;
      readStageValid_stageValid_2 <= 1'h0;
      readStageValid_readCounter_2 <= 4'h0;
      readStageValid_segPtr_3 <= 3'h0;
      readStageValid_readCount_3 <= 5'h0;
      readStageValid_stageValid_3 <= 1'h0;
      readStageValid_readCounter_3 <= 4'h0;
      readStageValid_segPtr_4 <= 3'h0;
      readStageValid_readCount_4 <= 5'h0;
      readStageValid_stageValid_4 <= 1'h0;
      readStageValid_readCounter_4 <= 4'h0;
      readStageValid_segPtr_5 <= 3'h0;
      readStageValid_readCount_5 <= 5'h0;
      readStageValid_stageValid_5 <= 1'h0;
      readStageValid_readCounter_5 <= 4'h0;
      readStageValid_segPtr_6 <= 3'h0;
      readStageValid_readCount_6 <= 5'h0;
      readStageValid_stageValid_6 <= 1'h0;
      readStageValid_readCounter_6 <= 4'h0;
      readStageValid_segPtr_7 <= 3'h0;
      readStageValid_readCount_7 <= 5'h0;
      readStageValid_stageValid_7 <= 1'h0;
      readStageValid_readCounter_7 <= 4'h0;
      readStageValid_segPtr_8 <= 3'h0;
      readStageValid_readCount_8 <= 5'h0;
      readStageValid_stageValid_8 <= 1'h0;
      readStageValid_readCounter_8 <= 4'h0;
      readStageValid_segPtr_9 <= 3'h0;
      readStageValid_readCount_9 <= 5'h0;
      readStageValid_stageValid_9 <= 1'h0;
      readStageValid_readCounter_9 <= 4'h0;
      readStageValid_segPtr_10 <= 3'h0;
      readStageValid_readCount_10 <= 5'h0;
      readStageValid_stageValid_10 <= 1'h0;
      readStageValid_readCounter_10 <= 4'h0;
      readStageValid_segPtr_11 <= 3'h0;
      readStageValid_readCount_11 <= 5'h0;
      readStageValid_stageValid_11 <= 1'h0;
      readStageValid_readCounter_11 <= 4'h0;
      readStageValid_segPtr_12 <= 3'h0;
      readStageValid_readCount_12 <= 5'h0;
      readStageValid_stageValid_12 <= 1'h0;
      readStageValid_readCounter_12 <= 4'h0;
      readStageValid_segPtr_13 <= 3'h0;
      readStageValid_readCount_13 <= 5'h0;
      readStageValid_stageValid_13 <= 1'h0;
      readStageValid_readCounter_13 <= 4'h0;
      readStageValid_segPtr_14 <= 3'h0;
      readStageValid_readCount_14 <= 5'h0;
      readStageValid_stageValid_14 <= 1'h0;
      readStageValid_readCounter_14 <= 4'h0;
      readStageValid_segPtr_15 <= 3'h0;
      readStageValid_readCount_15 <= 5'h0;
      readStageValid_stageValid_15 <= 1'h0;
      readStageValid_readCounter_15 <= 4'h0;
      bufferFull <= 1'h0;
      bufferValid <= 1'h0;
      maskForBufferData_0 <= 64'h0;
      maskForBufferData_1 <= 64'h0;
      maskForBufferData_2 <= 64'h0;
      maskForBufferData_3 <= 64'h0;
      maskForBufferData_4 <= 64'h0;
      maskForBufferData_5 <= 64'h0;
      maskForBufferData_6 <= 64'h0;
      maskForBufferData_7 <= 64'h0;
      lastDataGroupInDataBuffer <= 1'h0;
      cacheLineTemp <= 512'h0;
      maskTemp <= 64'h0;
      canSendTail <= 1'h0;
      idleNext <= 1'h1;
    end
    else begin
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[5:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
        lastDataGroupReg <= lastDataGroupForInstruction;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[11:6] == 6'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[11:6];
      end
      if (_GEN_565 & (_GEN_566 | lsuRequest_valid))
        maskGroupCounter <= _maskSelect_bits_output;
      if (_GEN_565) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        dataGroup <= nextDataGroup;
      end
      if (accessBufferDequeueFire | accessBufferEnqueueFire | requestFireNext) begin
        accessData_0 <= accessDataUpdate_0;
        accessData_1 <= accessDataUpdate_1;
        accessData_2 <= accessDataUpdate_2;
        accessData_3 <= accessDataUpdate_3;
        accessData_4 <= accessDataUpdate_4;
        accessData_5 <= accessDataUpdate_5;
        accessData_6 <= accessDataUpdate_6;
        accessData_7 <= accessDataUpdate_7;
        accessPtr <= accessBufferDequeueFire | lastPtr | requestFireNext ? lsuRequestReg_instructionInformation_nf - {2'h0, accessBufferEnqueueFire & ~lastPtr} : accessPtr - 3'h1;
      end
      if (accessBufferDequeueFire) begin
        automatic logic [4095:0] _GEN_570 =
          (dataEEWOH[0]
             ? (_fillBySeg_T[0] ? regroupLoadData_0_0 : 4096'h0) | (_fillBySeg_T[1] ? regroupLoadData_0_1 : 4096'h0) | (_fillBySeg_T[2] ? regroupLoadData_0_2 : 4096'h0) | (_fillBySeg_T[3] ? regroupLoadData_0_3 : 4096'h0)
               | (_fillBySeg_T[4] ? regroupLoadData_0_4 : 4096'h0) | (_fillBySeg_T[5] ? regroupLoadData_0_5 : 4096'h0) | (_fillBySeg_T[6] ? regroupLoadData_0_6 : 4096'h0) | (_fillBySeg_T[7] ? regroupLoadData_0_7 : 4096'h0)
             : 4096'h0)
          | (dataEEWOH[1]
               ? (_fillBySeg_T[0] ? regroupLoadData_1_0 : 4096'h0) | (_fillBySeg_T[1] ? regroupLoadData_1_1 : 4096'h0) | (_fillBySeg_T[2] ? regroupLoadData_1_2 : 4096'h0) | (_fillBySeg_T[3] ? regroupLoadData_1_3 : 4096'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_1_4 : 4096'h0) | (_fillBySeg_T[5] ? regroupLoadData_1_5 : 4096'h0) | (_fillBySeg_T[6] ? regroupLoadData_1_6 : 4096'h0) | (_fillBySeg_T[7] ? regroupLoadData_1_7 : 4096'h0)
               : 4096'h0)
          | (dataEEWOH[2]
               ? (_fillBySeg_T[0] ? regroupLoadData_2_0 : 4096'h0) | (_fillBySeg_T[1] ? regroupLoadData_2_1 : 4096'h0) | (_fillBySeg_T[2] ? regroupLoadData_2_2 : 4096'h0) | (_fillBySeg_T[3] ? regroupLoadData_2_3 : 4096'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_2_4 : 4096'h0) | (_fillBySeg_T[5] ? regroupLoadData_2_5 : 4096'h0) | (_fillBySeg_T[6] ? regroupLoadData_2_6 : 4096'h0) | (_fillBySeg_T[7] ? regroupLoadData_2_7 : 4096'h0)
               : 4096'h0);
        dataBuffer_0 <= _GEN_570[511:0];
        dataBuffer_1 <= _GEN_570[1023:512];
        dataBuffer_2 <= _GEN_570[1535:1024];
        dataBuffer_3 <= _GEN_570[2047:1536];
        dataBuffer_4 <= _GEN_570[2559:2048];
        dataBuffer_5 <= _GEN_570[3071:2560];
        dataBuffer_6 <= _GEN_570[3583:3072];
        dataBuffer_7 <= _GEN_570[4095:3584];
        maskForBufferData_0 <= fillBySeg[63:0];
        maskForBufferData_1 <= fillBySeg[127:64];
        maskForBufferData_2 <= fillBySeg[191:128];
        maskForBufferData_3 <= fillBySeg[255:192];
        maskForBufferData_4 <= fillBySeg[319:256];
        maskForBufferData_5 <= fillBySeg[383:320];
        maskForBufferData_6 <= fillBySeg[447:384];
        maskForBufferData_7 <= fillBySeg[511:448];
        lastDataGroupInDataBuffer <= isLastRead;
      end
      else if (alignedDequeueFire) begin
        dataBuffer_0 <= dataBuffer_1;
        dataBuffer_1 <= dataBuffer_2;
        dataBuffer_2 <= dataBuffer_3;
        dataBuffer_3 <= dataBuffer_4;
        dataBuffer_4 <= dataBuffer_5;
        dataBuffer_5 <= dataBuffer_6;
        dataBuffer_6 <= dataBuffer_7;
        dataBuffer_7 <= 512'h0;
      end
      if (lsuRequest_valid | alignedDequeueFire) begin
        bufferBaseCacheLineIndex <= lsuRequest_valid ? 6'h0 : bufferBaseCacheLineIndex + 6'h1;
        maskTemp <= lsuRequest_valid ? 64'h0 : _GEN_568;
        canSendTail <= ~lsuRequest_valid & bufferValid & isLastCacheLineInBuffer & lastDataGroupInDataBuffer;
      end
      if (accessBufferDequeueFire | alignedDequeueFire)
        cacheLineIndexInBuffer <= accessBufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      hazardCheck <= ~lsuRequest_valid;
      if (lsuRequest_valid | _readStageValid_T_11)
        readStageValid_segPtr <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_11 & readStageValid_lastReadPtr)
        readStageValid_readCount <= readStageValid_nextReadCount;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup & readStageValid_lastReadPtr & _readStageValid_T_11)
        readStageValid_stageValid <= lsuRequest_valid;
      if (_readStageValid_T_11 ^ vrfReadQueueVec_0_deq_ready & vrfReadQueueVec_0_deq_valid)
        readStageValid_readCounter <= readStageValid_readCounter + readStageValid_counterChange;
      if (lsuRequest_valid | _readStageValid_T_30)
        readStageValid_segPtr_1 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_1 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_1 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_30 & readStageValid_lastReadPtr_1)
        readStageValid_readCount_1 <= readStageValid_nextReadCount_1;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_1 & readStageValid_lastReadPtr_1 & _readStageValid_T_30)
        readStageValid_stageValid_1 <= lsuRequest_valid;
      if (_readStageValid_T_30 ^ vrfReadQueueVec_1_deq_ready & vrfReadQueueVec_1_deq_valid)
        readStageValid_readCounter_1 <= readStageValid_readCounter_1 + readStageValid_counterChange_1;
      if (lsuRequest_valid | _readStageValid_T_49)
        readStageValid_segPtr_2 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_2 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_2 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_49 & readStageValid_lastReadPtr_2)
        readStageValid_readCount_2 <= readStageValid_nextReadCount_2;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_2 & readStageValid_lastReadPtr_2 & _readStageValid_T_49)
        readStageValid_stageValid_2 <= lsuRequest_valid;
      if (_readStageValid_T_49 ^ vrfReadQueueVec_2_deq_ready & vrfReadQueueVec_2_deq_valid)
        readStageValid_readCounter_2 <= readStageValid_readCounter_2 + readStageValid_counterChange_2;
      if (lsuRequest_valid | _readStageValid_T_68)
        readStageValid_segPtr_3 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_3 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_3 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_68 & readStageValid_lastReadPtr_3)
        readStageValid_readCount_3 <= readStageValid_nextReadCount_3;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_3 & readStageValid_lastReadPtr_3 & _readStageValid_T_68)
        readStageValid_stageValid_3 <= lsuRequest_valid;
      if (_readStageValid_T_68 ^ vrfReadQueueVec_3_deq_ready & vrfReadQueueVec_3_deq_valid)
        readStageValid_readCounter_3 <= readStageValid_readCounter_3 + readStageValid_counterChange_3;
      if (lsuRequest_valid | _readStageValid_T_87)
        readStageValid_segPtr_4 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_4 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_4 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_87 & readStageValid_lastReadPtr_4)
        readStageValid_readCount_4 <= readStageValid_nextReadCount_4;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_4 & readStageValid_lastReadPtr_4 & _readStageValid_T_87)
        readStageValid_stageValid_4 <= lsuRequest_valid;
      if (_readStageValid_T_87 ^ vrfReadQueueVec_4_deq_ready & vrfReadQueueVec_4_deq_valid)
        readStageValid_readCounter_4 <= readStageValid_readCounter_4 + readStageValid_counterChange_4;
      if (lsuRequest_valid | _readStageValid_T_106)
        readStageValid_segPtr_5 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_5 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_5 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_106 & readStageValid_lastReadPtr_5)
        readStageValid_readCount_5 <= readStageValid_nextReadCount_5;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_5 & readStageValid_lastReadPtr_5 & _readStageValid_T_106)
        readStageValid_stageValid_5 <= lsuRequest_valid;
      if (_readStageValid_T_106 ^ vrfReadQueueVec_5_deq_ready & vrfReadQueueVec_5_deq_valid)
        readStageValid_readCounter_5 <= readStageValid_readCounter_5 + readStageValid_counterChange_5;
      if (lsuRequest_valid | _readStageValid_T_125)
        readStageValid_segPtr_6 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_6 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_6 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_125 & readStageValid_lastReadPtr_6)
        readStageValid_readCount_6 <= readStageValid_nextReadCount_6;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_6 & readStageValid_lastReadPtr_6 & _readStageValid_T_125)
        readStageValid_stageValid_6 <= lsuRequest_valid;
      if (_readStageValid_T_125 ^ vrfReadQueueVec_6_deq_ready & vrfReadQueueVec_6_deq_valid)
        readStageValid_readCounter_6 <= readStageValid_readCounter_6 + readStageValid_counterChange_6;
      if (lsuRequest_valid | _readStageValid_T_144)
        readStageValid_segPtr_7 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_7 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_7 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_144 & readStageValid_lastReadPtr_7)
        readStageValid_readCount_7 <= readStageValid_nextReadCount_7;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_7 & readStageValid_lastReadPtr_7 & _readStageValid_T_144)
        readStageValid_stageValid_7 <= lsuRequest_valid;
      if (_readStageValid_T_144 ^ vrfReadQueueVec_7_deq_ready & vrfReadQueueVec_7_deq_valid)
        readStageValid_readCounter_7 <= readStageValid_readCounter_7 + readStageValid_counterChange_7;
      if (lsuRequest_valid | _readStageValid_T_163)
        readStageValid_segPtr_8 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_8 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_8 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_163 & readStageValid_lastReadPtr_8)
        readStageValid_readCount_8 <= readStageValid_nextReadCount_8;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_8 & readStageValid_lastReadPtr_8 & _readStageValid_T_163)
        readStageValid_stageValid_8 <= lsuRequest_valid;
      if (_readStageValid_T_163 ^ vrfReadQueueVec_8_deq_ready & vrfReadQueueVec_8_deq_valid)
        readStageValid_readCounter_8 <= readStageValid_readCounter_8 + readStageValid_counterChange_8;
      if (lsuRequest_valid | _readStageValid_T_182)
        readStageValid_segPtr_9 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_9 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_9 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_182 & readStageValid_lastReadPtr_9)
        readStageValid_readCount_9 <= readStageValid_nextReadCount_9;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_9 & readStageValid_lastReadPtr_9 & _readStageValid_T_182)
        readStageValid_stageValid_9 <= lsuRequest_valid;
      if (_readStageValid_T_182 ^ vrfReadQueueVec_9_deq_ready & vrfReadQueueVec_9_deq_valid)
        readStageValid_readCounter_9 <= readStageValid_readCounter_9 + readStageValid_counterChange_9;
      if (lsuRequest_valid | _readStageValid_T_201)
        readStageValid_segPtr_10 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_10 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_10 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_201 & readStageValid_lastReadPtr_10)
        readStageValid_readCount_10 <= readStageValid_nextReadCount_10;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_10 & readStageValid_lastReadPtr_10 & _readStageValid_T_201)
        readStageValid_stageValid_10 <= lsuRequest_valid;
      if (_readStageValid_T_201 ^ vrfReadQueueVec_10_deq_ready & vrfReadQueueVec_10_deq_valid)
        readStageValid_readCounter_10 <= readStageValid_readCounter_10 + readStageValid_counterChange_10;
      if (lsuRequest_valid | _readStageValid_T_220)
        readStageValid_segPtr_11 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_11 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_11 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_220 & readStageValid_lastReadPtr_11)
        readStageValid_readCount_11 <= readStageValid_nextReadCount_11;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_11 & readStageValid_lastReadPtr_11 & _readStageValid_T_220)
        readStageValid_stageValid_11 <= lsuRequest_valid;
      if (_readStageValid_T_220 ^ vrfReadQueueVec_11_deq_ready & vrfReadQueueVec_11_deq_valid)
        readStageValid_readCounter_11 <= readStageValid_readCounter_11 + readStageValid_counterChange_11;
      if (lsuRequest_valid | _readStageValid_T_239)
        readStageValid_segPtr_12 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_12 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_12 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_239 & readStageValid_lastReadPtr_12)
        readStageValid_readCount_12 <= readStageValid_nextReadCount_12;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_12 & readStageValid_lastReadPtr_12 & _readStageValid_T_239)
        readStageValid_stageValid_12 <= lsuRequest_valid;
      if (_readStageValid_T_239 ^ vrfReadQueueVec_12_deq_ready & vrfReadQueueVec_12_deq_valid)
        readStageValid_readCounter_12 <= readStageValid_readCounter_12 + readStageValid_counterChange_12;
      if (lsuRequest_valid | _readStageValid_T_258)
        readStageValid_segPtr_13 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_13 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_13 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_258 & readStageValid_lastReadPtr_13)
        readStageValid_readCount_13 <= readStageValid_nextReadCount_13;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_13 & readStageValid_lastReadPtr_13 & _readStageValid_T_258)
        readStageValid_stageValid_13 <= lsuRequest_valid;
      if (_readStageValid_T_258 ^ vrfReadQueueVec_13_deq_ready & vrfReadQueueVec_13_deq_valid)
        readStageValid_readCounter_13 <= readStageValid_readCounter_13 + readStageValid_counterChange_13;
      if (lsuRequest_valid | _readStageValid_T_277)
        readStageValid_segPtr_14 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_14 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_14 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_277 & readStageValid_lastReadPtr_14)
        readStageValid_readCount_14 <= readStageValid_nextReadCount_14;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_14 & readStageValid_lastReadPtr_14 & _readStageValid_T_277)
        readStageValid_stageValid_14 <= lsuRequest_valid;
      if (_readStageValid_T_277 ^ vrfReadQueueVec_14_deq_ready & vrfReadQueueVec_14_deq_valid)
        readStageValid_readCounter_14 <= readStageValid_readCounter_14 + readStageValid_counterChange_14;
      if (lsuRequest_valid | _readStageValid_T_296)
        readStageValid_segPtr_15 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_15 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_15 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_296 & readStageValid_lastReadPtr_15)
        readStageValid_readCount_15 <= readStageValid_nextReadCount_15;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_15 & readStageValid_lastReadPtr_15 & _readStageValid_T_296)
        readStageValid_stageValid_15 <= lsuRequest_valid;
      if (_readStageValid_T_296 ^ vrfReadQueueVec_15_deq_ready & vrfReadQueueVec_15_deq_valid)
        readStageValid_readCounter_15 <= readStageValid_readCounter_15 + readStageValid_counterChange_15;
      if (lastPtrEnq ^ accessBufferDequeueFire)
        bufferFull <= lastPtrEnq;
      if (accessBufferDequeueFire ^ bufferWillClear)
        bufferValid <= accessBufferDequeueFire;
      if (alignedDequeueFire)
        cacheLineTemp <= dataBuffer_0;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:309];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h136; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[9'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[9'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[9'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[9'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[9'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[9'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[9'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[9'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[9'h0][31:20], _RANDOM[9'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[9'h1][31:20], _RANDOM[9'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[9'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[9'h2][31:23], _RANDOM[9'h3][2:0]};
        csrInterfaceReg_vStart = _RANDOM[9'h3][14:3];
        csrInterfaceReg_vlmul = _RANDOM[9'h3][17:15];
        csrInterfaceReg_vSew = _RANDOM[9'h3][19:18];
        csrInterfaceReg_vxrm = _RANDOM[9'h3][21:20];
        csrInterfaceReg_vta = _RANDOM[9'h3][22];
        csrInterfaceReg_vma = _RANDOM[9'h3][23];
        requestFireNext = _RANDOM[9'h3][24];
        dataEEW = _RANDOM[9'h3][26:25];
        maskReg = {_RANDOM[9'h3][31:27], _RANDOM[9'h4], _RANDOM[9'h5][26:0]};
        needAmend = _RANDOM[9'h5][27];
        lastMaskAmendReg = {_RANDOM[9'h5][31:28], _RANDOM[9'h6], _RANDOM[9'h7][26:0]};
        maskGroupCounter = _RANDOM[9'h7][31:27];
        maskCounterInGroup = _RANDOM[9'h8][1:0];
        isLastMaskGroup = _RANDOM[9'hA][2];
        accessData_0 =
          {_RANDOM[9'hA][31:3],
           _RANDOM[9'hB],
           _RANDOM[9'hC],
           _RANDOM[9'hD],
           _RANDOM[9'hE],
           _RANDOM[9'hF],
           _RANDOM[9'h10],
           _RANDOM[9'h11],
           _RANDOM[9'h12],
           _RANDOM[9'h13],
           _RANDOM[9'h14],
           _RANDOM[9'h15],
           _RANDOM[9'h16],
           _RANDOM[9'h17],
           _RANDOM[9'h18],
           _RANDOM[9'h19],
           _RANDOM[9'h1A][2:0]};
        accessData_1 =
          {_RANDOM[9'h1A][31:3],
           _RANDOM[9'h1B],
           _RANDOM[9'h1C],
           _RANDOM[9'h1D],
           _RANDOM[9'h1E],
           _RANDOM[9'h1F],
           _RANDOM[9'h20],
           _RANDOM[9'h21],
           _RANDOM[9'h22],
           _RANDOM[9'h23],
           _RANDOM[9'h24],
           _RANDOM[9'h25],
           _RANDOM[9'h26],
           _RANDOM[9'h27],
           _RANDOM[9'h28],
           _RANDOM[9'h29],
           _RANDOM[9'h2A][2:0]};
        accessData_2 =
          {_RANDOM[9'h2A][31:3],
           _RANDOM[9'h2B],
           _RANDOM[9'h2C],
           _RANDOM[9'h2D],
           _RANDOM[9'h2E],
           _RANDOM[9'h2F],
           _RANDOM[9'h30],
           _RANDOM[9'h31],
           _RANDOM[9'h32],
           _RANDOM[9'h33],
           _RANDOM[9'h34],
           _RANDOM[9'h35],
           _RANDOM[9'h36],
           _RANDOM[9'h37],
           _RANDOM[9'h38],
           _RANDOM[9'h39],
           _RANDOM[9'h3A][2:0]};
        accessData_3 =
          {_RANDOM[9'h3A][31:3],
           _RANDOM[9'h3B],
           _RANDOM[9'h3C],
           _RANDOM[9'h3D],
           _RANDOM[9'h3E],
           _RANDOM[9'h3F],
           _RANDOM[9'h40],
           _RANDOM[9'h41],
           _RANDOM[9'h42],
           _RANDOM[9'h43],
           _RANDOM[9'h44],
           _RANDOM[9'h45],
           _RANDOM[9'h46],
           _RANDOM[9'h47],
           _RANDOM[9'h48],
           _RANDOM[9'h49],
           _RANDOM[9'h4A][2:0]};
        accessData_4 =
          {_RANDOM[9'h4A][31:3],
           _RANDOM[9'h4B],
           _RANDOM[9'h4C],
           _RANDOM[9'h4D],
           _RANDOM[9'h4E],
           _RANDOM[9'h4F],
           _RANDOM[9'h50],
           _RANDOM[9'h51],
           _RANDOM[9'h52],
           _RANDOM[9'h53],
           _RANDOM[9'h54],
           _RANDOM[9'h55],
           _RANDOM[9'h56],
           _RANDOM[9'h57],
           _RANDOM[9'h58],
           _RANDOM[9'h59],
           _RANDOM[9'h5A][2:0]};
        accessData_5 =
          {_RANDOM[9'h5A][31:3],
           _RANDOM[9'h5B],
           _RANDOM[9'h5C],
           _RANDOM[9'h5D],
           _RANDOM[9'h5E],
           _RANDOM[9'h5F],
           _RANDOM[9'h60],
           _RANDOM[9'h61],
           _RANDOM[9'h62],
           _RANDOM[9'h63],
           _RANDOM[9'h64],
           _RANDOM[9'h65],
           _RANDOM[9'h66],
           _RANDOM[9'h67],
           _RANDOM[9'h68],
           _RANDOM[9'h69],
           _RANDOM[9'h6A][2:0]};
        accessData_6 =
          {_RANDOM[9'h6A][31:3],
           _RANDOM[9'h6B],
           _RANDOM[9'h6C],
           _RANDOM[9'h6D],
           _RANDOM[9'h6E],
           _RANDOM[9'h6F],
           _RANDOM[9'h70],
           _RANDOM[9'h71],
           _RANDOM[9'h72],
           _RANDOM[9'h73],
           _RANDOM[9'h74],
           _RANDOM[9'h75],
           _RANDOM[9'h76],
           _RANDOM[9'h77],
           _RANDOM[9'h78],
           _RANDOM[9'h79],
           _RANDOM[9'h7A][2:0]};
        accessData_7 =
          {_RANDOM[9'h7A][31:3],
           _RANDOM[9'h7B],
           _RANDOM[9'h7C],
           _RANDOM[9'h7D],
           _RANDOM[9'h7E],
           _RANDOM[9'h7F],
           _RANDOM[9'h80],
           _RANDOM[9'h81],
           _RANDOM[9'h82],
           _RANDOM[9'h83],
           _RANDOM[9'h84],
           _RANDOM[9'h85],
           _RANDOM[9'h86],
           _RANDOM[9'h87],
           _RANDOM[9'h88],
           _RANDOM[9'h89],
           _RANDOM[9'h8A][2:0]};
        accessPtr = _RANDOM[9'h8A][5:3];
        dataGroup = _RANDOM[9'h8A][26:22];
        dataBuffer_0 =
          {_RANDOM[9'h8A][31:27],
           _RANDOM[9'h8B],
           _RANDOM[9'h8C],
           _RANDOM[9'h8D],
           _RANDOM[9'h8E],
           _RANDOM[9'h8F],
           _RANDOM[9'h90],
           _RANDOM[9'h91],
           _RANDOM[9'h92],
           _RANDOM[9'h93],
           _RANDOM[9'h94],
           _RANDOM[9'h95],
           _RANDOM[9'h96],
           _RANDOM[9'h97],
           _RANDOM[9'h98],
           _RANDOM[9'h99],
           _RANDOM[9'h9A][26:0]};
        dataBuffer_1 =
          {_RANDOM[9'h9A][31:27],
           _RANDOM[9'h9B],
           _RANDOM[9'h9C],
           _RANDOM[9'h9D],
           _RANDOM[9'h9E],
           _RANDOM[9'h9F],
           _RANDOM[9'hA0],
           _RANDOM[9'hA1],
           _RANDOM[9'hA2],
           _RANDOM[9'hA3],
           _RANDOM[9'hA4],
           _RANDOM[9'hA5],
           _RANDOM[9'hA6],
           _RANDOM[9'hA7],
           _RANDOM[9'hA8],
           _RANDOM[9'hA9],
           _RANDOM[9'hAA][26:0]};
        dataBuffer_2 =
          {_RANDOM[9'hAA][31:27],
           _RANDOM[9'hAB],
           _RANDOM[9'hAC],
           _RANDOM[9'hAD],
           _RANDOM[9'hAE],
           _RANDOM[9'hAF],
           _RANDOM[9'hB0],
           _RANDOM[9'hB1],
           _RANDOM[9'hB2],
           _RANDOM[9'hB3],
           _RANDOM[9'hB4],
           _RANDOM[9'hB5],
           _RANDOM[9'hB6],
           _RANDOM[9'hB7],
           _RANDOM[9'hB8],
           _RANDOM[9'hB9],
           _RANDOM[9'hBA][26:0]};
        dataBuffer_3 =
          {_RANDOM[9'hBA][31:27],
           _RANDOM[9'hBB],
           _RANDOM[9'hBC],
           _RANDOM[9'hBD],
           _RANDOM[9'hBE],
           _RANDOM[9'hBF],
           _RANDOM[9'hC0],
           _RANDOM[9'hC1],
           _RANDOM[9'hC2],
           _RANDOM[9'hC3],
           _RANDOM[9'hC4],
           _RANDOM[9'hC5],
           _RANDOM[9'hC6],
           _RANDOM[9'hC7],
           _RANDOM[9'hC8],
           _RANDOM[9'hC9],
           _RANDOM[9'hCA][26:0]};
        dataBuffer_4 =
          {_RANDOM[9'hCA][31:27],
           _RANDOM[9'hCB],
           _RANDOM[9'hCC],
           _RANDOM[9'hCD],
           _RANDOM[9'hCE],
           _RANDOM[9'hCF],
           _RANDOM[9'hD0],
           _RANDOM[9'hD1],
           _RANDOM[9'hD2],
           _RANDOM[9'hD3],
           _RANDOM[9'hD4],
           _RANDOM[9'hD5],
           _RANDOM[9'hD6],
           _RANDOM[9'hD7],
           _RANDOM[9'hD8],
           _RANDOM[9'hD9],
           _RANDOM[9'hDA][26:0]};
        dataBuffer_5 =
          {_RANDOM[9'hDA][31:27],
           _RANDOM[9'hDB],
           _RANDOM[9'hDC],
           _RANDOM[9'hDD],
           _RANDOM[9'hDE],
           _RANDOM[9'hDF],
           _RANDOM[9'hE0],
           _RANDOM[9'hE1],
           _RANDOM[9'hE2],
           _RANDOM[9'hE3],
           _RANDOM[9'hE4],
           _RANDOM[9'hE5],
           _RANDOM[9'hE6],
           _RANDOM[9'hE7],
           _RANDOM[9'hE8],
           _RANDOM[9'hE9],
           _RANDOM[9'hEA][26:0]};
        dataBuffer_6 =
          {_RANDOM[9'hEA][31:27],
           _RANDOM[9'hEB],
           _RANDOM[9'hEC],
           _RANDOM[9'hED],
           _RANDOM[9'hEE],
           _RANDOM[9'hEF],
           _RANDOM[9'hF0],
           _RANDOM[9'hF1],
           _RANDOM[9'hF2],
           _RANDOM[9'hF3],
           _RANDOM[9'hF4],
           _RANDOM[9'hF5],
           _RANDOM[9'hF6],
           _RANDOM[9'hF7],
           _RANDOM[9'hF8],
           _RANDOM[9'hF9],
           _RANDOM[9'hFA][26:0]};
        dataBuffer_7 =
          {_RANDOM[9'hFA][31:27],
           _RANDOM[9'hFB],
           _RANDOM[9'hFC],
           _RANDOM[9'hFD],
           _RANDOM[9'hFE],
           _RANDOM[9'hFF],
           _RANDOM[9'h100],
           _RANDOM[9'h101],
           _RANDOM[9'h102],
           _RANDOM[9'h103],
           _RANDOM[9'h104],
           _RANDOM[9'h105],
           _RANDOM[9'h106],
           _RANDOM[9'h107],
           _RANDOM[9'h108],
           _RANDOM[9'h109],
           _RANDOM[9'h10A][26:0]};
        bufferBaseCacheLineIndex = {_RANDOM[9'h10A][31:27], _RANDOM[9'h10B][0]};
        cacheLineIndexInBuffer = _RANDOM[9'h10B][3:1];
        invalidInstructionNext = _RANDOM[9'h10B][4];
        segmentInstructionIndexInterval = _RANDOM[9'h10B][8:5];
        lastWriteVrfIndexReg = _RANDOM[9'h10B][21:9];
        lastCacheNeedPush = _RANDOM[9'h10B][22];
        cacheLineNumberReg = {_RANDOM[9'h10B][31:23], _RANDOM[9'h10C][3:0]};
        lastDataGroupReg = _RANDOM[9'h10C][12:4];
        hazardCheck = _RANDOM[9'h10C][13];
        readStageValid_segPtr = _RANDOM[9'h10C][16:14];
        readStageValid_readCount = _RANDOM[9'h10C][21:17];
        readStageValid_stageValid = _RANDOM[9'h10C][22];
        readStageValid_readCounter = _RANDOM[9'h10C][26:23];
        readStageValid_segPtr_1 = _RANDOM[9'h10C][29:27];
        readStageValid_readCount_1 = {_RANDOM[9'h10C][31:30], _RANDOM[9'h10D][2:0]};
        readStageValid_stageValid_1 = _RANDOM[9'h10D][3];
        readStageValid_readCounter_1 = _RANDOM[9'h10D][7:4];
        readStageValid_segPtr_2 = _RANDOM[9'h10D][10:8];
        readStageValid_readCount_2 = _RANDOM[9'h10D][15:11];
        readStageValid_stageValid_2 = _RANDOM[9'h10D][16];
        readStageValid_readCounter_2 = _RANDOM[9'h10D][20:17];
        readStageValid_segPtr_3 = _RANDOM[9'h10D][23:21];
        readStageValid_readCount_3 = _RANDOM[9'h10D][28:24];
        readStageValid_stageValid_3 = _RANDOM[9'h10D][29];
        readStageValid_readCounter_3 = {_RANDOM[9'h10D][31:30], _RANDOM[9'h10E][1:0]};
        readStageValid_segPtr_4 = _RANDOM[9'h10E][4:2];
        readStageValid_readCount_4 = _RANDOM[9'h10E][9:5];
        readStageValid_stageValid_4 = _RANDOM[9'h10E][10];
        readStageValid_readCounter_4 = _RANDOM[9'h10E][14:11];
        readStageValid_segPtr_5 = _RANDOM[9'h10E][17:15];
        readStageValid_readCount_5 = _RANDOM[9'h10E][22:18];
        readStageValid_stageValid_5 = _RANDOM[9'h10E][23];
        readStageValid_readCounter_5 = _RANDOM[9'h10E][27:24];
        readStageValid_segPtr_6 = _RANDOM[9'h10E][30:28];
        readStageValid_readCount_6 = {_RANDOM[9'h10E][31], _RANDOM[9'h10F][3:0]};
        readStageValid_stageValid_6 = _RANDOM[9'h10F][4];
        readStageValid_readCounter_6 = _RANDOM[9'h10F][8:5];
        readStageValid_segPtr_7 = _RANDOM[9'h10F][11:9];
        readStageValid_readCount_7 = _RANDOM[9'h10F][16:12];
        readStageValid_stageValid_7 = _RANDOM[9'h10F][17];
        readStageValid_readCounter_7 = _RANDOM[9'h10F][21:18];
        readStageValid_segPtr_8 = _RANDOM[9'h10F][24:22];
        readStageValid_readCount_8 = _RANDOM[9'h10F][29:25];
        readStageValid_stageValid_8 = _RANDOM[9'h10F][30];
        readStageValid_readCounter_8 = {_RANDOM[9'h10F][31], _RANDOM[9'h110][2:0]};
        readStageValid_segPtr_9 = _RANDOM[9'h110][5:3];
        readStageValid_readCount_9 = _RANDOM[9'h110][10:6];
        readStageValid_stageValid_9 = _RANDOM[9'h110][11];
        readStageValid_readCounter_9 = _RANDOM[9'h110][15:12];
        readStageValid_segPtr_10 = _RANDOM[9'h110][18:16];
        readStageValid_readCount_10 = _RANDOM[9'h110][23:19];
        readStageValid_stageValid_10 = _RANDOM[9'h110][24];
        readStageValid_readCounter_10 = _RANDOM[9'h110][28:25];
        readStageValid_segPtr_11 = _RANDOM[9'h110][31:29];
        readStageValid_readCount_11 = _RANDOM[9'h111][4:0];
        readStageValid_stageValid_11 = _RANDOM[9'h111][5];
        readStageValid_readCounter_11 = _RANDOM[9'h111][9:6];
        readStageValid_segPtr_12 = _RANDOM[9'h111][12:10];
        readStageValid_readCount_12 = _RANDOM[9'h111][17:13];
        readStageValid_stageValid_12 = _RANDOM[9'h111][18];
        readStageValid_readCounter_12 = _RANDOM[9'h111][22:19];
        readStageValid_segPtr_13 = _RANDOM[9'h111][25:23];
        readStageValid_readCount_13 = _RANDOM[9'h111][30:26];
        readStageValid_stageValid_13 = _RANDOM[9'h111][31];
        readStageValid_readCounter_13 = _RANDOM[9'h112][3:0];
        readStageValid_segPtr_14 = _RANDOM[9'h112][6:4];
        readStageValid_readCount_14 = _RANDOM[9'h112][11:7];
        readStageValid_stageValid_14 = _RANDOM[9'h112][12];
        readStageValid_readCounter_14 = _RANDOM[9'h112][16:13];
        readStageValid_segPtr_15 = _RANDOM[9'h112][19:17];
        readStageValid_readCount_15 = _RANDOM[9'h112][24:20];
        readStageValid_stageValid_15 = _RANDOM[9'h112][25];
        readStageValid_readCounter_15 = _RANDOM[9'h112][29:26];
        bufferFull = _RANDOM[9'h112][30];
        bufferValid = _RANDOM[9'h112][31];
        maskForBufferData_0 = {_RANDOM[9'h113], _RANDOM[9'h114]};
        maskForBufferData_1 = {_RANDOM[9'h115], _RANDOM[9'h116]};
        maskForBufferData_2 = {_RANDOM[9'h117], _RANDOM[9'h118]};
        maskForBufferData_3 = {_RANDOM[9'h119], _RANDOM[9'h11A]};
        maskForBufferData_4 = {_RANDOM[9'h11B], _RANDOM[9'h11C]};
        maskForBufferData_5 = {_RANDOM[9'h11D], _RANDOM[9'h11E]};
        maskForBufferData_6 = {_RANDOM[9'h11F], _RANDOM[9'h120]};
        maskForBufferData_7 = {_RANDOM[9'h121], _RANDOM[9'h122]};
        lastDataGroupInDataBuffer = _RANDOM[9'h123][0];
        cacheLineTemp =
          {_RANDOM[9'h123][31:1],
           _RANDOM[9'h124],
           _RANDOM[9'h125],
           _RANDOM[9'h126],
           _RANDOM[9'h127],
           _RANDOM[9'h128],
           _RANDOM[9'h129],
           _RANDOM[9'h12A],
           _RANDOM[9'h12B],
           _RANDOM[9'h12C],
           _RANDOM[9'h12D],
           _RANDOM[9'h12E],
           _RANDOM[9'h12F],
           _RANDOM[9'h130],
           _RANDOM[9'h131],
           _RANDOM[9'h132],
           _RANDOM[9'h133][0]};
        maskTemp = {_RANDOM[9'h133][31:1], _RANDOM[9'h134], _RANDOM[9'h135][0]};
        canSendTail = _RANDOM[9'h135][1];
        idleNext = _RANDOM[9'h135][2];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire             vrfReadQueueVec_0_empty;
  assign vrfReadQueueVec_0_empty = _vrfReadQueueVec_fifo_empty;
  wire             vrfReadQueueVec_0_full;
  assign vrfReadQueueVec_0_full = _vrfReadQueueVec_fifo_full;
  wire             vrfReadQueueVec_1_empty;
  assign vrfReadQueueVec_1_empty = _vrfReadQueueVec_fifo_1_empty;
  wire             vrfReadQueueVec_1_full;
  assign vrfReadQueueVec_1_full = _vrfReadQueueVec_fifo_1_full;
  wire             vrfReadQueueVec_2_empty;
  assign vrfReadQueueVec_2_empty = _vrfReadQueueVec_fifo_2_empty;
  wire             vrfReadQueueVec_2_full;
  assign vrfReadQueueVec_2_full = _vrfReadQueueVec_fifo_2_full;
  wire             vrfReadQueueVec_3_empty;
  assign vrfReadQueueVec_3_empty = _vrfReadQueueVec_fifo_3_empty;
  wire             vrfReadQueueVec_3_full;
  assign vrfReadQueueVec_3_full = _vrfReadQueueVec_fifo_3_full;
  wire             vrfReadQueueVec_4_empty;
  assign vrfReadQueueVec_4_empty = _vrfReadQueueVec_fifo_4_empty;
  wire             vrfReadQueueVec_4_full;
  assign vrfReadQueueVec_4_full = _vrfReadQueueVec_fifo_4_full;
  wire             vrfReadQueueVec_5_empty;
  assign vrfReadQueueVec_5_empty = _vrfReadQueueVec_fifo_5_empty;
  wire             vrfReadQueueVec_5_full;
  assign vrfReadQueueVec_5_full = _vrfReadQueueVec_fifo_5_full;
  wire             vrfReadQueueVec_6_empty;
  assign vrfReadQueueVec_6_empty = _vrfReadQueueVec_fifo_6_empty;
  wire             vrfReadQueueVec_6_full;
  assign vrfReadQueueVec_6_full = _vrfReadQueueVec_fifo_6_full;
  wire             vrfReadQueueVec_7_empty;
  assign vrfReadQueueVec_7_empty = _vrfReadQueueVec_fifo_7_empty;
  wire             vrfReadQueueVec_7_full;
  assign vrfReadQueueVec_7_full = _vrfReadQueueVec_fifo_7_full;
  wire             vrfReadQueueVec_8_empty;
  assign vrfReadQueueVec_8_empty = _vrfReadQueueVec_fifo_8_empty;
  wire             vrfReadQueueVec_8_full;
  assign vrfReadQueueVec_8_full = _vrfReadQueueVec_fifo_8_full;
  wire             vrfReadQueueVec_9_empty;
  assign vrfReadQueueVec_9_empty = _vrfReadQueueVec_fifo_9_empty;
  wire             vrfReadQueueVec_9_full;
  assign vrfReadQueueVec_9_full = _vrfReadQueueVec_fifo_9_full;
  wire             vrfReadQueueVec_10_empty;
  assign vrfReadQueueVec_10_empty = _vrfReadQueueVec_fifo_10_empty;
  wire             vrfReadQueueVec_10_full;
  assign vrfReadQueueVec_10_full = _vrfReadQueueVec_fifo_10_full;
  wire             vrfReadQueueVec_11_empty;
  assign vrfReadQueueVec_11_empty = _vrfReadQueueVec_fifo_11_empty;
  wire             vrfReadQueueVec_11_full;
  assign vrfReadQueueVec_11_full = _vrfReadQueueVec_fifo_11_full;
  wire             vrfReadQueueVec_12_empty;
  assign vrfReadQueueVec_12_empty = _vrfReadQueueVec_fifo_12_empty;
  wire             vrfReadQueueVec_12_full;
  assign vrfReadQueueVec_12_full = _vrfReadQueueVec_fifo_12_full;
  wire             vrfReadQueueVec_13_empty;
  assign vrfReadQueueVec_13_empty = _vrfReadQueueVec_fifo_13_empty;
  wire             vrfReadQueueVec_13_full;
  assign vrfReadQueueVec_13_full = _vrfReadQueueVec_fifo_13_full;
  wire             vrfReadQueueVec_14_empty;
  assign vrfReadQueueVec_14_empty = _vrfReadQueueVec_fifo_14_empty;
  wire             vrfReadQueueVec_14_full;
  assign vrfReadQueueVec_14_full = _vrfReadQueueVec_fifo_14_full;
  wire             vrfReadQueueVec_15_empty;
  assign vrfReadQueueVec_15_empty = _vrfReadQueueVec_fifo_15_empty;
  wire             vrfReadQueueVec_15_full;
  assign vrfReadQueueVec_15_full = _vrfReadQueueVec_fifo_15_full;
  wire             addressQueue_empty;
  assign addressQueue_empty = _addressQueue_fifo_empty;
  wire             addressQueue_full;
  assign addressQueue_full = _addressQueue_fifo_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_0_enq_ready & vrfReadQueueVec_0_enq_valid & ~(_vrfReadQueueVec_fifo_empty & vrfReadQueueVec_0_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_0_deq_ready & ~_vrfReadQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_0_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_empty),
    .almost_empty (vrfReadQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_0_almostFull),
    .full         (_vrfReadQueueVec_fifo_full),
    .error        (_vrfReadQueueVec_fifo_error),
    .data_out     (_vrfReadQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_1_enq_ready & vrfReadQueueVec_1_enq_valid & ~(_vrfReadQueueVec_fifo_1_empty & vrfReadQueueVec_1_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_1_deq_ready & ~_vrfReadQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_1_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_1_empty),
    .almost_empty (vrfReadQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_1_almostFull),
    .full         (_vrfReadQueueVec_fifo_1_full),
    .error        (_vrfReadQueueVec_fifo_1_error),
    .data_out     (_vrfReadQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_2_enq_ready & vrfReadQueueVec_2_enq_valid & ~(_vrfReadQueueVec_fifo_2_empty & vrfReadQueueVec_2_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_2_deq_ready & ~_vrfReadQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_2_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_2_empty),
    .almost_empty (vrfReadQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_2_almostFull),
    .full         (_vrfReadQueueVec_fifo_2_full),
    .error        (_vrfReadQueueVec_fifo_2_error),
    .data_out     (_vrfReadQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_3_enq_ready & vrfReadQueueVec_3_enq_valid & ~(_vrfReadQueueVec_fifo_3_empty & vrfReadQueueVec_3_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_3_deq_ready & ~_vrfReadQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_3_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_3_empty),
    .almost_empty (vrfReadQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_3_almostFull),
    .full         (_vrfReadQueueVec_fifo_3_full),
    .error        (_vrfReadQueueVec_fifo_3_error),
    .data_out     (_vrfReadQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_4_enq_ready & vrfReadQueueVec_4_enq_valid & ~(_vrfReadQueueVec_fifo_4_empty & vrfReadQueueVec_4_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_4_deq_ready & ~_vrfReadQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_4_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_4_empty),
    .almost_empty (vrfReadQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_4_almostFull),
    .full         (_vrfReadQueueVec_fifo_4_full),
    .error        (_vrfReadQueueVec_fifo_4_error),
    .data_out     (_vrfReadQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_5_enq_ready & vrfReadQueueVec_5_enq_valid & ~(_vrfReadQueueVec_fifo_5_empty & vrfReadQueueVec_5_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_5_deq_ready & ~_vrfReadQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_5_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_5_empty),
    .almost_empty (vrfReadQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_5_almostFull),
    .full         (_vrfReadQueueVec_fifo_5_full),
    .error        (_vrfReadQueueVec_fifo_5_error),
    .data_out     (_vrfReadQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_6_enq_ready & vrfReadQueueVec_6_enq_valid & ~(_vrfReadQueueVec_fifo_6_empty & vrfReadQueueVec_6_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_6_deq_ready & ~_vrfReadQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_6_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_6_empty),
    .almost_empty (vrfReadQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_6_almostFull),
    .full         (_vrfReadQueueVec_fifo_6_full),
    .error        (_vrfReadQueueVec_fifo_6_error),
    .data_out     (_vrfReadQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_7_enq_ready & vrfReadQueueVec_7_enq_valid & ~(_vrfReadQueueVec_fifo_7_empty & vrfReadQueueVec_7_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_7_deq_ready & ~_vrfReadQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_7_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_7_empty),
    .almost_empty (vrfReadQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_7_almostFull),
    .full         (_vrfReadQueueVec_fifo_7_full),
    .error        (_vrfReadQueueVec_fifo_7_error),
    .data_out     (_vrfReadQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_8_enq_ready & vrfReadQueueVec_8_enq_valid & ~(_vrfReadQueueVec_fifo_8_empty & vrfReadQueueVec_8_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_8_deq_ready & ~_vrfReadQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_8_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_8_empty),
    .almost_empty (vrfReadQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_8_almostFull),
    .full         (_vrfReadQueueVec_fifo_8_full),
    .error        (_vrfReadQueueVec_fifo_8_error),
    .data_out     (_vrfReadQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_9_enq_ready & vrfReadQueueVec_9_enq_valid & ~(_vrfReadQueueVec_fifo_9_empty & vrfReadQueueVec_9_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_9_deq_ready & ~_vrfReadQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_9_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_9_empty),
    .almost_empty (vrfReadQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_9_almostFull),
    .full         (_vrfReadQueueVec_fifo_9_full),
    .error        (_vrfReadQueueVec_fifo_9_error),
    .data_out     (_vrfReadQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_10_enq_ready & vrfReadQueueVec_10_enq_valid & ~(_vrfReadQueueVec_fifo_10_empty & vrfReadQueueVec_10_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_10_deq_ready & ~_vrfReadQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_10_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_10_empty),
    .almost_empty (vrfReadQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_10_almostFull),
    .full         (_vrfReadQueueVec_fifo_10_full),
    .error        (_vrfReadQueueVec_fifo_10_error),
    .data_out     (_vrfReadQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_11_enq_ready & vrfReadQueueVec_11_enq_valid & ~(_vrfReadQueueVec_fifo_11_empty & vrfReadQueueVec_11_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_11_deq_ready & ~_vrfReadQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_11_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_11_empty),
    .almost_empty (vrfReadQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_11_almostFull),
    .full         (_vrfReadQueueVec_fifo_11_full),
    .error        (_vrfReadQueueVec_fifo_11_error),
    .data_out     (_vrfReadQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_12_enq_ready & vrfReadQueueVec_12_enq_valid & ~(_vrfReadQueueVec_fifo_12_empty & vrfReadQueueVec_12_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_12_deq_ready & ~_vrfReadQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_12_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_12_empty),
    .almost_empty (vrfReadQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_12_almostFull),
    .full         (_vrfReadQueueVec_fifo_12_full),
    .error        (_vrfReadQueueVec_fifo_12_error),
    .data_out     (_vrfReadQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_13_enq_ready & vrfReadQueueVec_13_enq_valid & ~(_vrfReadQueueVec_fifo_13_empty & vrfReadQueueVec_13_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_13_deq_ready & ~_vrfReadQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_13_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_13_empty),
    .almost_empty (vrfReadQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_13_almostFull),
    .full         (_vrfReadQueueVec_fifo_13_full),
    .error        (_vrfReadQueueVec_fifo_13_error),
    .data_out     (_vrfReadQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_14_enq_ready & vrfReadQueueVec_14_enq_valid & ~(_vrfReadQueueVec_fifo_14_empty & vrfReadQueueVec_14_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_14_deq_ready & ~_vrfReadQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_14_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_14_empty),
    .almost_empty (vrfReadQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_14_almostFull),
    .full         (_vrfReadQueueVec_fifo_14_full),
    .error        (_vrfReadQueueVec_fifo_14_error),
    .data_out     (_vrfReadQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_15_enq_ready & vrfReadQueueVec_15_enq_valid & ~(_vrfReadQueueVec_fifo_15_empty & vrfReadQueueVec_15_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_15_deq_ready & ~_vrfReadQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_15_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_15_empty),
    .almost_empty (vrfReadQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_15_almostFull),
    .full         (_vrfReadQueueVec_fifo_15_full),
    .error        (_vrfReadQueueVec_fifo_15_error),
    .data_out     (_vrfReadQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) addressQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(addressQueue_enq_ready & addressQueue_enq_valid)),
    .pop_req_n    (~(addressQueue_deq_ready & ~_addressQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (addressQueue_enq_bits),
    .empty        (_addressQueue_fifo_empty),
    .almost_empty (addressQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (addressQueue_almostFull),
    .full         (_addressQueue_fifo_full),
    .error        (_addressQueue_fifo_error),
    .data_out     (addressQueue_deq_bits)
  );
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_data = memRequest_bits_data_0;
  assign memRequest_bits_mask = memRequest_bits_mask_0;
  assign memRequest_bits_index = memRequest_bits_index_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = addressQueue_deq_valid ? addressQueue_deq_bits : alignedDequeueAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:6] + {13'h0, cacheLineNumberReg}, 6'h0};
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfReadDataPorts_4_valid = vrfReadDataPorts_4_valid_0;
  assign vrfReadDataPorts_4_bits_vs = vrfReadDataPorts_4_bits_vs_0;
  assign vrfReadDataPorts_4_bits_offset = vrfReadDataPorts_4_bits_offset_0;
  assign vrfReadDataPorts_4_bits_instructionIndex = vrfReadDataPorts_4_bits_instructionIndex_0;
  assign vrfReadDataPorts_5_valid = vrfReadDataPorts_5_valid_0;
  assign vrfReadDataPorts_5_bits_vs = vrfReadDataPorts_5_bits_vs_0;
  assign vrfReadDataPorts_5_bits_offset = vrfReadDataPorts_5_bits_offset_0;
  assign vrfReadDataPorts_5_bits_instructionIndex = vrfReadDataPorts_5_bits_instructionIndex_0;
  assign vrfReadDataPorts_6_valid = vrfReadDataPorts_6_valid_0;
  assign vrfReadDataPorts_6_bits_vs = vrfReadDataPorts_6_bits_vs_0;
  assign vrfReadDataPorts_6_bits_offset = vrfReadDataPorts_6_bits_offset_0;
  assign vrfReadDataPorts_6_bits_instructionIndex = vrfReadDataPorts_6_bits_instructionIndex_0;
  assign vrfReadDataPorts_7_valid = vrfReadDataPorts_7_valid_0;
  assign vrfReadDataPorts_7_bits_vs = vrfReadDataPorts_7_bits_vs_0;
  assign vrfReadDataPorts_7_bits_offset = vrfReadDataPorts_7_bits_offset_0;
  assign vrfReadDataPorts_7_bits_instructionIndex = vrfReadDataPorts_7_bits_instructionIndex_0;
  assign vrfReadDataPorts_8_valid = vrfReadDataPorts_8_valid_0;
  assign vrfReadDataPorts_8_bits_vs = vrfReadDataPorts_8_bits_vs_0;
  assign vrfReadDataPorts_8_bits_offset = vrfReadDataPorts_8_bits_offset_0;
  assign vrfReadDataPorts_8_bits_instructionIndex = vrfReadDataPorts_8_bits_instructionIndex_0;
  assign vrfReadDataPorts_9_valid = vrfReadDataPorts_9_valid_0;
  assign vrfReadDataPorts_9_bits_vs = vrfReadDataPorts_9_bits_vs_0;
  assign vrfReadDataPorts_9_bits_offset = vrfReadDataPorts_9_bits_offset_0;
  assign vrfReadDataPorts_9_bits_instructionIndex = vrfReadDataPorts_9_bits_instructionIndex_0;
  assign vrfReadDataPorts_10_valid = vrfReadDataPorts_10_valid_0;
  assign vrfReadDataPorts_10_bits_vs = vrfReadDataPorts_10_bits_vs_0;
  assign vrfReadDataPorts_10_bits_offset = vrfReadDataPorts_10_bits_offset_0;
  assign vrfReadDataPorts_10_bits_instructionIndex = vrfReadDataPorts_10_bits_instructionIndex_0;
  assign vrfReadDataPorts_11_valid = vrfReadDataPorts_11_valid_0;
  assign vrfReadDataPorts_11_bits_vs = vrfReadDataPorts_11_bits_vs_0;
  assign vrfReadDataPorts_11_bits_offset = vrfReadDataPorts_11_bits_offset_0;
  assign vrfReadDataPorts_11_bits_instructionIndex = vrfReadDataPorts_11_bits_instructionIndex_0;
  assign vrfReadDataPorts_12_valid = vrfReadDataPorts_12_valid_0;
  assign vrfReadDataPorts_12_bits_vs = vrfReadDataPorts_12_bits_vs_0;
  assign vrfReadDataPorts_12_bits_offset = vrfReadDataPorts_12_bits_offset_0;
  assign vrfReadDataPorts_12_bits_instructionIndex = vrfReadDataPorts_12_bits_instructionIndex_0;
  assign vrfReadDataPorts_13_valid = vrfReadDataPorts_13_valid_0;
  assign vrfReadDataPorts_13_bits_vs = vrfReadDataPorts_13_bits_vs_0;
  assign vrfReadDataPorts_13_bits_offset = vrfReadDataPorts_13_bits_offset_0;
  assign vrfReadDataPorts_13_bits_instructionIndex = vrfReadDataPorts_13_bits_instructionIndex_0;
  assign vrfReadDataPorts_14_valid = vrfReadDataPorts_14_valid_0;
  assign vrfReadDataPorts_14_bits_vs = vrfReadDataPorts_14_bits_vs_0;
  assign vrfReadDataPorts_14_bits_offset = vrfReadDataPorts_14_bits_offset_0;
  assign vrfReadDataPorts_14_bits_instructionIndex = vrfReadDataPorts_14_bits_instructionIndex_0;
  assign vrfReadDataPorts_15_valid = vrfReadDataPorts_15_valid_0;
  assign vrfReadDataPorts_15_bits_vs = vrfReadDataPorts_15_bits_vs_0;
  assign vrfReadDataPorts_15_bits_offset = vrfReadDataPorts_15_bits_offset_0;
  assign vrfReadDataPorts_15_bits_instructionIndex = vrfReadDataPorts_15_bits_instructionIndex_0;
endmodule

