module CarrySaveAdder_28(
  input  [27:0] in_0,
                in_1,
                in_2,
  output [27:0] out_0,
                out_1
);

  wire        out_xor01 = in_0[0] ^ in_1[0];
  wire        out_0_0 = in_0[0] & in_1[0] | out_xor01 & in_2[0];
  wire        out_1_0 = out_xor01 ^ in_2[0];
  wire        out_xor01_1 = in_0[1] ^ in_1[1];
  wire        out_0_1 = in_0[1] & in_1[1] | out_xor01_1 & in_2[1];
  wire        out_1_1 = out_xor01_1 ^ in_2[1];
  wire        out_xor01_2 = in_0[2] ^ in_1[2];
  wire        out_0_2 = in_0[2] & in_1[2] | out_xor01_2 & in_2[2];
  wire        out_1_2 = out_xor01_2 ^ in_2[2];
  wire        out_xor01_3 = in_0[3] ^ in_1[3];
  wire        out_0_3 = in_0[3] & in_1[3] | out_xor01_3 & in_2[3];
  wire        out_1_3 = out_xor01_3 ^ in_2[3];
  wire        out_xor01_4 = in_0[4] ^ in_1[4];
  wire        out_0_4 = in_0[4] & in_1[4] | out_xor01_4 & in_2[4];
  wire        out_1_4 = out_xor01_4 ^ in_2[4];
  wire        out_xor01_5 = in_0[5] ^ in_1[5];
  wire        out_0_5 = in_0[5] & in_1[5] | out_xor01_5 & in_2[5];
  wire        out_1_5 = out_xor01_5 ^ in_2[5];
  wire        out_xor01_6 = in_0[6] ^ in_1[6];
  wire        out_0_6 = in_0[6] & in_1[6] | out_xor01_6 & in_2[6];
  wire        out_1_6 = out_xor01_6 ^ in_2[6];
  wire        out_xor01_7 = in_0[7] ^ in_1[7];
  wire        out_0_7 = in_0[7] & in_1[7] | out_xor01_7 & in_2[7];
  wire        out_1_7 = out_xor01_7 ^ in_2[7];
  wire        out_xor01_8 = in_0[8] ^ in_1[8];
  wire        out_0_8 = in_0[8] & in_1[8] | out_xor01_8 & in_2[8];
  wire        out_1_8 = out_xor01_8 ^ in_2[8];
  wire        out_xor01_9 = in_0[9] ^ in_1[9];
  wire        out_0_9 = in_0[9] & in_1[9] | out_xor01_9 & in_2[9];
  wire        out_1_9 = out_xor01_9 ^ in_2[9];
  wire        out_xor01_10 = in_0[10] ^ in_1[10];
  wire        out_0_10 = in_0[10] & in_1[10] | out_xor01_10 & in_2[10];
  wire        out_1_10 = out_xor01_10 ^ in_2[10];
  wire        out_xor01_11 = in_0[11] ^ in_1[11];
  wire        out_0_11 = in_0[11] & in_1[11] | out_xor01_11 & in_2[11];
  wire        out_1_11 = out_xor01_11 ^ in_2[11];
  wire        out_xor01_12 = in_0[12] ^ in_1[12];
  wire        out_0_12 = in_0[12] & in_1[12] | out_xor01_12 & in_2[12];
  wire        out_1_12 = out_xor01_12 ^ in_2[12];
  wire        out_xor01_13 = in_0[13] ^ in_1[13];
  wire        out_0_13 = in_0[13] & in_1[13] | out_xor01_13 & in_2[13];
  wire        out_1_13 = out_xor01_13 ^ in_2[13];
  wire        out_xor01_14 = in_0[14] ^ in_1[14];
  wire        out_0_14 = in_0[14] & in_1[14] | out_xor01_14 & in_2[14];
  wire        out_1_14 = out_xor01_14 ^ in_2[14];
  wire        out_xor01_15 = in_0[15] ^ in_1[15];
  wire        out_0_15 = in_0[15] & in_1[15] | out_xor01_15 & in_2[15];
  wire        out_1_15 = out_xor01_15 ^ in_2[15];
  wire        out_xor01_16 = in_0[16] ^ in_1[16];
  wire        out_0_16 = in_0[16] & in_1[16] | out_xor01_16 & in_2[16];
  wire        out_1_16 = out_xor01_16 ^ in_2[16];
  wire        out_xor01_17 = in_0[17] ^ in_1[17];
  wire        out_0_17 = in_0[17] & in_1[17] | out_xor01_17 & in_2[17];
  wire        out_1_17 = out_xor01_17 ^ in_2[17];
  wire        out_xor01_18 = in_0[18] ^ in_1[18];
  wire        out_0_18 = in_0[18] & in_1[18] | out_xor01_18 & in_2[18];
  wire        out_1_18 = out_xor01_18 ^ in_2[18];
  wire        out_xor01_19 = in_0[19] ^ in_1[19];
  wire        out_0_19 = in_0[19] & in_1[19] | out_xor01_19 & in_2[19];
  wire        out_1_19 = out_xor01_19 ^ in_2[19];
  wire        out_xor01_20 = in_0[20] ^ in_1[20];
  wire        out_0_20 = in_0[20] & in_1[20] | out_xor01_20 & in_2[20];
  wire        out_1_20 = out_xor01_20 ^ in_2[20];
  wire        out_xor01_21 = in_0[21] ^ in_1[21];
  wire        out_0_21 = in_0[21] & in_1[21] | out_xor01_21 & in_2[21];
  wire        out_1_21 = out_xor01_21 ^ in_2[21];
  wire        out_xor01_22 = in_0[22] ^ in_1[22];
  wire        out_0_22 = in_0[22] & in_1[22] | out_xor01_22 & in_2[22];
  wire        out_1_22 = out_xor01_22 ^ in_2[22];
  wire        out_xor01_23 = in_0[23] ^ in_1[23];
  wire        out_0_23 = in_0[23] & in_1[23] | out_xor01_23 & in_2[23];
  wire        out_1_23 = out_xor01_23 ^ in_2[23];
  wire        out_xor01_24 = in_0[24] ^ in_1[24];
  wire        out_0_24 = in_0[24] & in_1[24] | out_xor01_24 & in_2[24];
  wire        out_1_24 = out_xor01_24 ^ in_2[24];
  wire        out_xor01_25 = in_0[25] ^ in_1[25];
  wire        out_0_25 = in_0[25] & in_1[25] | out_xor01_25 & in_2[25];
  wire        out_1_25 = out_xor01_25 ^ in_2[25];
  wire        out_xor01_26 = in_0[26] ^ in_1[26];
  wire        out_0_26 = in_0[26] & in_1[26] | out_xor01_26 & in_2[26];
  wire        out_1_26 = out_xor01_26 ^ in_2[26];
  wire        out_xor01_27 = in_0[27] ^ in_1[27];
  wire        out_0_27 = in_0[27] & in_1[27] | out_xor01_27 & in_2[27];
  wire        out_1_27 = out_xor01_27 ^ in_2[27];
  wire [1:0]  out_0_lo_lo_lo_hi = {out_0_2, out_0_1};
  wire [2:0]  out_0_lo_lo_lo = {out_0_lo_lo_lo_hi, out_0_0};
  wire [1:0]  out_0_lo_lo_hi_lo = {out_0_4, out_0_3};
  wire [1:0]  out_0_lo_lo_hi_hi = {out_0_6, out_0_5};
  wire [3:0]  out_0_lo_lo_hi = {out_0_lo_lo_hi_hi, out_0_lo_lo_hi_lo};
  wire [6:0]  out_0_lo_lo = {out_0_lo_lo_hi, out_0_lo_lo_lo};
  wire [1:0]  out_0_lo_hi_lo_hi = {out_0_9, out_0_8};
  wire [2:0]  out_0_lo_hi_lo = {out_0_lo_hi_lo_hi, out_0_7};
  wire [1:0]  out_0_lo_hi_hi_lo = {out_0_11, out_0_10};
  wire [1:0]  out_0_lo_hi_hi_hi = {out_0_13, out_0_12};
  wire [3:0]  out_0_lo_hi_hi = {out_0_lo_hi_hi_hi, out_0_lo_hi_hi_lo};
  wire [6:0]  out_0_lo_hi = {out_0_lo_hi_hi, out_0_lo_hi_lo};
  wire [13:0] out_0_lo = {out_0_lo_hi, out_0_lo_lo};
  wire [1:0]  out_0_hi_lo_lo_hi = {out_0_16, out_0_15};
  wire [2:0]  out_0_hi_lo_lo = {out_0_hi_lo_lo_hi, out_0_14};
  wire [1:0]  out_0_hi_lo_hi_lo = {out_0_18, out_0_17};
  wire [1:0]  out_0_hi_lo_hi_hi = {out_0_20, out_0_19};
  wire [3:0]  out_0_hi_lo_hi = {out_0_hi_lo_hi_hi, out_0_hi_lo_hi_lo};
  wire [6:0]  out_0_hi_lo = {out_0_hi_lo_hi, out_0_hi_lo_lo};
  wire [1:0]  out_0_hi_hi_lo_hi = {out_0_23, out_0_22};
  wire [2:0]  out_0_hi_hi_lo = {out_0_hi_hi_lo_hi, out_0_21};
  wire [1:0]  out_0_hi_hi_hi_lo = {out_0_25, out_0_24};
  wire [1:0]  out_0_hi_hi_hi_hi = {out_0_27, out_0_26};
  wire [3:0]  out_0_hi_hi_hi = {out_0_hi_hi_hi_hi, out_0_hi_hi_hi_lo};
  wire [6:0]  out_0_hi_hi = {out_0_hi_hi_hi, out_0_hi_hi_lo};
  wire [13:0] out_0_hi = {out_0_hi_hi, out_0_hi_lo};
  wire [1:0]  out_1_lo_lo_lo_hi = {out_1_2, out_1_1};
  wire [2:0]  out_1_lo_lo_lo = {out_1_lo_lo_lo_hi, out_1_0};
  wire [1:0]  out_1_lo_lo_hi_lo = {out_1_4, out_1_3};
  wire [1:0]  out_1_lo_lo_hi_hi = {out_1_6, out_1_5};
  wire [3:0]  out_1_lo_lo_hi = {out_1_lo_lo_hi_hi, out_1_lo_lo_hi_lo};
  wire [6:0]  out_1_lo_lo = {out_1_lo_lo_hi, out_1_lo_lo_lo};
  wire [1:0]  out_1_lo_hi_lo_hi = {out_1_9, out_1_8};
  wire [2:0]  out_1_lo_hi_lo = {out_1_lo_hi_lo_hi, out_1_7};
  wire [1:0]  out_1_lo_hi_hi_lo = {out_1_11, out_1_10};
  wire [1:0]  out_1_lo_hi_hi_hi = {out_1_13, out_1_12};
  wire [3:0]  out_1_lo_hi_hi = {out_1_lo_hi_hi_hi, out_1_lo_hi_hi_lo};
  wire [6:0]  out_1_lo_hi = {out_1_lo_hi_hi, out_1_lo_hi_lo};
  wire [13:0] out_1_lo = {out_1_lo_hi, out_1_lo_lo};
  wire [1:0]  out_1_hi_lo_lo_hi = {out_1_16, out_1_15};
  wire [2:0]  out_1_hi_lo_lo = {out_1_hi_lo_lo_hi, out_1_14};
  wire [1:0]  out_1_hi_lo_hi_lo = {out_1_18, out_1_17};
  wire [1:0]  out_1_hi_lo_hi_hi = {out_1_20, out_1_19};
  wire [3:0]  out_1_hi_lo_hi = {out_1_hi_lo_hi_hi, out_1_hi_lo_hi_lo};
  wire [6:0]  out_1_hi_lo = {out_1_hi_lo_hi, out_1_hi_lo_lo};
  wire [1:0]  out_1_hi_hi_lo_hi = {out_1_23, out_1_22};
  wire [2:0]  out_1_hi_hi_lo = {out_1_hi_hi_lo_hi, out_1_21};
  wire [1:0]  out_1_hi_hi_hi_lo = {out_1_25, out_1_24};
  wire [1:0]  out_1_hi_hi_hi_hi = {out_1_27, out_1_26};
  wire [3:0]  out_1_hi_hi_hi = {out_1_hi_hi_hi_hi, out_1_hi_hi_hi_lo};
  wire [6:0]  out_1_hi_hi = {out_1_hi_hi_hi, out_1_hi_hi_lo};
  wire [13:0] out_1_hi = {out_1_hi_hi, out_1_hi_lo};
  assign out_0 = {out_0_hi, out_0_lo};
  assign out_1 = {out_1_hi, out_1_lo};
endmodule

