
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskCompress(
  input          clock,
                 reset,
                 in_valid,
                 in_bits_maskType,
  input  [1:0]   in_bits_eew,
  input  [2:0]   in_bits_uop,
  input  [31:0]  in_bits_readFromScalar,
                 in_bits_source1,
                 in_bits_mask,
  input  [255:0] in_bits_source2,
                 in_bits_pipeData,
  input  [5:0]   in_bits_groupCounter,
  input  [7:0]   in_bits_ffoInput,
                 in_bits_validInput,
  input          in_bits_lastCompress,
  output [255:0] out_data,
  output [31:0]  out_mask,
  output [5:0]   out_groupCounter,
  output [7:0]   out_ffoOutput,
  output         out_compressValid,
  input          newInstruction,
                 ffoInstruction,
  output [31:0]  writeData,
  output         stageValid
);

  wire         compressDataVec_useTail_31 = 1'h0;
  wire         compressTailMask_elementValid_31 = 1'h0;
  reg          in_1_valid;
  reg          in_1_bits_maskType;
  reg  [1:0]   in_1_bits_eew;
  reg  [2:0]   in_1_bits_uop;
  reg  [31:0]  in_1_bits_readFromScalar;
  reg  [31:0]  in_1_bits_source1;
  reg  [31:0]  in_1_bits_mask;
  reg  [255:0] in_1_bits_source2;
  reg  [255:0] in_1_bits_pipeData;
  reg  [5:0]   in_1_bits_groupCounter;
  reg  [7:0]   in_1_bits_ffoInput;
  reg  [7:0]   in_1_bits_validInput;
  reg          in_1_bits_lastCompress;
  wire         compress = in_1_bits_uop == 3'h1;
  wire         viota = in_1_bits_uop == 3'h0;
  wire         mv = in_1_bits_uop == 3'h2;
  wire         mvRd = in_1_bits_uop == 3'h3;
  wire         writeRD = &(in_1_bits_uop[1:0]);
  wire         ffoType = &(in_1_bits_uop[2:1]);
  wire [3:0]   _eew1H_T = 4'h1 << in_1_bits_eew;
  wire [2:0]   eew1H = _eew1H_T[2:0];
  reg  [9:0]   compressInit;
  wire [9:0]   compressVec_0 = compressInit;
  wire [31:0]  maskInput = in_1_bits_source1 & in_1_bits_mask;
  wire         compressMaskVec_0 = maskInput[0];
  wire         compressMaskVec_1 = maskInput[1];
  wire         compressMaskVec_2 = maskInput[2];
  wire         compressMaskVec_3 = maskInput[3];
  wire         compressMaskVec_4 = maskInput[4];
  wire         compressMaskVec_5 = maskInput[5];
  wire         compressMaskVec_6 = maskInput[6];
  wire         compressMaskVec_7 = maskInput[7];
  wire         compressMaskVec_8 = maskInput[8];
  wire         compressMaskVec_9 = maskInput[9];
  wire         compressMaskVec_10 = maskInput[10];
  wire         compressMaskVec_11 = maskInput[11];
  wire         compressMaskVec_12 = maskInput[12];
  wire         compressMaskVec_13 = maskInput[13];
  wire         compressMaskVec_14 = maskInput[14];
  wire         compressMaskVec_15 = maskInput[15];
  wire         compressMaskVec_16 = maskInput[16];
  wire         compressMaskVec_17 = maskInput[17];
  wire         compressMaskVec_18 = maskInput[18];
  wire         compressMaskVec_19 = maskInput[19];
  wire         compressMaskVec_20 = maskInput[20];
  wire         compressMaskVec_21 = maskInput[21];
  wire         compressMaskVec_22 = maskInput[22];
  wire         compressMaskVec_23 = maskInput[23];
  wire         compressMaskVec_24 = maskInput[24];
  wire         compressMaskVec_25 = maskInput[25];
  wire         compressMaskVec_26 = maskInput[26];
  wire         compressMaskVec_27 = maskInput[27];
  wire         compressMaskVec_28 = maskInput[28];
  wire         compressMaskVec_29 = maskInput[29];
  wire         compressMaskVec_30 = maskInput[30];
  wire         compressMaskVec_31 = maskInput[31];
  wire [9:0]   compressCount =
    compressInit
    + {4'h0,
       {1'h0,
        {1'h0,
         {1'h0, {1'h0, {1'h0, compressMaskVec_0} + {1'h0, compressMaskVec_1}} + {1'h0, {1'h0, compressMaskVec_2} + {1'h0, compressMaskVec_3}}}
           + {1'h0, {1'h0, {1'h0, compressMaskVec_4} + {1'h0, compressMaskVec_5}} + {1'h0, {1'h0, compressMaskVec_6} + {1'h0, compressMaskVec_7}}}}
          + {1'h0,
             {1'h0, {1'h0, {1'h0, compressMaskVec_8} + {1'h0, compressMaskVec_9}} + {1'h0, {1'h0, compressMaskVec_10} + {1'h0, compressMaskVec_11}}}
               + {1'h0, {1'h0, {1'h0, compressMaskVec_12} + {1'h0, compressMaskVec_13}} + {1'h0, {1'h0, compressMaskVec_14} + {1'h0, compressMaskVec_15}}}}}
         + {1'h0,
            {1'h0,
             {1'h0, {1'h0, {1'h0, compressMaskVec_16} + {1'h0, compressMaskVec_17}} + {1'h0, {1'h0, compressMaskVec_18} + {1'h0, compressMaskVec_19}}}
               + {1'h0, {1'h0, {1'h0, compressMaskVec_20} + {1'h0, compressMaskVec_21}} + {1'h0, {1'h0, compressMaskVec_22} + {1'h0, compressMaskVec_23}}}}
              + {1'h0,
                 {1'h0, {1'h0, {1'h0, compressMaskVec_24} + {1'h0, compressMaskVec_25}} + {1'h0, {1'h0, compressMaskVec_26} + {1'h0, compressMaskVec_27}}}
                   + {1'h0, {1'h0, {1'h0, compressMaskVec_28} + {1'h0, compressMaskVec_29}} + {1'h0, {1'h0, compressMaskVec_30} + {1'h0, compressMaskVec_31}}}}}};
  wire [9:0]   compressVec_1 = compressInit + {9'h0, compressMaskVec_0};
  wire [9:0]   compressVec_2 = compressVec_1 + {9'h0, compressMaskVec_1};
  wire [9:0]   compressVec_3 = compressVec_2 + {9'h0, compressMaskVec_2};
  wire [9:0]   compressVec_4 = compressVec_3 + {9'h0, compressMaskVec_3};
  wire [9:0]   compressVec_5 = compressVec_4 + {9'h0, compressMaskVec_4};
  wire [9:0]   compressVec_6 = compressVec_5 + {9'h0, compressMaskVec_5};
  wire [9:0]   compressVec_7 = compressVec_6 + {9'h0, compressMaskVec_6};
  wire [9:0]   compressVec_8 = compressVec_7 + {9'h0, compressMaskVec_7};
  wire [9:0]   compressVec_9 = compressVec_8 + {9'h0, compressMaskVec_8};
  wire [9:0]   compressVec_10 = compressVec_9 + {9'h0, compressMaskVec_9};
  wire [9:0]   compressVec_11 = compressVec_10 + {9'h0, compressMaskVec_10};
  wire [9:0]   compressVec_12 = compressVec_11 + {9'h0, compressMaskVec_11};
  wire [9:0]   compressVec_13 = compressVec_12 + {9'h0, compressMaskVec_12};
  wire [9:0]   compressVec_14 = compressVec_13 + {9'h0, compressMaskVec_13};
  wire [9:0]   compressVec_15 = compressVec_14 + {9'h0, compressMaskVec_14};
  wire [9:0]   compressVec_16 = compressVec_15 + {9'h0, compressMaskVec_15};
  wire [9:0]   compressVec_17 = compressVec_16 + {9'h0, compressMaskVec_16};
  wire [9:0]   compressVec_18 = compressVec_17 + {9'h0, compressMaskVec_17};
  wire [9:0]   compressVec_19 = compressVec_18 + {9'h0, compressMaskVec_18};
  wire [9:0]   compressVec_20 = compressVec_19 + {9'h0, compressMaskVec_19};
  wire [9:0]   compressVec_21 = compressVec_20 + {9'h0, compressMaskVec_20};
  wire [9:0]   compressVec_22 = compressVec_21 + {9'h0, compressMaskVec_21};
  wire [9:0]   compressVec_23 = compressVec_22 + {9'h0, compressMaskVec_22};
  wire [9:0]   compressVec_24 = compressVec_23 + {9'h0, compressMaskVec_23};
  wire [9:0]   compressVec_25 = compressVec_24 + {9'h0, compressMaskVec_24};
  wire [9:0]   compressVec_26 = compressVec_25 + {9'h0, compressMaskVec_25};
  wire [9:0]   compressVec_27 = compressVec_26 + {9'h0, compressMaskVec_26};
  wire [9:0]   compressVec_28 = compressVec_27 + {9'h0, compressMaskVec_27};
  wire [9:0]   compressVec_29 = compressVec_28 + {9'h0, compressMaskVec_28};
  wire [9:0]   compressVec_30 = compressVec_29 + {9'h0, compressMaskVec_29};
  wire [9:0]   compressVec_31 = compressVec_30 + {9'h0, compressMaskVec_30};
  reg  [31:0]  ffoIndex;
  reg          ffoValid;
  wire         countSplit_0_1 = compressCount[5];
  wire [4:0]   countSplit_0_2 = compressCount[4:0];
  wire         countSplit_1_1 = compressCount[4];
  wire [3:0]   countSplit_1_2 = compressCount[3:0];
  wire         countSplit_2_1 = compressCount[3];
  wire [2:0]   countSplit_2_2 = compressCount[2:0];
  wire         compressDeqValid = eew1H[0] & countSplit_0_1 | eew1H[1] & countSplit_1_1 | eew1H[2] & countSplit_2_1 | ~compress;
  wire [4:0]   _compressCountSelect_T_3 = eew1H[0] ? countSplit_0_2 : 5'h0;
  wire [3:0]   _GEN = _compressCountSelect_T_3[3:0] | (eew1H[1] ? countSplit_1_2 : 4'h0);
  wire [4:0]   compressCountSelect = {_compressCountSelect_T_3[4], _GEN[3], _GEN[2:0] | (eew1H[2] ? countSplit_2_2 : 3'h0)};
  reg  [9:0]   compressVecPipe_0;
  reg  [9:0]   compressVecPipe_1;
  reg  [9:0]   compressVecPipe_2;
  reg  [9:0]   compressVecPipe_3;
  reg  [9:0]   compressVecPipe_4;
  reg  [9:0]   compressVecPipe_5;
  reg  [9:0]   compressVecPipe_6;
  reg  [9:0]   compressVecPipe_7;
  reg  [9:0]   compressVecPipe_8;
  reg  [9:0]   compressVecPipe_9;
  reg  [9:0]   compressVecPipe_10;
  reg  [9:0]   compressVecPipe_11;
  reg  [9:0]   compressVecPipe_12;
  reg  [9:0]   compressVecPipe_13;
  reg  [9:0]   compressVecPipe_14;
  reg  [9:0]   compressVecPipe_15;
  reg  [9:0]   compressVecPipe_16;
  reg  [9:0]   compressVecPipe_17;
  reg  [9:0]   compressVecPipe_18;
  reg  [9:0]   compressVecPipe_19;
  reg  [9:0]   compressVecPipe_20;
  reg  [9:0]   compressVecPipe_21;
  reg  [9:0]   compressVecPipe_22;
  reg  [9:0]   compressVecPipe_23;
  reg  [9:0]   compressVecPipe_24;
  reg  [9:0]   compressVecPipe_25;
  reg  [9:0]   compressVecPipe_26;
  reg  [9:0]   compressVecPipe_27;
  reg  [9:0]   compressVecPipe_28;
  reg  [9:0]   compressVecPipe_29;
  reg  [9:0]   compressVecPipe_30;
  reg  [9:0]   compressVecPipe_31;
  reg          compressMaskVecPipe_0;
  reg          compressMaskVecPipe_1;
  reg          compressMaskVecPipe_2;
  reg          compressMaskVecPipe_3;
  reg          compressMaskVecPipe_4;
  reg          compressMaskVecPipe_5;
  reg          compressMaskVecPipe_6;
  reg          compressMaskVecPipe_7;
  reg          compressMaskVecPipe_8;
  reg          compressMaskVecPipe_9;
  reg          compressMaskVecPipe_10;
  reg          compressMaskVecPipe_11;
  reg          compressMaskVecPipe_12;
  reg          compressMaskVecPipe_13;
  reg          compressMaskVecPipe_14;
  reg          compressMaskVecPipe_15;
  reg          compressMaskVecPipe_16;
  reg          compressMaskVecPipe_17;
  reg          compressMaskVecPipe_18;
  reg          compressMaskVecPipe_19;
  reg          compressMaskVecPipe_20;
  reg          compressMaskVecPipe_21;
  reg          compressMaskVecPipe_22;
  reg          compressMaskVecPipe_23;
  reg          compressMaskVecPipe_24;
  reg          compressMaskVecPipe_25;
  reg          compressMaskVecPipe_26;
  reg          compressMaskVecPipe_27;
  reg          compressMaskVecPipe_28;
  reg          compressMaskVecPipe_29;
  reg          compressMaskVecPipe_30;
  reg          compressMaskVecPipe_31;
  reg  [31:0]  maskPipe;
  reg  [255:0] source2Pipe;
  reg          lastCompressPipe;
  reg          stage2Valid;
  reg          newInstructionPipe;
  reg  [9:0]   compressInitPipe;
  reg          compressDeqValidPipe;
  reg  [5:0]   groupCounterPipe;
  wire [7:0]   viotaResult_res_0 = compressVecPipe_0[7:0];
  wire [7:0]   viotaResult_res_1 = compressVecPipe_1[7:0];
  wire [7:0]   viotaResult_res_2 = compressVecPipe_2[7:0];
  wire [7:0]   viotaResult_res_3 = compressVecPipe_3[7:0];
  wire [15:0]  viotaResult_lo = {viotaResult_res_1, viotaResult_res_0};
  wire [15:0]  viotaResult_hi = {viotaResult_res_3, viotaResult_res_2};
  wire [7:0]   viotaResult_res_0_1 = compressVecPipe_4[7:0];
  wire [7:0]   viotaResult_res_1_1 = compressVecPipe_5[7:0];
  wire [7:0]   viotaResult_res_2_1 = compressVecPipe_6[7:0];
  wire [7:0]   viotaResult_res_3_1 = compressVecPipe_7[7:0];
  wire [15:0]  viotaResult_lo_1 = {viotaResult_res_1_1, viotaResult_res_0_1};
  wire [15:0]  viotaResult_hi_1 = {viotaResult_res_3_1, viotaResult_res_2_1};
  wire [7:0]   viotaResult_res_0_2 = compressVecPipe_8[7:0];
  wire [7:0]   viotaResult_res_1_2 = compressVecPipe_9[7:0];
  wire [7:0]   viotaResult_res_2_2 = compressVecPipe_10[7:0];
  wire [7:0]   viotaResult_res_3_2 = compressVecPipe_11[7:0];
  wire [15:0]  viotaResult_lo_2 = {viotaResult_res_1_2, viotaResult_res_0_2};
  wire [15:0]  viotaResult_hi_2 = {viotaResult_res_3_2, viotaResult_res_2_2};
  wire [7:0]   viotaResult_res_0_3 = compressVecPipe_12[7:0];
  wire [7:0]   viotaResult_res_1_3 = compressVecPipe_13[7:0];
  wire [7:0]   viotaResult_res_2_3 = compressVecPipe_14[7:0];
  wire [7:0]   viotaResult_res_3_3 = compressVecPipe_15[7:0];
  wire [15:0]  viotaResult_lo_3 = {viotaResult_res_1_3, viotaResult_res_0_3};
  wire [15:0]  viotaResult_hi_3 = {viotaResult_res_3_3, viotaResult_res_2_3};
  wire [7:0]   viotaResult_res_0_4 = compressVecPipe_16[7:0];
  wire [7:0]   viotaResult_res_1_4 = compressVecPipe_17[7:0];
  wire [7:0]   viotaResult_res_2_4 = compressVecPipe_18[7:0];
  wire [7:0]   viotaResult_res_3_4 = compressVecPipe_19[7:0];
  wire [15:0]  viotaResult_lo_4 = {viotaResult_res_1_4, viotaResult_res_0_4};
  wire [15:0]  viotaResult_hi_4 = {viotaResult_res_3_4, viotaResult_res_2_4};
  wire [7:0]   viotaResult_res_0_5 = compressVecPipe_20[7:0];
  wire [7:0]   viotaResult_res_1_5 = compressVecPipe_21[7:0];
  wire [7:0]   viotaResult_res_2_5 = compressVecPipe_22[7:0];
  wire [7:0]   viotaResult_res_3_5 = compressVecPipe_23[7:0];
  wire [15:0]  viotaResult_lo_5 = {viotaResult_res_1_5, viotaResult_res_0_5};
  wire [15:0]  viotaResult_hi_5 = {viotaResult_res_3_5, viotaResult_res_2_5};
  wire [7:0]   viotaResult_res_0_6 = compressVecPipe_24[7:0];
  wire [7:0]   viotaResult_res_1_6 = compressVecPipe_25[7:0];
  wire [7:0]   viotaResult_res_2_6 = compressVecPipe_26[7:0];
  wire [7:0]   viotaResult_res_3_6 = compressVecPipe_27[7:0];
  wire [15:0]  viotaResult_lo_6 = {viotaResult_res_1_6, viotaResult_res_0_6};
  wire [15:0]  viotaResult_hi_6 = {viotaResult_res_3_6, viotaResult_res_2_6};
  wire [7:0]   viotaResult_res_0_7 = compressVecPipe_28[7:0];
  wire [7:0]   viotaResult_res_1_7 = compressVecPipe_29[7:0];
  wire [7:0]   viotaResult_res_2_7 = compressVecPipe_30[7:0];
  wire [7:0]   viotaResult_res_3_7 = compressVecPipe_31[7:0];
  wire [15:0]  viotaResult_lo_7 = {viotaResult_res_1_7, viotaResult_res_0_7};
  wire [15:0]  viotaResult_hi_7 = {viotaResult_res_3_7, viotaResult_res_2_7};
  wire [63:0]  viotaResult_lo_lo = {viotaResult_hi_1, viotaResult_lo_1, viotaResult_hi, viotaResult_lo};
  wire [63:0]  viotaResult_lo_hi = {viotaResult_hi_3, viotaResult_lo_3, viotaResult_hi_2, viotaResult_lo_2};
  wire [127:0] viotaResult_lo_8 = {viotaResult_lo_hi, viotaResult_lo_lo};
  wire [63:0]  viotaResult_hi_lo = {viotaResult_hi_5, viotaResult_lo_5, viotaResult_hi_4, viotaResult_lo_4};
  wire [63:0]  viotaResult_hi_hi = {viotaResult_hi_7, viotaResult_lo_7, viotaResult_hi_6, viotaResult_lo_6};
  wire [127:0] viotaResult_hi_8 = {viotaResult_hi_hi, viotaResult_hi_lo};
  wire [15:0]  viotaResult_res_0_8 = {6'h0, compressVecPipe_0};
  wire [15:0]  viotaResult_res_1_8 = {6'h0, compressVecPipe_1};
  wire [15:0]  viotaResult_res_0_9 = {6'h0, compressVecPipe_2};
  wire [15:0]  viotaResult_res_1_9 = {6'h0, compressVecPipe_3};
  wire [15:0]  viotaResult_res_0_10 = {6'h0, compressVecPipe_4};
  wire [15:0]  viotaResult_res_1_10 = {6'h0, compressVecPipe_5};
  wire [15:0]  viotaResult_res_0_11 = {6'h0, compressVecPipe_6};
  wire [15:0]  viotaResult_res_1_11 = {6'h0, compressVecPipe_7};
  wire [15:0]  viotaResult_res_0_12 = {6'h0, compressVecPipe_8};
  wire [15:0]  viotaResult_res_1_12 = {6'h0, compressVecPipe_9};
  wire [15:0]  viotaResult_res_0_13 = {6'h0, compressVecPipe_10};
  wire [15:0]  viotaResult_res_1_13 = {6'h0, compressVecPipe_11};
  wire [15:0]  viotaResult_res_0_14 = {6'h0, compressVecPipe_12};
  wire [15:0]  viotaResult_res_1_14 = {6'h0, compressVecPipe_13};
  wire [15:0]  viotaResult_res_0_15 = {6'h0, compressVecPipe_14};
  wire [15:0]  viotaResult_res_1_15 = {6'h0, compressVecPipe_15};
  wire [63:0]  viotaResult_lo_lo_1 = {viotaResult_res_1_9, viotaResult_res_0_9, viotaResult_res_1_8, viotaResult_res_0_8};
  wire [63:0]  viotaResult_lo_hi_1 = {viotaResult_res_1_11, viotaResult_res_0_11, viotaResult_res_1_10, viotaResult_res_0_10};
  wire [127:0] viotaResult_lo_9 = {viotaResult_lo_hi_1, viotaResult_lo_lo_1};
  wire [63:0]  viotaResult_hi_lo_1 = {viotaResult_res_1_13, viotaResult_res_0_13, viotaResult_res_1_12, viotaResult_res_0_12};
  wire [63:0]  viotaResult_hi_hi_1 = {viotaResult_res_1_15, viotaResult_res_0_15, viotaResult_res_1_14, viotaResult_res_0_14};
  wire [127:0] viotaResult_hi_9 = {viotaResult_hi_hi_1, viotaResult_hi_lo_1};
  wire [31:0]  viotaResult_res_0_16 = {22'h0, compressVecPipe_0};
  wire [31:0]  viotaResult_res_0_17 = {22'h0, compressVecPipe_1};
  wire [31:0]  viotaResult_res_0_18 = {22'h0, compressVecPipe_2};
  wire [31:0]  viotaResult_res_0_19 = {22'h0, compressVecPipe_3};
  wire [31:0]  viotaResult_res_0_20 = {22'h0, compressVecPipe_4};
  wire [31:0]  viotaResult_res_0_21 = {22'h0, compressVecPipe_5};
  wire [31:0]  viotaResult_res_0_22 = {22'h0, compressVecPipe_6};
  wire [31:0]  viotaResult_res_0_23 = {22'h0, compressVecPipe_7};
  wire [63:0]  viotaResult_lo_lo_2 = {viotaResult_res_0_17, viotaResult_res_0_16};
  wire [63:0]  viotaResult_lo_hi_2 = {viotaResult_res_0_19, viotaResult_res_0_18};
  wire [127:0] viotaResult_lo_10 = {viotaResult_lo_hi_2, viotaResult_lo_lo_2};
  wire [63:0]  viotaResult_hi_lo_2 = {viotaResult_res_0_21, viotaResult_res_0_20};
  wire [63:0]  viotaResult_hi_hi_2 = {viotaResult_res_0_23, viotaResult_res_0_22};
  wire [127:0] viotaResult_hi_10 = {viotaResult_hi_hi_2, viotaResult_hi_lo_2};
  wire [255:0] viotaResult = (eew1H[0] ? {viotaResult_hi_8, viotaResult_lo_8} : 256'h0) | (eew1H[1] ? {viotaResult_hi_9, viotaResult_lo_9} : 256'h0) | (eew1H[2] ? {viotaResult_hi_10, viotaResult_lo_10} : 256'h0);
  wire         viotaMask_res_0 = maskPipe[0];
  wire         viotaMask_res_1 = maskPipe[1];
  wire         viotaMask_res_2 = maskPipe[2];
  wire         viotaMask_res_3 = maskPipe[3];
  wire [1:0]   viotaMask_lo = {viotaMask_res_1, viotaMask_res_0};
  wire [1:0]   viotaMask_hi = {viotaMask_res_3, viotaMask_res_2};
  wire         viotaMask_res_0_1 = maskPipe[4];
  wire         viotaMask_res_1_1 = maskPipe[5];
  wire         viotaMask_res_2_1 = maskPipe[6];
  wire         viotaMask_res_3_1 = maskPipe[7];
  wire [1:0]   viotaMask_lo_1 = {viotaMask_res_1_1, viotaMask_res_0_1};
  wire [1:0]   viotaMask_hi_1 = {viotaMask_res_3_1, viotaMask_res_2_1};
  wire         viotaMask_res_0_2 = maskPipe[8];
  wire         viotaMask_res_1_2 = maskPipe[9];
  wire         viotaMask_res_2_2 = maskPipe[10];
  wire         viotaMask_res_3_2 = maskPipe[11];
  wire [1:0]   viotaMask_lo_2 = {viotaMask_res_1_2, viotaMask_res_0_2};
  wire [1:0]   viotaMask_hi_2 = {viotaMask_res_3_2, viotaMask_res_2_2};
  wire         viotaMask_res_0_3 = maskPipe[12];
  wire         viotaMask_res_1_3 = maskPipe[13];
  wire         viotaMask_res_2_3 = maskPipe[14];
  wire         viotaMask_res_3_3 = maskPipe[15];
  wire [1:0]   viotaMask_lo_3 = {viotaMask_res_1_3, viotaMask_res_0_3};
  wire [1:0]   viotaMask_hi_3 = {viotaMask_res_3_3, viotaMask_res_2_3};
  wire         viotaMask_res_0_4 = maskPipe[16];
  wire         viotaMask_res_1_4 = maskPipe[17];
  wire         viotaMask_res_2_4 = maskPipe[18];
  wire         viotaMask_res_3_4 = maskPipe[19];
  wire [1:0]   viotaMask_lo_4 = {viotaMask_res_1_4, viotaMask_res_0_4};
  wire [1:0]   viotaMask_hi_4 = {viotaMask_res_3_4, viotaMask_res_2_4};
  wire         viotaMask_res_0_5 = maskPipe[20];
  wire         viotaMask_res_1_5 = maskPipe[21];
  wire         viotaMask_res_2_5 = maskPipe[22];
  wire         viotaMask_res_3_5 = maskPipe[23];
  wire [1:0]   viotaMask_lo_5 = {viotaMask_res_1_5, viotaMask_res_0_5};
  wire [1:0]   viotaMask_hi_5 = {viotaMask_res_3_5, viotaMask_res_2_5};
  wire         viotaMask_res_0_6 = maskPipe[24];
  wire         viotaMask_res_1_6 = maskPipe[25];
  wire         viotaMask_res_2_6 = maskPipe[26];
  wire         viotaMask_res_3_6 = maskPipe[27];
  wire [1:0]   viotaMask_lo_6 = {viotaMask_res_1_6, viotaMask_res_0_6};
  wire [1:0]   viotaMask_hi_6 = {viotaMask_res_3_6, viotaMask_res_2_6};
  wire         viotaMask_res_0_7 = maskPipe[28];
  wire         viotaMask_res_1_7 = maskPipe[29];
  wire         viotaMask_res_2_7 = maskPipe[30];
  wire         viotaMask_res_3_7 = maskPipe[31];
  wire [1:0]   viotaMask_lo_7 = {viotaMask_res_1_7, viotaMask_res_0_7};
  wire [1:0]   viotaMask_hi_7 = {viotaMask_res_3_7, viotaMask_res_2_7};
  wire [7:0]   viotaMask_lo_lo = {viotaMask_hi_1, viotaMask_lo_1, viotaMask_hi, viotaMask_lo};
  wire [7:0]   viotaMask_lo_hi = {viotaMask_hi_3, viotaMask_lo_3, viotaMask_hi_2, viotaMask_lo_2};
  wire [15:0]  viotaMask_lo_8 = {viotaMask_lo_hi, viotaMask_lo_lo};
  wire [7:0]   viotaMask_hi_lo = {viotaMask_hi_5, viotaMask_lo_5, viotaMask_hi_4, viotaMask_lo_4};
  wire [7:0]   viotaMask_hi_hi = {viotaMask_hi_7, viotaMask_lo_7, viotaMask_hi_6, viotaMask_lo_6};
  wire [15:0]  viotaMask_hi_8 = {viotaMask_hi_hi, viotaMask_hi_lo};
  wire [1:0]   viotaMask_res_0_8 = {2{viotaMask_res_0}};
  wire [1:0]   viotaMask_res_1_8 = {2{viotaMask_res_1}};
  wire [1:0]   viotaMask_res_0_9 = {2{viotaMask_res_2}};
  wire [1:0]   viotaMask_res_1_9 = {2{viotaMask_res_3}};
  wire [1:0]   viotaMask_res_0_10 = {2{viotaMask_res_0_1}};
  wire [1:0]   viotaMask_res_1_10 = {2{viotaMask_res_1_1}};
  wire [1:0]   viotaMask_res_0_11 = {2{viotaMask_res_2_1}};
  wire [1:0]   viotaMask_res_1_11 = {2{viotaMask_res_3_1}};
  wire [1:0]   viotaMask_res_0_12 = {2{viotaMask_res_0_2}};
  wire [1:0]   viotaMask_res_1_12 = {2{viotaMask_res_1_2}};
  wire [1:0]   viotaMask_res_0_13 = {2{viotaMask_res_2_2}};
  wire [1:0]   viotaMask_res_1_13 = {2{viotaMask_res_3_2}};
  wire [1:0]   viotaMask_res_0_14 = {2{viotaMask_res_0_3}};
  wire [1:0]   viotaMask_res_1_14 = {2{viotaMask_res_1_3}};
  wire [1:0]   viotaMask_res_0_15 = {2{viotaMask_res_2_3}};
  wire [1:0]   viotaMask_res_1_15 = {2{viotaMask_res_3_3}};
  wire [7:0]   viotaMask_lo_lo_1 = {viotaMask_res_1_9, viotaMask_res_0_9, viotaMask_res_1_8, viotaMask_res_0_8};
  wire [7:0]   viotaMask_lo_hi_1 = {viotaMask_res_1_11, viotaMask_res_0_11, viotaMask_res_1_10, viotaMask_res_0_10};
  wire [15:0]  viotaMask_lo_9 = {viotaMask_lo_hi_1, viotaMask_lo_lo_1};
  wire [7:0]   viotaMask_hi_lo_1 = {viotaMask_res_1_13, viotaMask_res_0_13, viotaMask_res_1_12, viotaMask_res_0_12};
  wire [7:0]   viotaMask_hi_hi_1 = {viotaMask_res_1_15, viotaMask_res_0_15, viotaMask_res_1_14, viotaMask_res_0_14};
  wire [15:0]  viotaMask_hi_9 = {viotaMask_hi_hi_1, viotaMask_hi_lo_1};
  wire [3:0]   viotaMask_res_0_16 = {4{viotaMask_res_0}};
  wire [3:0]   viotaMask_res_0_17 = {4{viotaMask_res_1}};
  wire [3:0]   viotaMask_res_0_18 = {4{viotaMask_res_2}};
  wire [3:0]   viotaMask_res_0_19 = {4{viotaMask_res_3}};
  wire [3:0]   viotaMask_res_0_20 = {4{viotaMask_res_0_1}};
  wire [3:0]   viotaMask_res_0_21 = {4{viotaMask_res_1_1}};
  wire [3:0]   viotaMask_res_0_22 = {4{viotaMask_res_2_1}};
  wire [3:0]   viotaMask_res_0_23 = {4{viotaMask_res_3_1}};
  wire [7:0]   viotaMask_lo_lo_2 = {viotaMask_res_0_17, viotaMask_res_0_16};
  wire [7:0]   viotaMask_lo_hi_2 = {viotaMask_res_0_19, viotaMask_res_0_18};
  wire [15:0]  viotaMask_lo_10 = {viotaMask_lo_hi_2, viotaMask_lo_lo_2};
  wire [7:0]   viotaMask_hi_lo_2 = {viotaMask_res_0_21, viotaMask_res_0_20};
  wire [7:0]   viotaMask_hi_hi_2 = {viotaMask_res_0_23, viotaMask_res_0_22};
  wire [15:0]  viotaMask_hi_10 = {viotaMask_hi_hi_2, viotaMask_hi_lo_2};
  wire [31:0]  viotaMask = (eew1H[0] ? {viotaMask_hi_8, viotaMask_lo_8} : 32'h0) | (eew1H[1] ? {viotaMask_hi_9, viotaMask_lo_9} : 32'h0) | (eew1H[2] ? {viotaMask_hi_10, viotaMask_lo_10} : 32'h0);
  wire [4:0]   tailCount = compressInitPipe[4:0];
  wire [4:0]   tailCountForMask = compressInit[4:0];
  reg  [255:0] compressDataReg;
  reg          compressTailValid;
  reg  [5:0]   compressWriteGroupCount;
  wire         _GEN_0 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h0;
  wire         compressDataVec_hitReq_0;
  assign compressDataVec_hitReq_0 = _GEN_0;
  wire         compressDataVec_hitReq_0_64;
  assign compressDataVec_hitReq_0_64 = _GEN_0;
  wire         compressDataVec_hitReq_0_96;
  assign compressDataVec_hitReq_0_96 = _GEN_0;
  wire         _GEN_1 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h0;
  wire         compressDataVec_hitReq_1;
  assign compressDataVec_hitReq_1 = _GEN_1;
  wire         compressDataVec_hitReq_1_64;
  assign compressDataVec_hitReq_1_64 = _GEN_1;
  wire         compressDataVec_hitReq_1_96;
  assign compressDataVec_hitReq_1_96 = _GEN_1;
  wire         _GEN_2 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h0;
  wire         compressDataVec_hitReq_2;
  assign compressDataVec_hitReq_2 = _GEN_2;
  wire         compressDataVec_hitReq_2_64;
  assign compressDataVec_hitReq_2_64 = _GEN_2;
  wire         compressDataVec_hitReq_2_96;
  assign compressDataVec_hitReq_2_96 = _GEN_2;
  wire         _GEN_3 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h0;
  wire         compressDataVec_hitReq_3;
  assign compressDataVec_hitReq_3 = _GEN_3;
  wire         compressDataVec_hitReq_3_64;
  assign compressDataVec_hitReq_3_64 = _GEN_3;
  wire         compressDataVec_hitReq_3_96;
  assign compressDataVec_hitReq_3_96 = _GEN_3;
  wire         _GEN_4 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h0;
  wire         compressDataVec_hitReq_4;
  assign compressDataVec_hitReq_4 = _GEN_4;
  wire         compressDataVec_hitReq_4_64;
  assign compressDataVec_hitReq_4_64 = _GEN_4;
  wire         compressDataVec_hitReq_4_96;
  assign compressDataVec_hitReq_4_96 = _GEN_4;
  wire         _GEN_5 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h0;
  wire         compressDataVec_hitReq_5;
  assign compressDataVec_hitReq_5 = _GEN_5;
  wire         compressDataVec_hitReq_5_64;
  assign compressDataVec_hitReq_5_64 = _GEN_5;
  wire         compressDataVec_hitReq_5_96;
  assign compressDataVec_hitReq_5_96 = _GEN_5;
  wire         _GEN_6 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h0;
  wire         compressDataVec_hitReq_6;
  assign compressDataVec_hitReq_6 = _GEN_6;
  wire         compressDataVec_hitReq_6_64;
  assign compressDataVec_hitReq_6_64 = _GEN_6;
  wire         compressDataVec_hitReq_6_96;
  assign compressDataVec_hitReq_6_96 = _GEN_6;
  wire         _GEN_7 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h0;
  wire         compressDataVec_hitReq_7;
  assign compressDataVec_hitReq_7 = _GEN_7;
  wire         compressDataVec_hitReq_7_64;
  assign compressDataVec_hitReq_7_64 = _GEN_7;
  wire         compressDataVec_hitReq_7_96;
  assign compressDataVec_hitReq_7_96 = _GEN_7;
  wire         _GEN_8 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h0;
  wire         compressDataVec_hitReq_8;
  assign compressDataVec_hitReq_8 = _GEN_8;
  wire         compressDataVec_hitReq_8_64;
  assign compressDataVec_hitReq_8_64 = _GEN_8;
  wire         _GEN_9 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h0;
  wire         compressDataVec_hitReq_9;
  assign compressDataVec_hitReq_9 = _GEN_9;
  wire         compressDataVec_hitReq_9_64;
  assign compressDataVec_hitReq_9_64 = _GEN_9;
  wire         _GEN_10 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h0;
  wire         compressDataVec_hitReq_10;
  assign compressDataVec_hitReq_10 = _GEN_10;
  wire         compressDataVec_hitReq_10_64;
  assign compressDataVec_hitReq_10_64 = _GEN_10;
  wire         _GEN_11 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h0;
  wire         compressDataVec_hitReq_11;
  assign compressDataVec_hitReq_11 = _GEN_11;
  wire         compressDataVec_hitReq_11_64;
  assign compressDataVec_hitReq_11_64 = _GEN_11;
  wire         _GEN_12 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h0;
  wire         compressDataVec_hitReq_12;
  assign compressDataVec_hitReq_12 = _GEN_12;
  wire         compressDataVec_hitReq_12_64;
  assign compressDataVec_hitReq_12_64 = _GEN_12;
  wire         _GEN_13 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h0;
  wire         compressDataVec_hitReq_13;
  assign compressDataVec_hitReq_13 = _GEN_13;
  wire         compressDataVec_hitReq_13_64;
  assign compressDataVec_hitReq_13_64 = _GEN_13;
  wire         _GEN_14 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h0;
  wire         compressDataVec_hitReq_14;
  assign compressDataVec_hitReq_14 = _GEN_14;
  wire         compressDataVec_hitReq_14_64;
  assign compressDataVec_hitReq_14_64 = _GEN_14;
  wire         _GEN_15 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h0;
  wire         compressDataVec_hitReq_15;
  assign compressDataVec_hitReq_15 = _GEN_15;
  wire         compressDataVec_hitReq_15_64;
  assign compressDataVec_hitReq_15_64 = _GEN_15;
  wire         compressDataVec_hitReq_16 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h0;
  wire         compressDataVec_hitReq_17 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h0;
  wire         compressDataVec_hitReq_18 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h0;
  wire         compressDataVec_hitReq_19 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h0;
  wire         compressDataVec_hitReq_20 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h0;
  wire         compressDataVec_hitReq_21 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h0;
  wire         compressDataVec_hitReq_22 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h0;
  wire         compressDataVec_hitReq_23 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h0;
  wire         compressDataVec_hitReq_24 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h0;
  wire         compressDataVec_hitReq_25 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h0;
  wire         compressDataVec_hitReq_26 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h0;
  wire         compressDataVec_hitReq_27 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h0;
  wire         compressDataVec_hitReq_28 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h0;
  wire         compressDataVec_hitReq_29 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h0;
  wire         compressDataVec_hitReq_30 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h0;
  wire         compressDataVec_hitReq_31 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h0;
  wire [7:0]   compressDataVec_selectReqData =
    (compressDataVec_hitReq_0 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail;
  assign compressDataVec_useTail = |tailCount;
  wire         _GEN_16 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1;
  wire         compressDataVec_hitReq_0_1;
  assign compressDataVec_hitReq_0_1 = _GEN_16;
  wire         compressDataVec_hitReq_0_65;
  assign compressDataVec_hitReq_0_65 = _GEN_16;
  wire         compressDataVec_hitReq_0_97;
  assign compressDataVec_hitReq_0_97 = _GEN_16;
  wire         _GEN_17 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1;
  wire         compressDataVec_hitReq_1_1;
  assign compressDataVec_hitReq_1_1 = _GEN_17;
  wire         compressDataVec_hitReq_1_65;
  assign compressDataVec_hitReq_1_65 = _GEN_17;
  wire         compressDataVec_hitReq_1_97;
  assign compressDataVec_hitReq_1_97 = _GEN_17;
  wire         _GEN_18 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1;
  wire         compressDataVec_hitReq_2_1;
  assign compressDataVec_hitReq_2_1 = _GEN_18;
  wire         compressDataVec_hitReq_2_65;
  assign compressDataVec_hitReq_2_65 = _GEN_18;
  wire         compressDataVec_hitReq_2_97;
  assign compressDataVec_hitReq_2_97 = _GEN_18;
  wire         _GEN_19 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1;
  wire         compressDataVec_hitReq_3_1;
  assign compressDataVec_hitReq_3_1 = _GEN_19;
  wire         compressDataVec_hitReq_3_65;
  assign compressDataVec_hitReq_3_65 = _GEN_19;
  wire         compressDataVec_hitReq_3_97;
  assign compressDataVec_hitReq_3_97 = _GEN_19;
  wire         _GEN_20 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1;
  wire         compressDataVec_hitReq_4_1;
  assign compressDataVec_hitReq_4_1 = _GEN_20;
  wire         compressDataVec_hitReq_4_65;
  assign compressDataVec_hitReq_4_65 = _GEN_20;
  wire         compressDataVec_hitReq_4_97;
  assign compressDataVec_hitReq_4_97 = _GEN_20;
  wire         _GEN_21 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1;
  wire         compressDataVec_hitReq_5_1;
  assign compressDataVec_hitReq_5_1 = _GEN_21;
  wire         compressDataVec_hitReq_5_65;
  assign compressDataVec_hitReq_5_65 = _GEN_21;
  wire         compressDataVec_hitReq_5_97;
  assign compressDataVec_hitReq_5_97 = _GEN_21;
  wire         _GEN_22 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1;
  wire         compressDataVec_hitReq_6_1;
  assign compressDataVec_hitReq_6_1 = _GEN_22;
  wire         compressDataVec_hitReq_6_65;
  assign compressDataVec_hitReq_6_65 = _GEN_22;
  wire         compressDataVec_hitReq_6_97;
  assign compressDataVec_hitReq_6_97 = _GEN_22;
  wire         _GEN_23 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1;
  wire         compressDataVec_hitReq_7_1;
  assign compressDataVec_hitReq_7_1 = _GEN_23;
  wire         compressDataVec_hitReq_7_65;
  assign compressDataVec_hitReq_7_65 = _GEN_23;
  wire         compressDataVec_hitReq_7_97;
  assign compressDataVec_hitReq_7_97 = _GEN_23;
  wire         _GEN_24 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1;
  wire         compressDataVec_hitReq_8_1;
  assign compressDataVec_hitReq_8_1 = _GEN_24;
  wire         compressDataVec_hitReq_8_65;
  assign compressDataVec_hitReq_8_65 = _GEN_24;
  wire         _GEN_25 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1;
  wire         compressDataVec_hitReq_9_1;
  assign compressDataVec_hitReq_9_1 = _GEN_25;
  wire         compressDataVec_hitReq_9_65;
  assign compressDataVec_hitReq_9_65 = _GEN_25;
  wire         _GEN_26 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1;
  wire         compressDataVec_hitReq_10_1;
  assign compressDataVec_hitReq_10_1 = _GEN_26;
  wire         compressDataVec_hitReq_10_65;
  assign compressDataVec_hitReq_10_65 = _GEN_26;
  wire         _GEN_27 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1;
  wire         compressDataVec_hitReq_11_1;
  assign compressDataVec_hitReq_11_1 = _GEN_27;
  wire         compressDataVec_hitReq_11_65;
  assign compressDataVec_hitReq_11_65 = _GEN_27;
  wire         _GEN_28 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1;
  wire         compressDataVec_hitReq_12_1;
  assign compressDataVec_hitReq_12_1 = _GEN_28;
  wire         compressDataVec_hitReq_12_65;
  assign compressDataVec_hitReq_12_65 = _GEN_28;
  wire         _GEN_29 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1;
  wire         compressDataVec_hitReq_13_1;
  assign compressDataVec_hitReq_13_1 = _GEN_29;
  wire         compressDataVec_hitReq_13_65;
  assign compressDataVec_hitReq_13_65 = _GEN_29;
  wire         _GEN_30 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1;
  wire         compressDataVec_hitReq_14_1;
  assign compressDataVec_hitReq_14_1 = _GEN_30;
  wire         compressDataVec_hitReq_14_65;
  assign compressDataVec_hitReq_14_65 = _GEN_30;
  wire         _GEN_31 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1;
  wire         compressDataVec_hitReq_15_1;
  assign compressDataVec_hitReq_15_1 = _GEN_31;
  wire         compressDataVec_hitReq_15_65;
  assign compressDataVec_hitReq_15_65 = _GEN_31;
  wire         compressDataVec_hitReq_16_1 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1;
  wire         compressDataVec_hitReq_17_1 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1;
  wire         compressDataVec_hitReq_18_1 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1;
  wire         compressDataVec_hitReq_19_1 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1;
  wire         compressDataVec_hitReq_20_1 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1;
  wire         compressDataVec_hitReq_21_1 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1;
  wire         compressDataVec_hitReq_22_1 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1;
  wire         compressDataVec_hitReq_23_1 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1;
  wire         compressDataVec_hitReq_24_1 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1;
  wire         compressDataVec_hitReq_25_1 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1;
  wire         compressDataVec_hitReq_26_1 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1;
  wire         compressDataVec_hitReq_27_1 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1;
  wire         compressDataVec_hitReq_28_1 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1;
  wire         compressDataVec_hitReq_29_1 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1;
  wire         compressDataVec_hitReq_30_1 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1;
  wire         compressDataVec_hitReq_31_1 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1;
  wire [7:0]   compressDataVec_selectReqData_1 =
    (compressDataVec_hitReq_0_1 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_1 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_1 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_1 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_1 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_1 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_1 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_1 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_1 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_1 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_1 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_1 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_1 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_1 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_1 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_1 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_1 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_1 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_1 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_1 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_1 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_1 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_1 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_1 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_1 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_1 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_1 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_1 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_1 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_1 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_1 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_1 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_1;
  assign compressDataVec_useTail_1 = |(tailCount[4:1]);
  wire         _GEN_32 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2;
  wire         compressDataVec_hitReq_0_2;
  assign compressDataVec_hitReq_0_2 = _GEN_32;
  wire         compressDataVec_hitReq_0_66;
  assign compressDataVec_hitReq_0_66 = _GEN_32;
  wire         compressDataVec_hitReq_0_98;
  assign compressDataVec_hitReq_0_98 = _GEN_32;
  wire         _GEN_33 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2;
  wire         compressDataVec_hitReq_1_2;
  assign compressDataVec_hitReq_1_2 = _GEN_33;
  wire         compressDataVec_hitReq_1_66;
  assign compressDataVec_hitReq_1_66 = _GEN_33;
  wire         compressDataVec_hitReq_1_98;
  assign compressDataVec_hitReq_1_98 = _GEN_33;
  wire         _GEN_34 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2;
  wire         compressDataVec_hitReq_2_2;
  assign compressDataVec_hitReq_2_2 = _GEN_34;
  wire         compressDataVec_hitReq_2_66;
  assign compressDataVec_hitReq_2_66 = _GEN_34;
  wire         compressDataVec_hitReq_2_98;
  assign compressDataVec_hitReq_2_98 = _GEN_34;
  wire         _GEN_35 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2;
  wire         compressDataVec_hitReq_3_2;
  assign compressDataVec_hitReq_3_2 = _GEN_35;
  wire         compressDataVec_hitReq_3_66;
  assign compressDataVec_hitReq_3_66 = _GEN_35;
  wire         compressDataVec_hitReq_3_98;
  assign compressDataVec_hitReq_3_98 = _GEN_35;
  wire         _GEN_36 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2;
  wire         compressDataVec_hitReq_4_2;
  assign compressDataVec_hitReq_4_2 = _GEN_36;
  wire         compressDataVec_hitReq_4_66;
  assign compressDataVec_hitReq_4_66 = _GEN_36;
  wire         compressDataVec_hitReq_4_98;
  assign compressDataVec_hitReq_4_98 = _GEN_36;
  wire         _GEN_37 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2;
  wire         compressDataVec_hitReq_5_2;
  assign compressDataVec_hitReq_5_2 = _GEN_37;
  wire         compressDataVec_hitReq_5_66;
  assign compressDataVec_hitReq_5_66 = _GEN_37;
  wire         compressDataVec_hitReq_5_98;
  assign compressDataVec_hitReq_5_98 = _GEN_37;
  wire         _GEN_38 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2;
  wire         compressDataVec_hitReq_6_2;
  assign compressDataVec_hitReq_6_2 = _GEN_38;
  wire         compressDataVec_hitReq_6_66;
  assign compressDataVec_hitReq_6_66 = _GEN_38;
  wire         compressDataVec_hitReq_6_98;
  assign compressDataVec_hitReq_6_98 = _GEN_38;
  wire         _GEN_39 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2;
  wire         compressDataVec_hitReq_7_2;
  assign compressDataVec_hitReq_7_2 = _GEN_39;
  wire         compressDataVec_hitReq_7_66;
  assign compressDataVec_hitReq_7_66 = _GEN_39;
  wire         compressDataVec_hitReq_7_98;
  assign compressDataVec_hitReq_7_98 = _GEN_39;
  wire         _GEN_40 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2;
  wire         compressDataVec_hitReq_8_2;
  assign compressDataVec_hitReq_8_2 = _GEN_40;
  wire         compressDataVec_hitReq_8_66;
  assign compressDataVec_hitReq_8_66 = _GEN_40;
  wire         _GEN_41 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2;
  wire         compressDataVec_hitReq_9_2;
  assign compressDataVec_hitReq_9_2 = _GEN_41;
  wire         compressDataVec_hitReq_9_66;
  assign compressDataVec_hitReq_9_66 = _GEN_41;
  wire         _GEN_42 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2;
  wire         compressDataVec_hitReq_10_2;
  assign compressDataVec_hitReq_10_2 = _GEN_42;
  wire         compressDataVec_hitReq_10_66;
  assign compressDataVec_hitReq_10_66 = _GEN_42;
  wire         _GEN_43 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2;
  wire         compressDataVec_hitReq_11_2;
  assign compressDataVec_hitReq_11_2 = _GEN_43;
  wire         compressDataVec_hitReq_11_66;
  assign compressDataVec_hitReq_11_66 = _GEN_43;
  wire         _GEN_44 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2;
  wire         compressDataVec_hitReq_12_2;
  assign compressDataVec_hitReq_12_2 = _GEN_44;
  wire         compressDataVec_hitReq_12_66;
  assign compressDataVec_hitReq_12_66 = _GEN_44;
  wire         _GEN_45 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2;
  wire         compressDataVec_hitReq_13_2;
  assign compressDataVec_hitReq_13_2 = _GEN_45;
  wire         compressDataVec_hitReq_13_66;
  assign compressDataVec_hitReq_13_66 = _GEN_45;
  wire         _GEN_46 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2;
  wire         compressDataVec_hitReq_14_2;
  assign compressDataVec_hitReq_14_2 = _GEN_46;
  wire         compressDataVec_hitReq_14_66;
  assign compressDataVec_hitReq_14_66 = _GEN_46;
  wire         _GEN_47 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2;
  wire         compressDataVec_hitReq_15_2;
  assign compressDataVec_hitReq_15_2 = _GEN_47;
  wire         compressDataVec_hitReq_15_66;
  assign compressDataVec_hitReq_15_66 = _GEN_47;
  wire         compressDataVec_hitReq_16_2 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2;
  wire         compressDataVec_hitReq_17_2 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2;
  wire         compressDataVec_hitReq_18_2 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2;
  wire         compressDataVec_hitReq_19_2 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2;
  wire         compressDataVec_hitReq_20_2 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2;
  wire         compressDataVec_hitReq_21_2 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2;
  wire         compressDataVec_hitReq_22_2 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2;
  wire         compressDataVec_hitReq_23_2 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2;
  wire         compressDataVec_hitReq_24_2 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2;
  wire         compressDataVec_hitReq_25_2 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2;
  wire         compressDataVec_hitReq_26_2 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2;
  wire         compressDataVec_hitReq_27_2 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2;
  wire         compressDataVec_hitReq_28_2 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2;
  wire         compressDataVec_hitReq_29_2 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2;
  wire         compressDataVec_hitReq_30_2 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2;
  wire         compressDataVec_hitReq_31_2 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2;
  wire [7:0]   compressDataVec_selectReqData_2 =
    (compressDataVec_hitReq_0_2 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_2 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_2 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_2 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_2 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_2 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_2 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_2 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_2 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_2 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_2 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_2 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_2 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_2 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_2 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_2 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_2 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_2 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_2 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_2 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_2 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_2 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_2 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_2 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_2 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_2 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_2 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_2 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_2 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_2 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_2 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_2 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_48 = tailCount > 5'h2;
  wire         compressDataVec_useTail_2;
  assign compressDataVec_useTail_2 = _GEN_48;
  wire         compressDataVec_useTail_34;
  assign compressDataVec_useTail_34 = _GEN_48;
  wire         compressDataVec_useTail_50;
  assign compressDataVec_useTail_50 = _GEN_48;
  wire         _GEN_49 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3;
  wire         compressDataVec_hitReq_0_3;
  assign compressDataVec_hitReq_0_3 = _GEN_49;
  wire         compressDataVec_hitReq_0_67;
  assign compressDataVec_hitReq_0_67 = _GEN_49;
  wire         compressDataVec_hitReq_0_99;
  assign compressDataVec_hitReq_0_99 = _GEN_49;
  wire         _GEN_50 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3;
  wire         compressDataVec_hitReq_1_3;
  assign compressDataVec_hitReq_1_3 = _GEN_50;
  wire         compressDataVec_hitReq_1_67;
  assign compressDataVec_hitReq_1_67 = _GEN_50;
  wire         compressDataVec_hitReq_1_99;
  assign compressDataVec_hitReq_1_99 = _GEN_50;
  wire         _GEN_51 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3;
  wire         compressDataVec_hitReq_2_3;
  assign compressDataVec_hitReq_2_3 = _GEN_51;
  wire         compressDataVec_hitReq_2_67;
  assign compressDataVec_hitReq_2_67 = _GEN_51;
  wire         compressDataVec_hitReq_2_99;
  assign compressDataVec_hitReq_2_99 = _GEN_51;
  wire         _GEN_52 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3;
  wire         compressDataVec_hitReq_3_3;
  assign compressDataVec_hitReq_3_3 = _GEN_52;
  wire         compressDataVec_hitReq_3_67;
  assign compressDataVec_hitReq_3_67 = _GEN_52;
  wire         compressDataVec_hitReq_3_99;
  assign compressDataVec_hitReq_3_99 = _GEN_52;
  wire         _GEN_53 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3;
  wire         compressDataVec_hitReq_4_3;
  assign compressDataVec_hitReq_4_3 = _GEN_53;
  wire         compressDataVec_hitReq_4_67;
  assign compressDataVec_hitReq_4_67 = _GEN_53;
  wire         compressDataVec_hitReq_4_99;
  assign compressDataVec_hitReq_4_99 = _GEN_53;
  wire         _GEN_54 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3;
  wire         compressDataVec_hitReq_5_3;
  assign compressDataVec_hitReq_5_3 = _GEN_54;
  wire         compressDataVec_hitReq_5_67;
  assign compressDataVec_hitReq_5_67 = _GEN_54;
  wire         compressDataVec_hitReq_5_99;
  assign compressDataVec_hitReq_5_99 = _GEN_54;
  wire         _GEN_55 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3;
  wire         compressDataVec_hitReq_6_3;
  assign compressDataVec_hitReq_6_3 = _GEN_55;
  wire         compressDataVec_hitReq_6_67;
  assign compressDataVec_hitReq_6_67 = _GEN_55;
  wire         compressDataVec_hitReq_6_99;
  assign compressDataVec_hitReq_6_99 = _GEN_55;
  wire         _GEN_56 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3;
  wire         compressDataVec_hitReq_7_3;
  assign compressDataVec_hitReq_7_3 = _GEN_56;
  wire         compressDataVec_hitReq_7_67;
  assign compressDataVec_hitReq_7_67 = _GEN_56;
  wire         compressDataVec_hitReq_7_99;
  assign compressDataVec_hitReq_7_99 = _GEN_56;
  wire         _GEN_57 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3;
  wire         compressDataVec_hitReq_8_3;
  assign compressDataVec_hitReq_8_3 = _GEN_57;
  wire         compressDataVec_hitReq_8_67;
  assign compressDataVec_hitReq_8_67 = _GEN_57;
  wire         _GEN_58 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3;
  wire         compressDataVec_hitReq_9_3;
  assign compressDataVec_hitReq_9_3 = _GEN_58;
  wire         compressDataVec_hitReq_9_67;
  assign compressDataVec_hitReq_9_67 = _GEN_58;
  wire         _GEN_59 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3;
  wire         compressDataVec_hitReq_10_3;
  assign compressDataVec_hitReq_10_3 = _GEN_59;
  wire         compressDataVec_hitReq_10_67;
  assign compressDataVec_hitReq_10_67 = _GEN_59;
  wire         _GEN_60 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3;
  wire         compressDataVec_hitReq_11_3;
  assign compressDataVec_hitReq_11_3 = _GEN_60;
  wire         compressDataVec_hitReq_11_67;
  assign compressDataVec_hitReq_11_67 = _GEN_60;
  wire         _GEN_61 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3;
  wire         compressDataVec_hitReq_12_3;
  assign compressDataVec_hitReq_12_3 = _GEN_61;
  wire         compressDataVec_hitReq_12_67;
  assign compressDataVec_hitReq_12_67 = _GEN_61;
  wire         _GEN_62 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3;
  wire         compressDataVec_hitReq_13_3;
  assign compressDataVec_hitReq_13_3 = _GEN_62;
  wire         compressDataVec_hitReq_13_67;
  assign compressDataVec_hitReq_13_67 = _GEN_62;
  wire         _GEN_63 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3;
  wire         compressDataVec_hitReq_14_3;
  assign compressDataVec_hitReq_14_3 = _GEN_63;
  wire         compressDataVec_hitReq_14_67;
  assign compressDataVec_hitReq_14_67 = _GEN_63;
  wire         _GEN_64 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3;
  wire         compressDataVec_hitReq_15_3;
  assign compressDataVec_hitReq_15_3 = _GEN_64;
  wire         compressDataVec_hitReq_15_67;
  assign compressDataVec_hitReq_15_67 = _GEN_64;
  wire         compressDataVec_hitReq_16_3 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3;
  wire         compressDataVec_hitReq_17_3 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3;
  wire         compressDataVec_hitReq_18_3 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3;
  wire         compressDataVec_hitReq_19_3 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3;
  wire         compressDataVec_hitReq_20_3 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3;
  wire         compressDataVec_hitReq_21_3 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3;
  wire         compressDataVec_hitReq_22_3 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3;
  wire         compressDataVec_hitReq_23_3 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3;
  wire         compressDataVec_hitReq_24_3 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3;
  wire         compressDataVec_hitReq_25_3 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3;
  wire         compressDataVec_hitReq_26_3 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3;
  wire         compressDataVec_hitReq_27_3 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3;
  wire         compressDataVec_hitReq_28_3 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3;
  wire         compressDataVec_hitReq_29_3 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3;
  wire         compressDataVec_hitReq_30_3 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3;
  wire         compressDataVec_hitReq_31_3 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3;
  wire [7:0]   compressDataVec_selectReqData_3 =
    (compressDataVec_hitReq_0_3 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_3 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_3 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_3 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_3 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_3 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_3 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_3 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_3 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_3 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_3 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_3 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_3 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_3 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_3 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_3 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_3 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_3 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_3 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_3 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_3 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_3 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_3 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_3 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_3 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_3 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_3 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_3 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_3 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_3 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_3 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_3 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_3;
  assign compressDataVec_useTail_3 = |(tailCount[4:2]);
  wire         _GEN_65 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h4;
  wire         compressDataVec_hitReq_0_4;
  assign compressDataVec_hitReq_0_4 = _GEN_65;
  wire         compressDataVec_hitReq_0_68;
  assign compressDataVec_hitReq_0_68 = _GEN_65;
  wire         compressDataVec_hitReq_0_100;
  assign compressDataVec_hitReq_0_100 = _GEN_65;
  wire         _GEN_66 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h4;
  wire         compressDataVec_hitReq_1_4;
  assign compressDataVec_hitReq_1_4 = _GEN_66;
  wire         compressDataVec_hitReq_1_68;
  assign compressDataVec_hitReq_1_68 = _GEN_66;
  wire         compressDataVec_hitReq_1_100;
  assign compressDataVec_hitReq_1_100 = _GEN_66;
  wire         _GEN_67 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h4;
  wire         compressDataVec_hitReq_2_4;
  assign compressDataVec_hitReq_2_4 = _GEN_67;
  wire         compressDataVec_hitReq_2_68;
  assign compressDataVec_hitReq_2_68 = _GEN_67;
  wire         compressDataVec_hitReq_2_100;
  assign compressDataVec_hitReq_2_100 = _GEN_67;
  wire         _GEN_68 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h4;
  wire         compressDataVec_hitReq_3_4;
  assign compressDataVec_hitReq_3_4 = _GEN_68;
  wire         compressDataVec_hitReq_3_68;
  assign compressDataVec_hitReq_3_68 = _GEN_68;
  wire         compressDataVec_hitReq_3_100;
  assign compressDataVec_hitReq_3_100 = _GEN_68;
  wire         _GEN_69 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h4;
  wire         compressDataVec_hitReq_4_4;
  assign compressDataVec_hitReq_4_4 = _GEN_69;
  wire         compressDataVec_hitReq_4_68;
  assign compressDataVec_hitReq_4_68 = _GEN_69;
  wire         compressDataVec_hitReq_4_100;
  assign compressDataVec_hitReq_4_100 = _GEN_69;
  wire         _GEN_70 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h4;
  wire         compressDataVec_hitReq_5_4;
  assign compressDataVec_hitReq_5_4 = _GEN_70;
  wire         compressDataVec_hitReq_5_68;
  assign compressDataVec_hitReq_5_68 = _GEN_70;
  wire         compressDataVec_hitReq_5_100;
  assign compressDataVec_hitReq_5_100 = _GEN_70;
  wire         _GEN_71 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h4;
  wire         compressDataVec_hitReq_6_4;
  assign compressDataVec_hitReq_6_4 = _GEN_71;
  wire         compressDataVec_hitReq_6_68;
  assign compressDataVec_hitReq_6_68 = _GEN_71;
  wire         compressDataVec_hitReq_6_100;
  assign compressDataVec_hitReq_6_100 = _GEN_71;
  wire         _GEN_72 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h4;
  wire         compressDataVec_hitReq_7_4;
  assign compressDataVec_hitReq_7_4 = _GEN_72;
  wire         compressDataVec_hitReq_7_68;
  assign compressDataVec_hitReq_7_68 = _GEN_72;
  wire         compressDataVec_hitReq_7_100;
  assign compressDataVec_hitReq_7_100 = _GEN_72;
  wire         _GEN_73 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h4;
  wire         compressDataVec_hitReq_8_4;
  assign compressDataVec_hitReq_8_4 = _GEN_73;
  wire         compressDataVec_hitReq_8_68;
  assign compressDataVec_hitReq_8_68 = _GEN_73;
  wire         _GEN_74 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h4;
  wire         compressDataVec_hitReq_9_4;
  assign compressDataVec_hitReq_9_4 = _GEN_74;
  wire         compressDataVec_hitReq_9_68;
  assign compressDataVec_hitReq_9_68 = _GEN_74;
  wire         _GEN_75 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h4;
  wire         compressDataVec_hitReq_10_4;
  assign compressDataVec_hitReq_10_4 = _GEN_75;
  wire         compressDataVec_hitReq_10_68;
  assign compressDataVec_hitReq_10_68 = _GEN_75;
  wire         _GEN_76 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h4;
  wire         compressDataVec_hitReq_11_4;
  assign compressDataVec_hitReq_11_4 = _GEN_76;
  wire         compressDataVec_hitReq_11_68;
  assign compressDataVec_hitReq_11_68 = _GEN_76;
  wire         _GEN_77 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h4;
  wire         compressDataVec_hitReq_12_4;
  assign compressDataVec_hitReq_12_4 = _GEN_77;
  wire         compressDataVec_hitReq_12_68;
  assign compressDataVec_hitReq_12_68 = _GEN_77;
  wire         _GEN_78 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h4;
  wire         compressDataVec_hitReq_13_4;
  assign compressDataVec_hitReq_13_4 = _GEN_78;
  wire         compressDataVec_hitReq_13_68;
  assign compressDataVec_hitReq_13_68 = _GEN_78;
  wire         _GEN_79 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h4;
  wire         compressDataVec_hitReq_14_4;
  assign compressDataVec_hitReq_14_4 = _GEN_79;
  wire         compressDataVec_hitReq_14_68;
  assign compressDataVec_hitReq_14_68 = _GEN_79;
  wire         _GEN_80 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h4;
  wire         compressDataVec_hitReq_15_4;
  assign compressDataVec_hitReq_15_4 = _GEN_80;
  wire         compressDataVec_hitReq_15_68;
  assign compressDataVec_hitReq_15_68 = _GEN_80;
  wire         compressDataVec_hitReq_16_4 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h4;
  wire         compressDataVec_hitReq_17_4 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h4;
  wire         compressDataVec_hitReq_18_4 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h4;
  wire         compressDataVec_hitReq_19_4 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h4;
  wire         compressDataVec_hitReq_20_4 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h4;
  wire         compressDataVec_hitReq_21_4 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h4;
  wire         compressDataVec_hitReq_22_4 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h4;
  wire         compressDataVec_hitReq_23_4 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h4;
  wire         compressDataVec_hitReq_24_4 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h4;
  wire         compressDataVec_hitReq_25_4 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h4;
  wire         compressDataVec_hitReq_26_4 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h4;
  wire         compressDataVec_hitReq_27_4 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h4;
  wire         compressDataVec_hitReq_28_4 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h4;
  wire         compressDataVec_hitReq_29_4 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h4;
  wire         compressDataVec_hitReq_30_4 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h4;
  wire         compressDataVec_hitReq_31_4 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h4;
  wire [7:0]   compressDataVec_selectReqData_4 =
    (compressDataVec_hitReq_0_4 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_4 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_4 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_4 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_4 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_4 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_4 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_4 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_4 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_4 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_4 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_4 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_4 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_4 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_4 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_4 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_4 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_4 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_4 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_4 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_4 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_4 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_4 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_4 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_4 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_4 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_4 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_4 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_4 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_4 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_4 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_4 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_81 = tailCount > 5'h4;
  wire         compressDataVec_useTail_4;
  assign compressDataVec_useTail_4 = _GEN_81;
  wire         compressDataVec_useTail_36;
  assign compressDataVec_useTail_36 = _GEN_81;
  wire         compressDataVec_useTail_52;
  assign compressDataVec_useTail_52 = _GEN_81;
  wire         _GEN_82 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h5;
  wire         compressDataVec_hitReq_0_5;
  assign compressDataVec_hitReq_0_5 = _GEN_82;
  wire         compressDataVec_hitReq_0_69;
  assign compressDataVec_hitReq_0_69 = _GEN_82;
  wire         compressDataVec_hitReq_0_101;
  assign compressDataVec_hitReq_0_101 = _GEN_82;
  wire         _GEN_83 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h5;
  wire         compressDataVec_hitReq_1_5;
  assign compressDataVec_hitReq_1_5 = _GEN_83;
  wire         compressDataVec_hitReq_1_69;
  assign compressDataVec_hitReq_1_69 = _GEN_83;
  wire         compressDataVec_hitReq_1_101;
  assign compressDataVec_hitReq_1_101 = _GEN_83;
  wire         _GEN_84 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h5;
  wire         compressDataVec_hitReq_2_5;
  assign compressDataVec_hitReq_2_5 = _GEN_84;
  wire         compressDataVec_hitReq_2_69;
  assign compressDataVec_hitReq_2_69 = _GEN_84;
  wire         compressDataVec_hitReq_2_101;
  assign compressDataVec_hitReq_2_101 = _GEN_84;
  wire         _GEN_85 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h5;
  wire         compressDataVec_hitReq_3_5;
  assign compressDataVec_hitReq_3_5 = _GEN_85;
  wire         compressDataVec_hitReq_3_69;
  assign compressDataVec_hitReq_3_69 = _GEN_85;
  wire         compressDataVec_hitReq_3_101;
  assign compressDataVec_hitReq_3_101 = _GEN_85;
  wire         _GEN_86 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h5;
  wire         compressDataVec_hitReq_4_5;
  assign compressDataVec_hitReq_4_5 = _GEN_86;
  wire         compressDataVec_hitReq_4_69;
  assign compressDataVec_hitReq_4_69 = _GEN_86;
  wire         compressDataVec_hitReq_4_101;
  assign compressDataVec_hitReq_4_101 = _GEN_86;
  wire         _GEN_87 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h5;
  wire         compressDataVec_hitReq_5_5;
  assign compressDataVec_hitReq_5_5 = _GEN_87;
  wire         compressDataVec_hitReq_5_69;
  assign compressDataVec_hitReq_5_69 = _GEN_87;
  wire         compressDataVec_hitReq_5_101;
  assign compressDataVec_hitReq_5_101 = _GEN_87;
  wire         _GEN_88 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h5;
  wire         compressDataVec_hitReq_6_5;
  assign compressDataVec_hitReq_6_5 = _GEN_88;
  wire         compressDataVec_hitReq_6_69;
  assign compressDataVec_hitReq_6_69 = _GEN_88;
  wire         compressDataVec_hitReq_6_101;
  assign compressDataVec_hitReq_6_101 = _GEN_88;
  wire         _GEN_89 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h5;
  wire         compressDataVec_hitReq_7_5;
  assign compressDataVec_hitReq_7_5 = _GEN_89;
  wire         compressDataVec_hitReq_7_69;
  assign compressDataVec_hitReq_7_69 = _GEN_89;
  wire         compressDataVec_hitReq_7_101;
  assign compressDataVec_hitReq_7_101 = _GEN_89;
  wire         _GEN_90 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h5;
  wire         compressDataVec_hitReq_8_5;
  assign compressDataVec_hitReq_8_5 = _GEN_90;
  wire         compressDataVec_hitReq_8_69;
  assign compressDataVec_hitReq_8_69 = _GEN_90;
  wire         _GEN_91 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h5;
  wire         compressDataVec_hitReq_9_5;
  assign compressDataVec_hitReq_9_5 = _GEN_91;
  wire         compressDataVec_hitReq_9_69;
  assign compressDataVec_hitReq_9_69 = _GEN_91;
  wire         _GEN_92 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h5;
  wire         compressDataVec_hitReq_10_5;
  assign compressDataVec_hitReq_10_5 = _GEN_92;
  wire         compressDataVec_hitReq_10_69;
  assign compressDataVec_hitReq_10_69 = _GEN_92;
  wire         _GEN_93 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h5;
  wire         compressDataVec_hitReq_11_5;
  assign compressDataVec_hitReq_11_5 = _GEN_93;
  wire         compressDataVec_hitReq_11_69;
  assign compressDataVec_hitReq_11_69 = _GEN_93;
  wire         _GEN_94 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h5;
  wire         compressDataVec_hitReq_12_5;
  assign compressDataVec_hitReq_12_5 = _GEN_94;
  wire         compressDataVec_hitReq_12_69;
  assign compressDataVec_hitReq_12_69 = _GEN_94;
  wire         _GEN_95 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h5;
  wire         compressDataVec_hitReq_13_5;
  assign compressDataVec_hitReq_13_5 = _GEN_95;
  wire         compressDataVec_hitReq_13_69;
  assign compressDataVec_hitReq_13_69 = _GEN_95;
  wire         _GEN_96 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h5;
  wire         compressDataVec_hitReq_14_5;
  assign compressDataVec_hitReq_14_5 = _GEN_96;
  wire         compressDataVec_hitReq_14_69;
  assign compressDataVec_hitReq_14_69 = _GEN_96;
  wire         _GEN_97 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h5;
  wire         compressDataVec_hitReq_15_5;
  assign compressDataVec_hitReq_15_5 = _GEN_97;
  wire         compressDataVec_hitReq_15_69;
  assign compressDataVec_hitReq_15_69 = _GEN_97;
  wire         compressDataVec_hitReq_16_5 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h5;
  wire         compressDataVec_hitReq_17_5 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h5;
  wire         compressDataVec_hitReq_18_5 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h5;
  wire         compressDataVec_hitReq_19_5 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h5;
  wire         compressDataVec_hitReq_20_5 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h5;
  wire         compressDataVec_hitReq_21_5 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h5;
  wire         compressDataVec_hitReq_22_5 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h5;
  wire         compressDataVec_hitReq_23_5 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h5;
  wire         compressDataVec_hitReq_24_5 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h5;
  wire         compressDataVec_hitReq_25_5 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h5;
  wire         compressDataVec_hitReq_26_5 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h5;
  wire         compressDataVec_hitReq_27_5 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h5;
  wire         compressDataVec_hitReq_28_5 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h5;
  wire         compressDataVec_hitReq_29_5 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h5;
  wire         compressDataVec_hitReq_30_5 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h5;
  wire         compressDataVec_hitReq_31_5 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h5;
  wire [7:0]   compressDataVec_selectReqData_5 =
    (compressDataVec_hitReq_0_5 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_5 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_5 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_5 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_5 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_5 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_5 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_5 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_5 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_5 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_5 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_5 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_5 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_5 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_5 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_5 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_5 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_5 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_5 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_5 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_5 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_5 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_5 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_5 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_5 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_5 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_5 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_5 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_5 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_5 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_5 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_5 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_98 = tailCount > 5'h5;
  wire         compressDataVec_useTail_5;
  assign compressDataVec_useTail_5 = _GEN_98;
  wire         compressDataVec_useTail_37;
  assign compressDataVec_useTail_37 = _GEN_98;
  wire         compressDataVec_useTail_53;
  assign compressDataVec_useTail_53 = _GEN_98;
  wire         _GEN_99 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h6;
  wire         compressDataVec_hitReq_0_6;
  assign compressDataVec_hitReq_0_6 = _GEN_99;
  wire         compressDataVec_hitReq_0_70;
  assign compressDataVec_hitReq_0_70 = _GEN_99;
  wire         compressDataVec_hitReq_0_102;
  assign compressDataVec_hitReq_0_102 = _GEN_99;
  wire         _GEN_100 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h6;
  wire         compressDataVec_hitReq_1_6;
  assign compressDataVec_hitReq_1_6 = _GEN_100;
  wire         compressDataVec_hitReq_1_70;
  assign compressDataVec_hitReq_1_70 = _GEN_100;
  wire         compressDataVec_hitReq_1_102;
  assign compressDataVec_hitReq_1_102 = _GEN_100;
  wire         _GEN_101 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h6;
  wire         compressDataVec_hitReq_2_6;
  assign compressDataVec_hitReq_2_6 = _GEN_101;
  wire         compressDataVec_hitReq_2_70;
  assign compressDataVec_hitReq_2_70 = _GEN_101;
  wire         compressDataVec_hitReq_2_102;
  assign compressDataVec_hitReq_2_102 = _GEN_101;
  wire         _GEN_102 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h6;
  wire         compressDataVec_hitReq_3_6;
  assign compressDataVec_hitReq_3_6 = _GEN_102;
  wire         compressDataVec_hitReq_3_70;
  assign compressDataVec_hitReq_3_70 = _GEN_102;
  wire         compressDataVec_hitReq_3_102;
  assign compressDataVec_hitReq_3_102 = _GEN_102;
  wire         _GEN_103 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h6;
  wire         compressDataVec_hitReq_4_6;
  assign compressDataVec_hitReq_4_6 = _GEN_103;
  wire         compressDataVec_hitReq_4_70;
  assign compressDataVec_hitReq_4_70 = _GEN_103;
  wire         compressDataVec_hitReq_4_102;
  assign compressDataVec_hitReq_4_102 = _GEN_103;
  wire         _GEN_104 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h6;
  wire         compressDataVec_hitReq_5_6;
  assign compressDataVec_hitReq_5_6 = _GEN_104;
  wire         compressDataVec_hitReq_5_70;
  assign compressDataVec_hitReq_5_70 = _GEN_104;
  wire         compressDataVec_hitReq_5_102;
  assign compressDataVec_hitReq_5_102 = _GEN_104;
  wire         _GEN_105 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h6;
  wire         compressDataVec_hitReq_6_6;
  assign compressDataVec_hitReq_6_6 = _GEN_105;
  wire         compressDataVec_hitReq_6_70;
  assign compressDataVec_hitReq_6_70 = _GEN_105;
  wire         compressDataVec_hitReq_6_102;
  assign compressDataVec_hitReq_6_102 = _GEN_105;
  wire         _GEN_106 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h6;
  wire         compressDataVec_hitReq_7_6;
  assign compressDataVec_hitReq_7_6 = _GEN_106;
  wire         compressDataVec_hitReq_7_70;
  assign compressDataVec_hitReq_7_70 = _GEN_106;
  wire         compressDataVec_hitReq_7_102;
  assign compressDataVec_hitReq_7_102 = _GEN_106;
  wire         _GEN_107 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h6;
  wire         compressDataVec_hitReq_8_6;
  assign compressDataVec_hitReq_8_6 = _GEN_107;
  wire         compressDataVec_hitReq_8_70;
  assign compressDataVec_hitReq_8_70 = _GEN_107;
  wire         _GEN_108 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h6;
  wire         compressDataVec_hitReq_9_6;
  assign compressDataVec_hitReq_9_6 = _GEN_108;
  wire         compressDataVec_hitReq_9_70;
  assign compressDataVec_hitReq_9_70 = _GEN_108;
  wire         _GEN_109 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h6;
  wire         compressDataVec_hitReq_10_6;
  assign compressDataVec_hitReq_10_6 = _GEN_109;
  wire         compressDataVec_hitReq_10_70;
  assign compressDataVec_hitReq_10_70 = _GEN_109;
  wire         _GEN_110 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h6;
  wire         compressDataVec_hitReq_11_6;
  assign compressDataVec_hitReq_11_6 = _GEN_110;
  wire         compressDataVec_hitReq_11_70;
  assign compressDataVec_hitReq_11_70 = _GEN_110;
  wire         _GEN_111 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h6;
  wire         compressDataVec_hitReq_12_6;
  assign compressDataVec_hitReq_12_6 = _GEN_111;
  wire         compressDataVec_hitReq_12_70;
  assign compressDataVec_hitReq_12_70 = _GEN_111;
  wire         _GEN_112 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h6;
  wire         compressDataVec_hitReq_13_6;
  assign compressDataVec_hitReq_13_6 = _GEN_112;
  wire         compressDataVec_hitReq_13_70;
  assign compressDataVec_hitReq_13_70 = _GEN_112;
  wire         _GEN_113 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h6;
  wire         compressDataVec_hitReq_14_6;
  assign compressDataVec_hitReq_14_6 = _GEN_113;
  wire         compressDataVec_hitReq_14_70;
  assign compressDataVec_hitReq_14_70 = _GEN_113;
  wire         _GEN_114 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h6;
  wire         compressDataVec_hitReq_15_6;
  assign compressDataVec_hitReq_15_6 = _GEN_114;
  wire         compressDataVec_hitReq_15_70;
  assign compressDataVec_hitReq_15_70 = _GEN_114;
  wire         compressDataVec_hitReq_16_6 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h6;
  wire         compressDataVec_hitReq_17_6 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h6;
  wire         compressDataVec_hitReq_18_6 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h6;
  wire         compressDataVec_hitReq_19_6 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h6;
  wire         compressDataVec_hitReq_20_6 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h6;
  wire         compressDataVec_hitReq_21_6 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h6;
  wire         compressDataVec_hitReq_22_6 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h6;
  wire         compressDataVec_hitReq_23_6 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h6;
  wire         compressDataVec_hitReq_24_6 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h6;
  wire         compressDataVec_hitReq_25_6 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h6;
  wire         compressDataVec_hitReq_26_6 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h6;
  wire         compressDataVec_hitReq_27_6 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h6;
  wire         compressDataVec_hitReq_28_6 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h6;
  wire         compressDataVec_hitReq_29_6 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h6;
  wire         compressDataVec_hitReq_30_6 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h6;
  wire         compressDataVec_hitReq_31_6 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h6;
  wire [7:0]   compressDataVec_selectReqData_6 =
    (compressDataVec_hitReq_0_6 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_6 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_6 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_6 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_6 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_6 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_6 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_6 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_6 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_6 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_6 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_6 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_6 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_6 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_6 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_6 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_6 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_6 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_6 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_6 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_6 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_6 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_6 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_6 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_6 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_6 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_6 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_6 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_6 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_6 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_6 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_6 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_115 = tailCount > 5'h6;
  wire         compressDataVec_useTail_6;
  assign compressDataVec_useTail_6 = _GEN_115;
  wire         compressDataVec_useTail_38;
  assign compressDataVec_useTail_38 = _GEN_115;
  wire         compressDataVec_useTail_54;
  assign compressDataVec_useTail_54 = _GEN_115;
  wire         _GEN_116 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h7;
  wire         compressDataVec_hitReq_0_7;
  assign compressDataVec_hitReq_0_7 = _GEN_116;
  wire         compressDataVec_hitReq_0_71;
  assign compressDataVec_hitReq_0_71 = _GEN_116;
  wire         compressDataVec_hitReq_0_103;
  assign compressDataVec_hitReq_0_103 = _GEN_116;
  wire         _GEN_117 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h7;
  wire         compressDataVec_hitReq_1_7;
  assign compressDataVec_hitReq_1_7 = _GEN_117;
  wire         compressDataVec_hitReq_1_71;
  assign compressDataVec_hitReq_1_71 = _GEN_117;
  wire         compressDataVec_hitReq_1_103;
  assign compressDataVec_hitReq_1_103 = _GEN_117;
  wire         _GEN_118 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h7;
  wire         compressDataVec_hitReq_2_7;
  assign compressDataVec_hitReq_2_7 = _GEN_118;
  wire         compressDataVec_hitReq_2_71;
  assign compressDataVec_hitReq_2_71 = _GEN_118;
  wire         compressDataVec_hitReq_2_103;
  assign compressDataVec_hitReq_2_103 = _GEN_118;
  wire         _GEN_119 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h7;
  wire         compressDataVec_hitReq_3_7;
  assign compressDataVec_hitReq_3_7 = _GEN_119;
  wire         compressDataVec_hitReq_3_71;
  assign compressDataVec_hitReq_3_71 = _GEN_119;
  wire         compressDataVec_hitReq_3_103;
  assign compressDataVec_hitReq_3_103 = _GEN_119;
  wire         _GEN_120 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h7;
  wire         compressDataVec_hitReq_4_7;
  assign compressDataVec_hitReq_4_7 = _GEN_120;
  wire         compressDataVec_hitReq_4_71;
  assign compressDataVec_hitReq_4_71 = _GEN_120;
  wire         compressDataVec_hitReq_4_103;
  assign compressDataVec_hitReq_4_103 = _GEN_120;
  wire         _GEN_121 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h7;
  wire         compressDataVec_hitReq_5_7;
  assign compressDataVec_hitReq_5_7 = _GEN_121;
  wire         compressDataVec_hitReq_5_71;
  assign compressDataVec_hitReq_5_71 = _GEN_121;
  wire         compressDataVec_hitReq_5_103;
  assign compressDataVec_hitReq_5_103 = _GEN_121;
  wire         _GEN_122 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h7;
  wire         compressDataVec_hitReq_6_7;
  assign compressDataVec_hitReq_6_7 = _GEN_122;
  wire         compressDataVec_hitReq_6_71;
  assign compressDataVec_hitReq_6_71 = _GEN_122;
  wire         compressDataVec_hitReq_6_103;
  assign compressDataVec_hitReq_6_103 = _GEN_122;
  wire         _GEN_123 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h7;
  wire         compressDataVec_hitReq_7_7;
  assign compressDataVec_hitReq_7_7 = _GEN_123;
  wire         compressDataVec_hitReq_7_71;
  assign compressDataVec_hitReq_7_71 = _GEN_123;
  wire         compressDataVec_hitReq_7_103;
  assign compressDataVec_hitReq_7_103 = _GEN_123;
  wire         _GEN_124 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h7;
  wire         compressDataVec_hitReq_8_7;
  assign compressDataVec_hitReq_8_7 = _GEN_124;
  wire         compressDataVec_hitReq_8_71;
  assign compressDataVec_hitReq_8_71 = _GEN_124;
  wire         _GEN_125 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h7;
  wire         compressDataVec_hitReq_9_7;
  assign compressDataVec_hitReq_9_7 = _GEN_125;
  wire         compressDataVec_hitReq_9_71;
  assign compressDataVec_hitReq_9_71 = _GEN_125;
  wire         _GEN_126 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h7;
  wire         compressDataVec_hitReq_10_7;
  assign compressDataVec_hitReq_10_7 = _GEN_126;
  wire         compressDataVec_hitReq_10_71;
  assign compressDataVec_hitReq_10_71 = _GEN_126;
  wire         _GEN_127 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h7;
  wire         compressDataVec_hitReq_11_7;
  assign compressDataVec_hitReq_11_7 = _GEN_127;
  wire         compressDataVec_hitReq_11_71;
  assign compressDataVec_hitReq_11_71 = _GEN_127;
  wire         _GEN_128 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h7;
  wire         compressDataVec_hitReq_12_7;
  assign compressDataVec_hitReq_12_7 = _GEN_128;
  wire         compressDataVec_hitReq_12_71;
  assign compressDataVec_hitReq_12_71 = _GEN_128;
  wire         _GEN_129 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h7;
  wire         compressDataVec_hitReq_13_7;
  assign compressDataVec_hitReq_13_7 = _GEN_129;
  wire         compressDataVec_hitReq_13_71;
  assign compressDataVec_hitReq_13_71 = _GEN_129;
  wire         _GEN_130 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h7;
  wire         compressDataVec_hitReq_14_7;
  assign compressDataVec_hitReq_14_7 = _GEN_130;
  wire         compressDataVec_hitReq_14_71;
  assign compressDataVec_hitReq_14_71 = _GEN_130;
  wire         _GEN_131 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h7;
  wire         compressDataVec_hitReq_15_7;
  assign compressDataVec_hitReq_15_7 = _GEN_131;
  wire         compressDataVec_hitReq_15_71;
  assign compressDataVec_hitReq_15_71 = _GEN_131;
  wire         compressDataVec_hitReq_16_7 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h7;
  wire         compressDataVec_hitReq_17_7 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h7;
  wire         compressDataVec_hitReq_18_7 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h7;
  wire         compressDataVec_hitReq_19_7 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h7;
  wire         compressDataVec_hitReq_20_7 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h7;
  wire         compressDataVec_hitReq_21_7 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h7;
  wire         compressDataVec_hitReq_22_7 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h7;
  wire         compressDataVec_hitReq_23_7 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h7;
  wire         compressDataVec_hitReq_24_7 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h7;
  wire         compressDataVec_hitReq_25_7 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h7;
  wire         compressDataVec_hitReq_26_7 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h7;
  wire         compressDataVec_hitReq_27_7 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h7;
  wire         compressDataVec_hitReq_28_7 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h7;
  wire         compressDataVec_hitReq_29_7 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h7;
  wire         compressDataVec_hitReq_30_7 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h7;
  wire         compressDataVec_hitReq_31_7 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h7;
  wire [7:0]   compressDataVec_selectReqData_7 =
    (compressDataVec_hitReq_0_7 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_7 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_7 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_7 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_7 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_7 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_7 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_7 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_7 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_7 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_7 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_7 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_7 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_7 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_7 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_7 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_7 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_7 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_7 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_7 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_7 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_7 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_7 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_7 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_7 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_7 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_7 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_7 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_7 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_7 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_7 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_7 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_7;
  assign compressDataVec_useTail_7 = |(tailCount[4:3]);
  wire         _GEN_132 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h8;
  wire         compressDataVec_hitReq_0_8;
  assign compressDataVec_hitReq_0_8 = _GEN_132;
  wire         compressDataVec_hitReq_0_72;
  assign compressDataVec_hitReq_0_72 = _GEN_132;
  wire         compressDataVec_hitReq_0_104;
  assign compressDataVec_hitReq_0_104 = _GEN_132;
  wire         _GEN_133 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h8;
  wire         compressDataVec_hitReq_1_8;
  assign compressDataVec_hitReq_1_8 = _GEN_133;
  wire         compressDataVec_hitReq_1_72;
  assign compressDataVec_hitReq_1_72 = _GEN_133;
  wire         compressDataVec_hitReq_1_104;
  assign compressDataVec_hitReq_1_104 = _GEN_133;
  wire         _GEN_134 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h8;
  wire         compressDataVec_hitReq_2_8;
  assign compressDataVec_hitReq_2_8 = _GEN_134;
  wire         compressDataVec_hitReq_2_72;
  assign compressDataVec_hitReq_2_72 = _GEN_134;
  wire         compressDataVec_hitReq_2_104;
  assign compressDataVec_hitReq_2_104 = _GEN_134;
  wire         _GEN_135 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h8;
  wire         compressDataVec_hitReq_3_8;
  assign compressDataVec_hitReq_3_8 = _GEN_135;
  wire         compressDataVec_hitReq_3_72;
  assign compressDataVec_hitReq_3_72 = _GEN_135;
  wire         compressDataVec_hitReq_3_104;
  assign compressDataVec_hitReq_3_104 = _GEN_135;
  wire         _GEN_136 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h8;
  wire         compressDataVec_hitReq_4_8;
  assign compressDataVec_hitReq_4_8 = _GEN_136;
  wire         compressDataVec_hitReq_4_72;
  assign compressDataVec_hitReq_4_72 = _GEN_136;
  wire         compressDataVec_hitReq_4_104;
  assign compressDataVec_hitReq_4_104 = _GEN_136;
  wire         _GEN_137 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h8;
  wire         compressDataVec_hitReq_5_8;
  assign compressDataVec_hitReq_5_8 = _GEN_137;
  wire         compressDataVec_hitReq_5_72;
  assign compressDataVec_hitReq_5_72 = _GEN_137;
  wire         compressDataVec_hitReq_5_104;
  assign compressDataVec_hitReq_5_104 = _GEN_137;
  wire         _GEN_138 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h8;
  wire         compressDataVec_hitReq_6_8;
  assign compressDataVec_hitReq_6_8 = _GEN_138;
  wire         compressDataVec_hitReq_6_72;
  assign compressDataVec_hitReq_6_72 = _GEN_138;
  wire         compressDataVec_hitReq_6_104;
  assign compressDataVec_hitReq_6_104 = _GEN_138;
  wire         _GEN_139 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h8;
  wire         compressDataVec_hitReq_7_8;
  assign compressDataVec_hitReq_7_8 = _GEN_139;
  wire         compressDataVec_hitReq_7_72;
  assign compressDataVec_hitReq_7_72 = _GEN_139;
  wire         compressDataVec_hitReq_7_104;
  assign compressDataVec_hitReq_7_104 = _GEN_139;
  wire         _GEN_140 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h8;
  wire         compressDataVec_hitReq_8_8;
  assign compressDataVec_hitReq_8_8 = _GEN_140;
  wire         compressDataVec_hitReq_8_72;
  assign compressDataVec_hitReq_8_72 = _GEN_140;
  wire         _GEN_141 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h8;
  wire         compressDataVec_hitReq_9_8;
  assign compressDataVec_hitReq_9_8 = _GEN_141;
  wire         compressDataVec_hitReq_9_72;
  assign compressDataVec_hitReq_9_72 = _GEN_141;
  wire         _GEN_142 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h8;
  wire         compressDataVec_hitReq_10_8;
  assign compressDataVec_hitReq_10_8 = _GEN_142;
  wire         compressDataVec_hitReq_10_72;
  assign compressDataVec_hitReq_10_72 = _GEN_142;
  wire         _GEN_143 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h8;
  wire         compressDataVec_hitReq_11_8;
  assign compressDataVec_hitReq_11_8 = _GEN_143;
  wire         compressDataVec_hitReq_11_72;
  assign compressDataVec_hitReq_11_72 = _GEN_143;
  wire         _GEN_144 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h8;
  wire         compressDataVec_hitReq_12_8;
  assign compressDataVec_hitReq_12_8 = _GEN_144;
  wire         compressDataVec_hitReq_12_72;
  assign compressDataVec_hitReq_12_72 = _GEN_144;
  wire         _GEN_145 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h8;
  wire         compressDataVec_hitReq_13_8;
  assign compressDataVec_hitReq_13_8 = _GEN_145;
  wire         compressDataVec_hitReq_13_72;
  assign compressDataVec_hitReq_13_72 = _GEN_145;
  wire         _GEN_146 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h8;
  wire         compressDataVec_hitReq_14_8;
  assign compressDataVec_hitReq_14_8 = _GEN_146;
  wire         compressDataVec_hitReq_14_72;
  assign compressDataVec_hitReq_14_72 = _GEN_146;
  wire         _GEN_147 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h8;
  wire         compressDataVec_hitReq_15_8;
  assign compressDataVec_hitReq_15_8 = _GEN_147;
  wire         compressDataVec_hitReq_15_72;
  assign compressDataVec_hitReq_15_72 = _GEN_147;
  wire         compressDataVec_hitReq_16_8 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h8;
  wire         compressDataVec_hitReq_17_8 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h8;
  wire         compressDataVec_hitReq_18_8 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h8;
  wire         compressDataVec_hitReq_19_8 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h8;
  wire         compressDataVec_hitReq_20_8 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h8;
  wire         compressDataVec_hitReq_21_8 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h8;
  wire         compressDataVec_hitReq_22_8 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h8;
  wire         compressDataVec_hitReq_23_8 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h8;
  wire         compressDataVec_hitReq_24_8 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h8;
  wire         compressDataVec_hitReq_25_8 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h8;
  wire         compressDataVec_hitReq_26_8 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h8;
  wire         compressDataVec_hitReq_27_8 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h8;
  wire         compressDataVec_hitReq_28_8 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h8;
  wire         compressDataVec_hitReq_29_8 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h8;
  wire         compressDataVec_hitReq_30_8 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h8;
  wire         compressDataVec_hitReq_31_8 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h8;
  wire [7:0]   compressDataVec_selectReqData_8 =
    (compressDataVec_hitReq_0_8 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_8 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_8 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_8 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_8 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_8 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_8 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_8 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_8 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_8 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_8 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_8 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_8 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_8 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_8 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_8 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_8 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_8 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_8 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_8 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_8 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_8 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_8 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_8 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_8 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_8 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_8 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_8 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_8 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_8 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_8 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_8 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_148 = tailCount > 5'h8;
  wire         compressDataVec_useTail_8;
  assign compressDataVec_useTail_8 = _GEN_148;
  wire         compressDataVec_useTail_40;
  assign compressDataVec_useTail_40 = _GEN_148;
  wire         _GEN_149 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h9;
  wire         compressDataVec_hitReq_0_9;
  assign compressDataVec_hitReq_0_9 = _GEN_149;
  wire         compressDataVec_hitReq_0_73;
  assign compressDataVec_hitReq_0_73 = _GEN_149;
  wire         compressDataVec_hitReq_0_105;
  assign compressDataVec_hitReq_0_105 = _GEN_149;
  wire         _GEN_150 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h9;
  wire         compressDataVec_hitReq_1_9;
  assign compressDataVec_hitReq_1_9 = _GEN_150;
  wire         compressDataVec_hitReq_1_73;
  assign compressDataVec_hitReq_1_73 = _GEN_150;
  wire         compressDataVec_hitReq_1_105;
  assign compressDataVec_hitReq_1_105 = _GEN_150;
  wire         _GEN_151 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h9;
  wire         compressDataVec_hitReq_2_9;
  assign compressDataVec_hitReq_2_9 = _GEN_151;
  wire         compressDataVec_hitReq_2_73;
  assign compressDataVec_hitReq_2_73 = _GEN_151;
  wire         compressDataVec_hitReq_2_105;
  assign compressDataVec_hitReq_2_105 = _GEN_151;
  wire         _GEN_152 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h9;
  wire         compressDataVec_hitReq_3_9;
  assign compressDataVec_hitReq_3_9 = _GEN_152;
  wire         compressDataVec_hitReq_3_73;
  assign compressDataVec_hitReq_3_73 = _GEN_152;
  wire         compressDataVec_hitReq_3_105;
  assign compressDataVec_hitReq_3_105 = _GEN_152;
  wire         _GEN_153 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h9;
  wire         compressDataVec_hitReq_4_9;
  assign compressDataVec_hitReq_4_9 = _GEN_153;
  wire         compressDataVec_hitReq_4_73;
  assign compressDataVec_hitReq_4_73 = _GEN_153;
  wire         compressDataVec_hitReq_4_105;
  assign compressDataVec_hitReq_4_105 = _GEN_153;
  wire         _GEN_154 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h9;
  wire         compressDataVec_hitReq_5_9;
  assign compressDataVec_hitReq_5_9 = _GEN_154;
  wire         compressDataVec_hitReq_5_73;
  assign compressDataVec_hitReq_5_73 = _GEN_154;
  wire         compressDataVec_hitReq_5_105;
  assign compressDataVec_hitReq_5_105 = _GEN_154;
  wire         _GEN_155 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h9;
  wire         compressDataVec_hitReq_6_9;
  assign compressDataVec_hitReq_6_9 = _GEN_155;
  wire         compressDataVec_hitReq_6_73;
  assign compressDataVec_hitReq_6_73 = _GEN_155;
  wire         compressDataVec_hitReq_6_105;
  assign compressDataVec_hitReq_6_105 = _GEN_155;
  wire         _GEN_156 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h9;
  wire         compressDataVec_hitReq_7_9;
  assign compressDataVec_hitReq_7_9 = _GEN_156;
  wire         compressDataVec_hitReq_7_73;
  assign compressDataVec_hitReq_7_73 = _GEN_156;
  wire         compressDataVec_hitReq_7_105;
  assign compressDataVec_hitReq_7_105 = _GEN_156;
  wire         _GEN_157 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h9;
  wire         compressDataVec_hitReq_8_9;
  assign compressDataVec_hitReq_8_9 = _GEN_157;
  wire         compressDataVec_hitReq_8_73;
  assign compressDataVec_hitReq_8_73 = _GEN_157;
  wire         _GEN_158 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h9;
  wire         compressDataVec_hitReq_9_9;
  assign compressDataVec_hitReq_9_9 = _GEN_158;
  wire         compressDataVec_hitReq_9_73;
  assign compressDataVec_hitReq_9_73 = _GEN_158;
  wire         _GEN_159 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h9;
  wire         compressDataVec_hitReq_10_9;
  assign compressDataVec_hitReq_10_9 = _GEN_159;
  wire         compressDataVec_hitReq_10_73;
  assign compressDataVec_hitReq_10_73 = _GEN_159;
  wire         _GEN_160 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h9;
  wire         compressDataVec_hitReq_11_9;
  assign compressDataVec_hitReq_11_9 = _GEN_160;
  wire         compressDataVec_hitReq_11_73;
  assign compressDataVec_hitReq_11_73 = _GEN_160;
  wire         _GEN_161 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h9;
  wire         compressDataVec_hitReq_12_9;
  assign compressDataVec_hitReq_12_9 = _GEN_161;
  wire         compressDataVec_hitReq_12_73;
  assign compressDataVec_hitReq_12_73 = _GEN_161;
  wire         _GEN_162 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h9;
  wire         compressDataVec_hitReq_13_9;
  assign compressDataVec_hitReq_13_9 = _GEN_162;
  wire         compressDataVec_hitReq_13_73;
  assign compressDataVec_hitReq_13_73 = _GEN_162;
  wire         _GEN_163 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h9;
  wire         compressDataVec_hitReq_14_9;
  assign compressDataVec_hitReq_14_9 = _GEN_163;
  wire         compressDataVec_hitReq_14_73;
  assign compressDataVec_hitReq_14_73 = _GEN_163;
  wire         _GEN_164 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h9;
  wire         compressDataVec_hitReq_15_9;
  assign compressDataVec_hitReq_15_9 = _GEN_164;
  wire         compressDataVec_hitReq_15_73;
  assign compressDataVec_hitReq_15_73 = _GEN_164;
  wire         compressDataVec_hitReq_16_9 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h9;
  wire         compressDataVec_hitReq_17_9 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h9;
  wire         compressDataVec_hitReq_18_9 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h9;
  wire         compressDataVec_hitReq_19_9 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h9;
  wire         compressDataVec_hitReq_20_9 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h9;
  wire         compressDataVec_hitReq_21_9 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h9;
  wire         compressDataVec_hitReq_22_9 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h9;
  wire         compressDataVec_hitReq_23_9 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h9;
  wire         compressDataVec_hitReq_24_9 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h9;
  wire         compressDataVec_hitReq_25_9 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h9;
  wire         compressDataVec_hitReq_26_9 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h9;
  wire         compressDataVec_hitReq_27_9 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h9;
  wire         compressDataVec_hitReq_28_9 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h9;
  wire         compressDataVec_hitReq_29_9 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h9;
  wire         compressDataVec_hitReq_30_9 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h9;
  wire         compressDataVec_hitReq_31_9 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h9;
  wire [7:0]   compressDataVec_selectReqData_9 =
    (compressDataVec_hitReq_0_9 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_9 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_9 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_9 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_9 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_9 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_9 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_9 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_9 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_9 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_9 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_9 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_9 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_9 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_9 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_9 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_9 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_9 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_9 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_9 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_9 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_9 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_9 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_9 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_9 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_9 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_9 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_9 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_9 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_9 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_9 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_9 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_165 = tailCount > 5'h9;
  wire         compressDataVec_useTail_9;
  assign compressDataVec_useTail_9 = _GEN_165;
  wire         compressDataVec_useTail_41;
  assign compressDataVec_useTail_41 = _GEN_165;
  wire         _GEN_166 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hA;
  wire         compressDataVec_hitReq_0_10;
  assign compressDataVec_hitReq_0_10 = _GEN_166;
  wire         compressDataVec_hitReq_0_74;
  assign compressDataVec_hitReq_0_74 = _GEN_166;
  wire         compressDataVec_hitReq_0_106;
  assign compressDataVec_hitReq_0_106 = _GEN_166;
  wire         _GEN_167 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hA;
  wire         compressDataVec_hitReq_1_10;
  assign compressDataVec_hitReq_1_10 = _GEN_167;
  wire         compressDataVec_hitReq_1_74;
  assign compressDataVec_hitReq_1_74 = _GEN_167;
  wire         compressDataVec_hitReq_1_106;
  assign compressDataVec_hitReq_1_106 = _GEN_167;
  wire         _GEN_168 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hA;
  wire         compressDataVec_hitReq_2_10;
  assign compressDataVec_hitReq_2_10 = _GEN_168;
  wire         compressDataVec_hitReq_2_74;
  assign compressDataVec_hitReq_2_74 = _GEN_168;
  wire         compressDataVec_hitReq_2_106;
  assign compressDataVec_hitReq_2_106 = _GEN_168;
  wire         _GEN_169 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hA;
  wire         compressDataVec_hitReq_3_10;
  assign compressDataVec_hitReq_3_10 = _GEN_169;
  wire         compressDataVec_hitReq_3_74;
  assign compressDataVec_hitReq_3_74 = _GEN_169;
  wire         compressDataVec_hitReq_3_106;
  assign compressDataVec_hitReq_3_106 = _GEN_169;
  wire         _GEN_170 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hA;
  wire         compressDataVec_hitReq_4_10;
  assign compressDataVec_hitReq_4_10 = _GEN_170;
  wire         compressDataVec_hitReq_4_74;
  assign compressDataVec_hitReq_4_74 = _GEN_170;
  wire         compressDataVec_hitReq_4_106;
  assign compressDataVec_hitReq_4_106 = _GEN_170;
  wire         _GEN_171 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hA;
  wire         compressDataVec_hitReq_5_10;
  assign compressDataVec_hitReq_5_10 = _GEN_171;
  wire         compressDataVec_hitReq_5_74;
  assign compressDataVec_hitReq_5_74 = _GEN_171;
  wire         compressDataVec_hitReq_5_106;
  assign compressDataVec_hitReq_5_106 = _GEN_171;
  wire         _GEN_172 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hA;
  wire         compressDataVec_hitReq_6_10;
  assign compressDataVec_hitReq_6_10 = _GEN_172;
  wire         compressDataVec_hitReq_6_74;
  assign compressDataVec_hitReq_6_74 = _GEN_172;
  wire         compressDataVec_hitReq_6_106;
  assign compressDataVec_hitReq_6_106 = _GEN_172;
  wire         _GEN_173 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hA;
  wire         compressDataVec_hitReq_7_10;
  assign compressDataVec_hitReq_7_10 = _GEN_173;
  wire         compressDataVec_hitReq_7_74;
  assign compressDataVec_hitReq_7_74 = _GEN_173;
  wire         compressDataVec_hitReq_7_106;
  assign compressDataVec_hitReq_7_106 = _GEN_173;
  wire         _GEN_174 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hA;
  wire         compressDataVec_hitReq_8_10;
  assign compressDataVec_hitReq_8_10 = _GEN_174;
  wire         compressDataVec_hitReq_8_74;
  assign compressDataVec_hitReq_8_74 = _GEN_174;
  wire         _GEN_175 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hA;
  wire         compressDataVec_hitReq_9_10;
  assign compressDataVec_hitReq_9_10 = _GEN_175;
  wire         compressDataVec_hitReq_9_74;
  assign compressDataVec_hitReq_9_74 = _GEN_175;
  wire         _GEN_176 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hA;
  wire         compressDataVec_hitReq_10_10;
  assign compressDataVec_hitReq_10_10 = _GEN_176;
  wire         compressDataVec_hitReq_10_74;
  assign compressDataVec_hitReq_10_74 = _GEN_176;
  wire         _GEN_177 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hA;
  wire         compressDataVec_hitReq_11_10;
  assign compressDataVec_hitReq_11_10 = _GEN_177;
  wire         compressDataVec_hitReq_11_74;
  assign compressDataVec_hitReq_11_74 = _GEN_177;
  wire         _GEN_178 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hA;
  wire         compressDataVec_hitReq_12_10;
  assign compressDataVec_hitReq_12_10 = _GEN_178;
  wire         compressDataVec_hitReq_12_74;
  assign compressDataVec_hitReq_12_74 = _GEN_178;
  wire         _GEN_179 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hA;
  wire         compressDataVec_hitReq_13_10;
  assign compressDataVec_hitReq_13_10 = _GEN_179;
  wire         compressDataVec_hitReq_13_74;
  assign compressDataVec_hitReq_13_74 = _GEN_179;
  wire         _GEN_180 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hA;
  wire         compressDataVec_hitReq_14_10;
  assign compressDataVec_hitReq_14_10 = _GEN_180;
  wire         compressDataVec_hitReq_14_74;
  assign compressDataVec_hitReq_14_74 = _GEN_180;
  wire         _GEN_181 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hA;
  wire         compressDataVec_hitReq_15_10;
  assign compressDataVec_hitReq_15_10 = _GEN_181;
  wire         compressDataVec_hitReq_15_74;
  assign compressDataVec_hitReq_15_74 = _GEN_181;
  wire         compressDataVec_hitReq_16_10 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hA;
  wire         compressDataVec_hitReq_17_10 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hA;
  wire         compressDataVec_hitReq_18_10 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hA;
  wire         compressDataVec_hitReq_19_10 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hA;
  wire         compressDataVec_hitReq_20_10 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hA;
  wire         compressDataVec_hitReq_21_10 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hA;
  wire         compressDataVec_hitReq_22_10 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hA;
  wire         compressDataVec_hitReq_23_10 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hA;
  wire         compressDataVec_hitReq_24_10 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hA;
  wire         compressDataVec_hitReq_25_10 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hA;
  wire         compressDataVec_hitReq_26_10 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hA;
  wire         compressDataVec_hitReq_27_10 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hA;
  wire         compressDataVec_hitReq_28_10 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hA;
  wire         compressDataVec_hitReq_29_10 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hA;
  wire         compressDataVec_hitReq_30_10 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hA;
  wire         compressDataVec_hitReq_31_10 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hA;
  wire [7:0]   compressDataVec_selectReqData_10 =
    (compressDataVec_hitReq_0_10 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_10 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_10 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_10 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_10 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_10 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_10 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_10 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_10 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_10 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_10 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_10 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_10 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_10 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_10 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_10 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_10 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_10 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_10 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_10 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_10 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_10 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_10 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_10 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_10 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_10 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_10 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_10 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_10 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_10 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_10 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_10 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_182 = tailCount > 5'hA;
  wire         compressDataVec_useTail_10;
  assign compressDataVec_useTail_10 = _GEN_182;
  wire         compressDataVec_useTail_42;
  assign compressDataVec_useTail_42 = _GEN_182;
  wire         _GEN_183 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hB;
  wire         compressDataVec_hitReq_0_11;
  assign compressDataVec_hitReq_0_11 = _GEN_183;
  wire         compressDataVec_hitReq_0_75;
  assign compressDataVec_hitReq_0_75 = _GEN_183;
  wire         compressDataVec_hitReq_0_107;
  assign compressDataVec_hitReq_0_107 = _GEN_183;
  wire         _GEN_184 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hB;
  wire         compressDataVec_hitReq_1_11;
  assign compressDataVec_hitReq_1_11 = _GEN_184;
  wire         compressDataVec_hitReq_1_75;
  assign compressDataVec_hitReq_1_75 = _GEN_184;
  wire         compressDataVec_hitReq_1_107;
  assign compressDataVec_hitReq_1_107 = _GEN_184;
  wire         _GEN_185 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hB;
  wire         compressDataVec_hitReq_2_11;
  assign compressDataVec_hitReq_2_11 = _GEN_185;
  wire         compressDataVec_hitReq_2_75;
  assign compressDataVec_hitReq_2_75 = _GEN_185;
  wire         compressDataVec_hitReq_2_107;
  assign compressDataVec_hitReq_2_107 = _GEN_185;
  wire         _GEN_186 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hB;
  wire         compressDataVec_hitReq_3_11;
  assign compressDataVec_hitReq_3_11 = _GEN_186;
  wire         compressDataVec_hitReq_3_75;
  assign compressDataVec_hitReq_3_75 = _GEN_186;
  wire         compressDataVec_hitReq_3_107;
  assign compressDataVec_hitReq_3_107 = _GEN_186;
  wire         _GEN_187 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hB;
  wire         compressDataVec_hitReq_4_11;
  assign compressDataVec_hitReq_4_11 = _GEN_187;
  wire         compressDataVec_hitReq_4_75;
  assign compressDataVec_hitReq_4_75 = _GEN_187;
  wire         compressDataVec_hitReq_4_107;
  assign compressDataVec_hitReq_4_107 = _GEN_187;
  wire         _GEN_188 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hB;
  wire         compressDataVec_hitReq_5_11;
  assign compressDataVec_hitReq_5_11 = _GEN_188;
  wire         compressDataVec_hitReq_5_75;
  assign compressDataVec_hitReq_5_75 = _GEN_188;
  wire         compressDataVec_hitReq_5_107;
  assign compressDataVec_hitReq_5_107 = _GEN_188;
  wire         _GEN_189 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hB;
  wire         compressDataVec_hitReq_6_11;
  assign compressDataVec_hitReq_6_11 = _GEN_189;
  wire         compressDataVec_hitReq_6_75;
  assign compressDataVec_hitReq_6_75 = _GEN_189;
  wire         compressDataVec_hitReq_6_107;
  assign compressDataVec_hitReq_6_107 = _GEN_189;
  wire         _GEN_190 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hB;
  wire         compressDataVec_hitReq_7_11;
  assign compressDataVec_hitReq_7_11 = _GEN_190;
  wire         compressDataVec_hitReq_7_75;
  assign compressDataVec_hitReq_7_75 = _GEN_190;
  wire         compressDataVec_hitReq_7_107;
  assign compressDataVec_hitReq_7_107 = _GEN_190;
  wire         _GEN_191 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hB;
  wire         compressDataVec_hitReq_8_11;
  assign compressDataVec_hitReq_8_11 = _GEN_191;
  wire         compressDataVec_hitReq_8_75;
  assign compressDataVec_hitReq_8_75 = _GEN_191;
  wire         _GEN_192 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hB;
  wire         compressDataVec_hitReq_9_11;
  assign compressDataVec_hitReq_9_11 = _GEN_192;
  wire         compressDataVec_hitReq_9_75;
  assign compressDataVec_hitReq_9_75 = _GEN_192;
  wire         _GEN_193 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hB;
  wire         compressDataVec_hitReq_10_11;
  assign compressDataVec_hitReq_10_11 = _GEN_193;
  wire         compressDataVec_hitReq_10_75;
  assign compressDataVec_hitReq_10_75 = _GEN_193;
  wire         _GEN_194 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hB;
  wire         compressDataVec_hitReq_11_11;
  assign compressDataVec_hitReq_11_11 = _GEN_194;
  wire         compressDataVec_hitReq_11_75;
  assign compressDataVec_hitReq_11_75 = _GEN_194;
  wire         _GEN_195 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hB;
  wire         compressDataVec_hitReq_12_11;
  assign compressDataVec_hitReq_12_11 = _GEN_195;
  wire         compressDataVec_hitReq_12_75;
  assign compressDataVec_hitReq_12_75 = _GEN_195;
  wire         _GEN_196 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hB;
  wire         compressDataVec_hitReq_13_11;
  assign compressDataVec_hitReq_13_11 = _GEN_196;
  wire         compressDataVec_hitReq_13_75;
  assign compressDataVec_hitReq_13_75 = _GEN_196;
  wire         _GEN_197 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hB;
  wire         compressDataVec_hitReq_14_11;
  assign compressDataVec_hitReq_14_11 = _GEN_197;
  wire         compressDataVec_hitReq_14_75;
  assign compressDataVec_hitReq_14_75 = _GEN_197;
  wire         _GEN_198 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hB;
  wire         compressDataVec_hitReq_15_11;
  assign compressDataVec_hitReq_15_11 = _GEN_198;
  wire         compressDataVec_hitReq_15_75;
  assign compressDataVec_hitReq_15_75 = _GEN_198;
  wire         compressDataVec_hitReq_16_11 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hB;
  wire         compressDataVec_hitReq_17_11 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hB;
  wire         compressDataVec_hitReq_18_11 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hB;
  wire         compressDataVec_hitReq_19_11 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hB;
  wire         compressDataVec_hitReq_20_11 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hB;
  wire         compressDataVec_hitReq_21_11 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hB;
  wire         compressDataVec_hitReq_22_11 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hB;
  wire         compressDataVec_hitReq_23_11 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hB;
  wire         compressDataVec_hitReq_24_11 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hB;
  wire         compressDataVec_hitReq_25_11 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hB;
  wire         compressDataVec_hitReq_26_11 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hB;
  wire         compressDataVec_hitReq_27_11 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hB;
  wire         compressDataVec_hitReq_28_11 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hB;
  wire         compressDataVec_hitReq_29_11 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hB;
  wire         compressDataVec_hitReq_30_11 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hB;
  wire         compressDataVec_hitReq_31_11 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hB;
  wire [7:0]   compressDataVec_selectReqData_11 =
    (compressDataVec_hitReq_0_11 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_11 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_11 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_11 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_11 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_11 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_11 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_11 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_11 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_11 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_11 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_11 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_11 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_11 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_11 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_11 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_11 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_11 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_11 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_11 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_11 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_11 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_11 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_11 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_11 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_11 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_11 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_11 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_11 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_11 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_11 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_11 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_199 = tailCount > 5'hB;
  wire         compressDataVec_useTail_11;
  assign compressDataVec_useTail_11 = _GEN_199;
  wire         compressDataVec_useTail_43;
  assign compressDataVec_useTail_43 = _GEN_199;
  wire         _GEN_200 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hC;
  wire         compressDataVec_hitReq_0_12;
  assign compressDataVec_hitReq_0_12 = _GEN_200;
  wire         compressDataVec_hitReq_0_76;
  assign compressDataVec_hitReq_0_76 = _GEN_200;
  wire         compressDataVec_hitReq_0_108;
  assign compressDataVec_hitReq_0_108 = _GEN_200;
  wire         _GEN_201 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hC;
  wire         compressDataVec_hitReq_1_12;
  assign compressDataVec_hitReq_1_12 = _GEN_201;
  wire         compressDataVec_hitReq_1_76;
  assign compressDataVec_hitReq_1_76 = _GEN_201;
  wire         compressDataVec_hitReq_1_108;
  assign compressDataVec_hitReq_1_108 = _GEN_201;
  wire         _GEN_202 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hC;
  wire         compressDataVec_hitReq_2_12;
  assign compressDataVec_hitReq_2_12 = _GEN_202;
  wire         compressDataVec_hitReq_2_76;
  assign compressDataVec_hitReq_2_76 = _GEN_202;
  wire         compressDataVec_hitReq_2_108;
  assign compressDataVec_hitReq_2_108 = _GEN_202;
  wire         _GEN_203 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hC;
  wire         compressDataVec_hitReq_3_12;
  assign compressDataVec_hitReq_3_12 = _GEN_203;
  wire         compressDataVec_hitReq_3_76;
  assign compressDataVec_hitReq_3_76 = _GEN_203;
  wire         compressDataVec_hitReq_3_108;
  assign compressDataVec_hitReq_3_108 = _GEN_203;
  wire         _GEN_204 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hC;
  wire         compressDataVec_hitReq_4_12;
  assign compressDataVec_hitReq_4_12 = _GEN_204;
  wire         compressDataVec_hitReq_4_76;
  assign compressDataVec_hitReq_4_76 = _GEN_204;
  wire         compressDataVec_hitReq_4_108;
  assign compressDataVec_hitReq_4_108 = _GEN_204;
  wire         _GEN_205 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hC;
  wire         compressDataVec_hitReq_5_12;
  assign compressDataVec_hitReq_5_12 = _GEN_205;
  wire         compressDataVec_hitReq_5_76;
  assign compressDataVec_hitReq_5_76 = _GEN_205;
  wire         compressDataVec_hitReq_5_108;
  assign compressDataVec_hitReq_5_108 = _GEN_205;
  wire         _GEN_206 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hC;
  wire         compressDataVec_hitReq_6_12;
  assign compressDataVec_hitReq_6_12 = _GEN_206;
  wire         compressDataVec_hitReq_6_76;
  assign compressDataVec_hitReq_6_76 = _GEN_206;
  wire         compressDataVec_hitReq_6_108;
  assign compressDataVec_hitReq_6_108 = _GEN_206;
  wire         _GEN_207 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hC;
  wire         compressDataVec_hitReq_7_12;
  assign compressDataVec_hitReq_7_12 = _GEN_207;
  wire         compressDataVec_hitReq_7_76;
  assign compressDataVec_hitReq_7_76 = _GEN_207;
  wire         compressDataVec_hitReq_7_108;
  assign compressDataVec_hitReq_7_108 = _GEN_207;
  wire         _GEN_208 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hC;
  wire         compressDataVec_hitReq_8_12;
  assign compressDataVec_hitReq_8_12 = _GEN_208;
  wire         compressDataVec_hitReq_8_76;
  assign compressDataVec_hitReq_8_76 = _GEN_208;
  wire         _GEN_209 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hC;
  wire         compressDataVec_hitReq_9_12;
  assign compressDataVec_hitReq_9_12 = _GEN_209;
  wire         compressDataVec_hitReq_9_76;
  assign compressDataVec_hitReq_9_76 = _GEN_209;
  wire         _GEN_210 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hC;
  wire         compressDataVec_hitReq_10_12;
  assign compressDataVec_hitReq_10_12 = _GEN_210;
  wire         compressDataVec_hitReq_10_76;
  assign compressDataVec_hitReq_10_76 = _GEN_210;
  wire         _GEN_211 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hC;
  wire         compressDataVec_hitReq_11_12;
  assign compressDataVec_hitReq_11_12 = _GEN_211;
  wire         compressDataVec_hitReq_11_76;
  assign compressDataVec_hitReq_11_76 = _GEN_211;
  wire         _GEN_212 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hC;
  wire         compressDataVec_hitReq_12_12;
  assign compressDataVec_hitReq_12_12 = _GEN_212;
  wire         compressDataVec_hitReq_12_76;
  assign compressDataVec_hitReq_12_76 = _GEN_212;
  wire         _GEN_213 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hC;
  wire         compressDataVec_hitReq_13_12;
  assign compressDataVec_hitReq_13_12 = _GEN_213;
  wire         compressDataVec_hitReq_13_76;
  assign compressDataVec_hitReq_13_76 = _GEN_213;
  wire         _GEN_214 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hC;
  wire         compressDataVec_hitReq_14_12;
  assign compressDataVec_hitReq_14_12 = _GEN_214;
  wire         compressDataVec_hitReq_14_76;
  assign compressDataVec_hitReq_14_76 = _GEN_214;
  wire         _GEN_215 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hC;
  wire         compressDataVec_hitReq_15_12;
  assign compressDataVec_hitReq_15_12 = _GEN_215;
  wire         compressDataVec_hitReq_15_76;
  assign compressDataVec_hitReq_15_76 = _GEN_215;
  wire         compressDataVec_hitReq_16_12 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hC;
  wire         compressDataVec_hitReq_17_12 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hC;
  wire         compressDataVec_hitReq_18_12 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hC;
  wire         compressDataVec_hitReq_19_12 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hC;
  wire         compressDataVec_hitReq_20_12 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hC;
  wire         compressDataVec_hitReq_21_12 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hC;
  wire         compressDataVec_hitReq_22_12 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hC;
  wire         compressDataVec_hitReq_23_12 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hC;
  wire         compressDataVec_hitReq_24_12 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hC;
  wire         compressDataVec_hitReq_25_12 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hC;
  wire         compressDataVec_hitReq_26_12 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hC;
  wire         compressDataVec_hitReq_27_12 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hC;
  wire         compressDataVec_hitReq_28_12 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hC;
  wire         compressDataVec_hitReq_29_12 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hC;
  wire         compressDataVec_hitReq_30_12 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hC;
  wire         compressDataVec_hitReq_31_12 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hC;
  wire [7:0]   compressDataVec_selectReqData_12 =
    (compressDataVec_hitReq_0_12 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_12 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_12 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_12 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_12 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_12 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_12 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_12 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_12 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_12 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_12 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_12 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_12 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_12 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_12 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_12 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_12 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_12 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_12 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_12 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_12 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_12 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_12 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_12 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_12 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_12 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_12 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_12 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_12 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_12 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_12 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_12 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_216 = tailCount > 5'hC;
  wire         compressDataVec_useTail_12;
  assign compressDataVec_useTail_12 = _GEN_216;
  wire         compressDataVec_useTail_44;
  assign compressDataVec_useTail_44 = _GEN_216;
  wire         _GEN_217 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hD;
  wire         compressDataVec_hitReq_0_13;
  assign compressDataVec_hitReq_0_13 = _GEN_217;
  wire         compressDataVec_hitReq_0_77;
  assign compressDataVec_hitReq_0_77 = _GEN_217;
  wire         compressDataVec_hitReq_0_109;
  assign compressDataVec_hitReq_0_109 = _GEN_217;
  wire         _GEN_218 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hD;
  wire         compressDataVec_hitReq_1_13;
  assign compressDataVec_hitReq_1_13 = _GEN_218;
  wire         compressDataVec_hitReq_1_77;
  assign compressDataVec_hitReq_1_77 = _GEN_218;
  wire         compressDataVec_hitReq_1_109;
  assign compressDataVec_hitReq_1_109 = _GEN_218;
  wire         _GEN_219 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hD;
  wire         compressDataVec_hitReq_2_13;
  assign compressDataVec_hitReq_2_13 = _GEN_219;
  wire         compressDataVec_hitReq_2_77;
  assign compressDataVec_hitReq_2_77 = _GEN_219;
  wire         compressDataVec_hitReq_2_109;
  assign compressDataVec_hitReq_2_109 = _GEN_219;
  wire         _GEN_220 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hD;
  wire         compressDataVec_hitReq_3_13;
  assign compressDataVec_hitReq_3_13 = _GEN_220;
  wire         compressDataVec_hitReq_3_77;
  assign compressDataVec_hitReq_3_77 = _GEN_220;
  wire         compressDataVec_hitReq_3_109;
  assign compressDataVec_hitReq_3_109 = _GEN_220;
  wire         _GEN_221 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hD;
  wire         compressDataVec_hitReq_4_13;
  assign compressDataVec_hitReq_4_13 = _GEN_221;
  wire         compressDataVec_hitReq_4_77;
  assign compressDataVec_hitReq_4_77 = _GEN_221;
  wire         compressDataVec_hitReq_4_109;
  assign compressDataVec_hitReq_4_109 = _GEN_221;
  wire         _GEN_222 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hD;
  wire         compressDataVec_hitReq_5_13;
  assign compressDataVec_hitReq_5_13 = _GEN_222;
  wire         compressDataVec_hitReq_5_77;
  assign compressDataVec_hitReq_5_77 = _GEN_222;
  wire         compressDataVec_hitReq_5_109;
  assign compressDataVec_hitReq_5_109 = _GEN_222;
  wire         _GEN_223 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hD;
  wire         compressDataVec_hitReq_6_13;
  assign compressDataVec_hitReq_6_13 = _GEN_223;
  wire         compressDataVec_hitReq_6_77;
  assign compressDataVec_hitReq_6_77 = _GEN_223;
  wire         compressDataVec_hitReq_6_109;
  assign compressDataVec_hitReq_6_109 = _GEN_223;
  wire         _GEN_224 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hD;
  wire         compressDataVec_hitReq_7_13;
  assign compressDataVec_hitReq_7_13 = _GEN_224;
  wire         compressDataVec_hitReq_7_77;
  assign compressDataVec_hitReq_7_77 = _GEN_224;
  wire         compressDataVec_hitReq_7_109;
  assign compressDataVec_hitReq_7_109 = _GEN_224;
  wire         _GEN_225 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hD;
  wire         compressDataVec_hitReq_8_13;
  assign compressDataVec_hitReq_8_13 = _GEN_225;
  wire         compressDataVec_hitReq_8_77;
  assign compressDataVec_hitReq_8_77 = _GEN_225;
  wire         _GEN_226 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hD;
  wire         compressDataVec_hitReq_9_13;
  assign compressDataVec_hitReq_9_13 = _GEN_226;
  wire         compressDataVec_hitReq_9_77;
  assign compressDataVec_hitReq_9_77 = _GEN_226;
  wire         _GEN_227 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hD;
  wire         compressDataVec_hitReq_10_13;
  assign compressDataVec_hitReq_10_13 = _GEN_227;
  wire         compressDataVec_hitReq_10_77;
  assign compressDataVec_hitReq_10_77 = _GEN_227;
  wire         _GEN_228 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hD;
  wire         compressDataVec_hitReq_11_13;
  assign compressDataVec_hitReq_11_13 = _GEN_228;
  wire         compressDataVec_hitReq_11_77;
  assign compressDataVec_hitReq_11_77 = _GEN_228;
  wire         _GEN_229 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hD;
  wire         compressDataVec_hitReq_12_13;
  assign compressDataVec_hitReq_12_13 = _GEN_229;
  wire         compressDataVec_hitReq_12_77;
  assign compressDataVec_hitReq_12_77 = _GEN_229;
  wire         _GEN_230 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hD;
  wire         compressDataVec_hitReq_13_13;
  assign compressDataVec_hitReq_13_13 = _GEN_230;
  wire         compressDataVec_hitReq_13_77;
  assign compressDataVec_hitReq_13_77 = _GEN_230;
  wire         _GEN_231 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hD;
  wire         compressDataVec_hitReq_14_13;
  assign compressDataVec_hitReq_14_13 = _GEN_231;
  wire         compressDataVec_hitReq_14_77;
  assign compressDataVec_hitReq_14_77 = _GEN_231;
  wire         _GEN_232 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hD;
  wire         compressDataVec_hitReq_15_13;
  assign compressDataVec_hitReq_15_13 = _GEN_232;
  wire         compressDataVec_hitReq_15_77;
  assign compressDataVec_hitReq_15_77 = _GEN_232;
  wire         compressDataVec_hitReq_16_13 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hD;
  wire         compressDataVec_hitReq_17_13 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hD;
  wire         compressDataVec_hitReq_18_13 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hD;
  wire         compressDataVec_hitReq_19_13 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hD;
  wire         compressDataVec_hitReq_20_13 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hD;
  wire         compressDataVec_hitReq_21_13 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hD;
  wire         compressDataVec_hitReq_22_13 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hD;
  wire         compressDataVec_hitReq_23_13 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hD;
  wire         compressDataVec_hitReq_24_13 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hD;
  wire         compressDataVec_hitReq_25_13 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hD;
  wire         compressDataVec_hitReq_26_13 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hD;
  wire         compressDataVec_hitReq_27_13 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hD;
  wire         compressDataVec_hitReq_28_13 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hD;
  wire         compressDataVec_hitReq_29_13 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hD;
  wire         compressDataVec_hitReq_30_13 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hD;
  wire         compressDataVec_hitReq_31_13 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hD;
  wire [7:0]   compressDataVec_selectReqData_13 =
    (compressDataVec_hitReq_0_13 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_13 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_13 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_13 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_13 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_13 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_13 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_13 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_13 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_13 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_13 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_13 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_13 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_13 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_13 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_13 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_13 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_13 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_13 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_13 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_13 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_13 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_13 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_13 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_13 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_13 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_13 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_13 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_13 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_13 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_13 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_13 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_233 = tailCount > 5'hD;
  wire         compressDataVec_useTail_13;
  assign compressDataVec_useTail_13 = _GEN_233;
  wire         compressDataVec_useTail_45;
  assign compressDataVec_useTail_45 = _GEN_233;
  wire         _GEN_234 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hE;
  wire         compressDataVec_hitReq_0_14;
  assign compressDataVec_hitReq_0_14 = _GEN_234;
  wire         compressDataVec_hitReq_0_78;
  assign compressDataVec_hitReq_0_78 = _GEN_234;
  wire         compressDataVec_hitReq_0_110;
  assign compressDataVec_hitReq_0_110 = _GEN_234;
  wire         _GEN_235 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hE;
  wire         compressDataVec_hitReq_1_14;
  assign compressDataVec_hitReq_1_14 = _GEN_235;
  wire         compressDataVec_hitReq_1_78;
  assign compressDataVec_hitReq_1_78 = _GEN_235;
  wire         compressDataVec_hitReq_1_110;
  assign compressDataVec_hitReq_1_110 = _GEN_235;
  wire         _GEN_236 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hE;
  wire         compressDataVec_hitReq_2_14;
  assign compressDataVec_hitReq_2_14 = _GEN_236;
  wire         compressDataVec_hitReq_2_78;
  assign compressDataVec_hitReq_2_78 = _GEN_236;
  wire         compressDataVec_hitReq_2_110;
  assign compressDataVec_hitReq_2_110 = _GEN_236;
  wire         _GEN_237 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hE;
  wire         compressDataVec_hitReq_3_14;
  assign compressDataVec_hitReq_3_14 = _GEN_237;
  wire         compressDataVec_hitReq_3_78;
  assign compressDataVec_hitReq_3_78 = _GEN_237;
  wire         compressDataVec_hitReq_3_110;
  assign compressDataVec_hitReq_3_110 = _GEN_237;
  wire         _GEN_238 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hE;
  wire         compressDataVec_hitReq_4_14;
  assign compressDataVec_hitReq_4_14 = _GEN_238;
  wire         compressDataVec_hitReq_4_78;
  assign compressDataVec_hitReq_4_78 = _GEN_238;
  wire         compressDataVec_hitReq_4_110;
  assign compressDataVec_hitReq_4_110 = _GEN_238;
  wire         _GEN_239 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hE;
  wire         compressDataVec_hitReq_5_14;
  assign compressDataVec_hitReq_5_14 = _GEN_239;
  wire         compressDataVec_hitReq_5_78;
  assign compressDataVec_hitReq_5_78 = _GEN_239;
  wire         compressDataVec_hitReq_5_110;
  assign compressDataVec_hitReq_5_110 = _GEN_239;
  wire         _GEN_240 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hE;
  wire         compressDataVec_hitReq_6_14;
  assign compressDataVec_hitReq_6_14 = _GEN_240;
  wire         compressDataVec_hitReq_6_78;
  assign compressDataVec_hitReq_6_78 = _GEN_240;
  wire         compressDataVec_hitReq_6_110;
  assign compressDataVec_hitReq_6_110 = _GEN_240;
  wire         _GEN_241 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hE;
  wire         compressDataVec_hitReq_7_14;
  assign compressDataVec_hitReq_7_14 = _GEN_241;
  wire         compressDataVec_hitReq_7_78;
  assign compressDataVec_hitReq_7_78 = _GEN_241;
  wire         compressDataVec_hitReq_7_110;
  assign compressDataVec_hitReq_7_110 = _GEN_241;
  wire         _GEN_242 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hE;
  wire         compressDataVec_hitReq_8_14;
  assign compressDataVec_hitReq_8_14 = _GEN_242;
  wire         compressDataVec_hitReq_8_78;
  assign compressDataVec_hitReq_8_78 = _GEN_242;
  wire         _GEN_243 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hE;
  wire         compressDataVec_hitReq_9_14;
  assign compressDataVec_hitReq_9_14 = _GEN_243;
  wire         compressDataVec_hitReq_9_78;
  assign compressDataVec_hitReq_9_78 = _GEN_243;
  wire         _GEN_244 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hE;
  wire         compressDataVec_hitReq_10_14;
  assign compressDataVec_hitReq_10_14 = _GEN_244;
  wire         compressDataVec_hitReq_10_78;
  assign compressDataVec_hitReq_10_78 = _GEN_244;
  wire         _GEN_245 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hE;
  wire         compressDataVec_hitReq_11_14;
  assign compressDataVec_hitReq_11_14 = _GEN_245;
  wire         compressDataVec_hitReq_11_78;
  assign compressDataVec_hitReq_11_78 = _GEN_245;
  wire         _GEN_246 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hE;
  wire         compressDataVec_hitReq_12_14;
  assign compressDataVec_hitReq_12_14 = _GEN_246;
  wire         compressDataVec_hitReq_12_78;
  assign compressDataVec_hitReq_12_78 = _GEN_246;
  wire         _GEN_247 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hE;
  wire         compressDataVec_hitReq_13_14;
  assign compressDataVec_hitReq_13_14 = _GEN_247;
  wire         compressDataVec_hitReq_13_78;
  assign compressDataVec_hitReq_13_78 = _GEN_247;
  wire         _GEN_248 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hE;
  wire         compressDataVec_hitReq_14_14;
  assign compressDataVec_hitReq_14_14 = _GEN_248;
  wire         compressDataVec_hitReq_14_78;
  assign compressDataVec_hitReq_14_78 = _GEN_248;
  wire         _GEN_249 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hE;
  wire         compressDataVec_hitReq_15_14;
  assign compressDataVec_hitReq_15_14 = _GEN_249;
  wire         compressDataVec_hitReq_15_78;
  assign compressDataVec_hitReq_15_78 = _GEN_249;
  wire         compressDataVec_hitReq_16_14 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hE;
  wire         compressDataVec_hitReq_17_14 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hE;
  wire         compressDataVec_hitReq_18_14 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hE;
  wire         compressDataVec_hitReq_19_14 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hE;
  wire         compressDataVec_hitReq_20_14 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hE;
  wire         compressDataVec_hitReq_21_14 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hE;
  wire         compressDataVec_hitReq_22_14 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hE;
  wire         compressDataVec_hitReq_23_14 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hE;
  wire         compressDataVec_hitReq_24_14 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hE;
  wire         compressDataVec_hitReq_25_14 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hE;
  wire         compressDataVec_hitReq_26_14 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hE;
  wire         compressDataVec_hitReq_27_14 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hE;
  wire         compressDataVec_hitReq_28_14 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hE;
  wire         compressDataVec_hitReq_29_14 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hE;
  wire         compressDataVec_hitReq_30_14 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hE;
  wire         compressDataVec_hitReq_31_14 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hE;
  wire [7:0]   compressDataVec_selectReqData_14 =
    (compressDataVec_hitReq_0_14 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_14 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_14 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_14 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_14 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_14 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_14 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_14 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_14 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_14 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_14 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_14 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_14 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_14 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_14 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_14 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_14 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_14 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_14 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_14 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_14 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_14 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_14 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_14 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_14 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_14 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_14 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_14 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_14 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_14 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_14 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_14 ? source2Pipe[255:248] : 8'h0);
  wire         _GEN_250 = tailCount > 5'hE;
  wire         compressDataVec_useTail_14;
  assign compressDataVec_useTail_14 = _GEN_250;
  wire         compressDataVec_useTail_46;
  assign compressDataVec_useTail_46 = _GEN_250;
  wire         _GEN_251 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'hF;
  wire         compressDataVec_hitReq_0_15;
  assign compressDataVec_hitReq_0_15 = _GEN_251;
  wire         compressDataVec_hitReq_0_79;
  assign compressDataVec_hitReq_0_79 = _GEN_251;
  wire         compressDataVec_hitReq_0_111;
  assign compressDataVec_hitReq_0_111 = _GEN_251;
  wire         _GEN_252 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'hF;
  wire         compressDataVec_hitReq_1_15;
  assign compressDataVec_hitReq_1_15 = _GEN_252;
  wire         compressDataVec_hitReq_1_79;
  assign compressDataVec_hitReq_1_79 = _GEN_252;
  wire         compressDataVec_hitReq_1_111;
  assign compressDataVec_hitReq_1_111 = _GEN_252;
  wire         _GEN_253 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'hF;
  wire         compressDataVec_hitReq_2_15;
  assign compressDataVec_hitReq_2_15 = _GEN_253;
  wire         compressDataVec_hitReq_2_79;
  assign compressDataVec_hitReq_2_79 = _GEN_253;
  wire         compressDataVec_hitReq_2_111;
  assign compressDataVec_hitReq_2_111 = _GEN_253;
  wire         _GEN_254 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'hF;
  wire         compressDataVec_hitReq_3_15;
  assign compressDataVec_hitReq_3_15 = _GEN_254;
  wire         compressDataVec_hitReq_3_79;
  assign compressDataVec_hitReq_3_79 = _GEN_254;
  wire         compressDataVec_hitReq_3_111;
  assign compressDataVec_hitReq_3_111 = _GEN_254;
  wire         _GEN_255 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'hF;
  wire         compressDataVec_hitReq_4_15;
  assign compressDataVec_hitReq_4_15 = _GEN_255;
  wire         compressDataVec_hitReq_4_79;
  assign compressDataVec_hitReq_4_79 = _GEN_255;
  wire         compressDataVec_hitReq_4_111;
  assign compressDataVec_hitReq_4_111 = _GEN_255;
  wire         _GEN_256 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'hF;
  wire         compressDataVec_hitReq_5_15;
  assign compressDataVec_hitReq_5_15 = _GEN_256;
  wire         compressDataVec_hitReq_5_79;
  assign compressDataVec_hitReq_5_79 = _GEN_256;
  wire         compressDataVec_hitReq_5_111;
  assign compressDataVec_hitReq_5_111 = _GEN_256;
  wire         _GEN_257 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'hF;
  wire         compressDataVec_hitReq_6_15;
  assign compressDataVec_hitReq_6_15 = _GEN_257;
  wire         compressDataVec_hitReq_6_79;
  assign compressDataVec_hitReq_6_79 = _GEN_257;
  wire         compressDataVec_hitReq_6_111;
  assign compressDataVec_hitReq_6_111 = _GEN_257;
  wire         _GEN_258 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'hF;
  wire         compressDataVec_hitReq_7_15;
  assign compressDataVec_hitReq_7_15 = _GEN_258;
  wire         compressDataVec_hitReq_7_79;
  assign compressDataVec_hitReq_7_79 = _GEN_258;
  wire         compressDataVec_hitReq_7_111;
  assign compressDataVec_hitReq_7_111 = _GEN_258;
  wire         _GEN_259 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'hF;
  wire         compressDataVec_hitReq_8_15;
  assign compressDataVec_hitReq_8_15 = _GEN_259;
  wire         compressDataVec_hitReq_8_79;
  assign compressDataVec_hitReq_8_79 = _GEN_259;
  wire         _GEN_260 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'hF;
  wire         compressDataVec_hitReq_9_15;
  assign compressDataVec_hitReq_9_15 = _GEN_260;
  wire         compressDataVec_hitReq_9_79;
  assign compressDataVec_hitReq_9_79 = _GEN_260;
  wire         _GEN_261 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'hF;
  wire         compressDataVec_hitReq_10_15;
  assign compressDataVec_hitReq_10_15 = _GEN_261;
  wire         compressDataVec_hitReq_10_79;
  assign compressDataVec_hitReq_10_79 = _GEN_261;
  wire         _GEN_262 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'hF;
  wire         compressDataVec_hitReq_11_15;
  assign compressDataVec_hitReq_11_15 = _GEN_262;
  wire         compressDataVec_hitReq_11_79;
  assign compressDataVec_hitReq_11_79 = _GEN_262;
  wire         _GEN_263 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'hF;
  wire         compressDataVec_hitReq_12_15;
  assign compressDataVec_hitReq_12_15 = _GEN_263;
  wire         compressDataVec_hitReq_12_79;
  assign compressDataVec_hitReq_12_79 = _GEN_263;
  wire         _GEN_264 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'hF;
  wire         compressDataVec_hitReq_13_15;
  assign compressDataVec_hitReq_13_15 = _GEN_264;
  wire         compressDataVec_hitReq_13_79;
  assign compressDataVec_hitReq_13_79 = _GEN_264;
  wire         _GEN_265 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'hF;
  wire         compressDataVec_hitReq_14_15;
  assign compressDataVec_hitReq_14_15 = _GEN_265;
  wire         compressDataVec_hitReq_14_79;
  assign compressDataVec_hitReq_14_79 = _GEN_265;
  wire         _GEN_266 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'hF;
  wire         compressDataVec_hitReq_15_15;
  assign compressDataVec_hitReq_15_15 = _GEN_266;
  wire         compressDataVec_hitReq_15_79;
  assign compressDataVec_hitReq_15_79 = _GEN_266;
  wire         compressDataVec_hitReq_16_15 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'hF;
  wire         compressDataVec_hitReq_17_15 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'hF;
  wire         compressDataVec_hitReq_18_15 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'hF;
  wire         compressDataVec_hitReq_19_15 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'hF;
  wire         compressDataVec_hitReq_20_15 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'hF;
  wire         compressDataVec_hitReq_21_15 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'hF;
  wire         compressDataVec_hitReq_22_15 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'hF;
  wire         compressDataVec_hitReq_23_15 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'hF;
  wire         compressDataVec_hitReq_24_15 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'hF;
  wire         compressDataVec_hitReq_25_15 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'hF;
  wire         compressDataVec_hitReq_26_15 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'hF;
  wire         compressDataVec_hitReq_27_15 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'hF;
  wire         compressDataVec_hitReq_28_15 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'hF;
  wire         compressDataVec_hitReq_29_15 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'hF;
  wire         compressDataVec_hitReq_30_15 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'hF;
  wire         compressDataVec_hitReq_31_15 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'hF;
  wire [7:0]   compressDataVec_selectReqData_15 =
    (compressDataVec_hitReq_0_15 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_15 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_15 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_15 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_15 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_15 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_15 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_15 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_15 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_15 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_15 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_15 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_15 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_15 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_15 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_15 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_15 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_15 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_15 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_15 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_15 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_15 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_15 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_15 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_15 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_15 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_15 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_15 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_15 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_15 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_15 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_15 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_15 = tailCount[4];
  wire         compressDataVec_useTail_47 = tailCount[4];
  wire         _GEN_267 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h10;
  wire         compressDataVec_hitReq_0_16;
  assign compressDataVec_hitReq_0_16 = _GEN_267;
  wire         compressDataVec_hitReq_0_80;
  assign compressDataVec_hitReq_0_80 = _GEN_267;
  wire         _GEN_268 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h10;
  wire         compressDataVec_hitReq_1_16;
  assign compressDataVec_hitReq_1_16 = _GEN_268;
  wire         compressDataVec_hitReq_1_80;
  assign compressDataVec_hitReq_1_80 = _GEN_268;
  wire         _GEN_269 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h10;
  wire         compressDataVec_hitReq_2_16;
  assign compressDataVec_hitReq_2_16 = _GEN_269;
  wire         compressDataVec_hitReq_2_80;
  assign compressDataVec_hitReq_2_80 = _GEN_269;
  wire         _GEN_270 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h10;
  wire         compressDataVec_hitReq_3_16;
  assign compressDataVec_hitReq_3_16 = _GEN_270;
  wire         compressDataVec_hitReq_3_80;
  assign compressDataVec_hitReq_3_80 = _GEN_270;
  wire         _GEN_271 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h10;
  wire         compressDataVec_hitReq_4_16;
  assign compressDataVec_hitReq_4_16 = _GEN_271;
  wire         compressDataVec_hitReq_4_80;
  assign compressDataVec_hitReq_4_80 = _GEN_271;
  wire         _GEN_272 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h10;
  wire         compressDataVec_hitReq_5_16;
  assign compressDataVec_hitReq_5_16 = _GEN_272;
  wire         compressDataVec_hitReq_5_80;
  assign compressDataVec_hitReq_5_80 = _GEN_272;
  wire         _GEN_273 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h10;
  wire         compressDataVec_hitReq_6_16;
  assign compressDataVec_hitReq_6_16 = _GEN_273;
  wire         compressDataVec_hitReq_6_80;
  assign compressDataVec_hitReq_6_80 = _GEN_273;
  wire         _GEN_274 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h10;
  wire         compressDataVec_hitReq_7_16;
  assign compressDataVec_hitReq_7_16 = _GEN_274;
  wire         compressDataVec_hitReq_7_80;
  assign compressDataVec_hitReq_7_80 = _GEN_274;
  wire         _GEN_275 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h10;
  wire         compressDataVec_hitReq_8_16;
  assign compressDataVec_hitReq_8_16 = _GEN_275;
  wire         compressDataVec_hitReq_8_80;
  assign compressDataVec_hitReq_8_80 = _GEN_275;
  wire         _GEN_276 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h10;
  wire         compressDataVec_hitReq_9_16;
  assign compressDataVec_hitReq_9_16 = _GEN_276;
  wire         compressDataVec_hitReq_9_80;
  assign compressDataVec_hitReq_9_80 = _GEN_276;
  wire         _GEN_277 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h10;
  wire         compressDataVec_hitReq_10_16;
  assign compressDataVec_hitReq_10_16 = _GEN_277;
  wire         compressDataVec_hitReq_10_80;
  assign compressDataVec_hitReq_10_80 = _GEN_277;
  wire         _GEN_278 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h10;
  wire         compressDataVec_hitReq_11_16;
  assign compressDataVec_hitReq_11_16 = _GEN_278;
  wire         compressDataVec_hitReq_11_80;
  assign compressDataVec_hitReq_11_80 = _GEN_278;
  wire         _GEN_279 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h10;
  wire         compressDataVec_hitReq_12_16;
  assign compressDataVec_hitReq_12_16 = _GEN_279;
  wire         compressDataVec_hitReq_12_80;
  assign compressDataVec_hitReq_12_80 = _GEN_279;
  wire         _GEN_280 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h10;
  wire         compressDataVec_hitReq_13_16;
  assign compressDataVec_hitReq_13_16 = _GEN_280;
  wire         compressDataVec_hitReq_13_80;
  assign compressDataVec_hitReq_13_80 = _GEN_280;
  wire         _GEN_281 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h10;
  wire         compressDataVec_hitReq_14_16;
  assign compressDataVec_hitReq_14_16 = _GEN_281;
  wire         compressDataVec_hitReq_14_80;
  assign compressDataVec_hitReq_14_80 = _GEN_281;
  wire         _GEN_282 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h10;
  wire         compressDataVec_hitReq_15_16;
  assign compressDataVec_hitReq_15_16 = _GEN_282;
  wire         compressDataVec_hitReq_15_80;
  assign compressDataVec_hitReq_15_80 = _GEN_282;
  wire         compressDataVec_hitReq_16_16 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h10;
  wire         compressDataVec_hitReq_17_16 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h10;
  wire         compressDataVec_hitReq_18_16 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h10;
  wire         compressDataVec_hitReq_19_16 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h10;
  wire         compressDataVec_hitReq_20_16 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h10;
  wire         compressDataVec_hitReq_21_16 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h10;
  wire         compressDataVec_hitReq_22_16 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h10;
  wire         compressDataVec_hitReq_23_16 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h10;
  wire         compressDataVec_hitReq_24_16 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h10;
  wire         compressDataVec_hitReq_25_16 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h10;
  wire         compressDataVec_hitReq_26_16 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h10;
  wire         compressDataVec_hitReq_27_16 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h10;
  wire         compressDataVec_hitReq_28_16 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h10;
  wire         compressDataVec_hitReq_29_16 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h10;
  wire         compressDataVec_hitReq_30_16 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h10;
  wire         compressDataVec_hitReq_31_16 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h10;
  wire [7:0]   compressDataVec_selectReqData_16 =
    (compressDataVec_hitReq_0_16 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_16 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_16 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_16 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_16 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_16 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_16 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_16 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_16 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_16 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_16 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_16 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_16 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_16 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_16 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_16 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_16 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_16 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_16 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_16 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_16 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_16 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_16 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_16 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_16 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_16 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_16 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_16 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_16 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_16 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_16 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_16 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_16 = tailCount > 5'h10;
  wire         _GEN_283 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h11;
  wire         compressDataVec_hitReq_0_17;
  assign compressDataVec_hitReq_0_17 = _GEN_283;
  wire         compressDataVec_hitReq_0_81;
  assign compressDataVec_hitReq_0_81 = _GEN_283;
  wire         _GEN_284 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h11;
  wire         compressDataVec_hitReq_1_17;
  assign compressDataVec_hitReq_1_17 = _GEN_284;
  wire         compressDataVec_hitReq_1_81;
  assign compressDataVec_hitReq_1_81 = _GEN_284;
  wire         _GEN_285 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h11;
  wire         compressDataVec_hitReq_2_17;
  assign compressDataVec_hitReq_2_17 = _GEN_285;
  wire         compressDataVec_hitReq_2_81;
  assign compressDataVec_hitReq_2_81 = _GEN_285;
  wire         _GEN_286 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h11;
  wire         compressDataVec_hitReq_3_17;
  assign compressDataVec_hitReq_3_17 = _GEN_286;
  wire         compressDataVec_hitReq_3_81;
  assign compressDataVec_hitReq_3_81 = _GEN_286;
  wire         _GEN_287 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h11;
  wire         compressDataVec_hitReq_4_17;
  assign compressDataVec_hitReq_4_17 = _GEN_287;
  wire         compressDataVec_hitReq_4_81;
  assign compressDataVec_hitReq_4_81 = _GEN_287;
  wire         _GEN_288 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h11;
  wire         compressDataVec_hitReq_5_17;
  assign compressDataVec_hitReq_5_17 = _GEN_288;
  wire         compressDataVec_hitReq_5_81;
  assign compressDataVec_hitReq_5_81 = _GEN_288;
  wire         _GEN_289 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h11;
  wire         compressDataVec_hitReq_6_17;
  assign compressDataVec_hitReq_6_17 = _GEN_289;
  wire         compressDataVec_hitReq_6_81;
  assign compressDataVec_hitReq_6_81 = _GEN_289;
  wire         _GEN_290 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h11;
  wire         compressDataVec_hitReq_7_17;
  assign compressDataVec_hitReq_7_17 = _GEN_290;
  wire         compressDataVec_hitReq_7_81;
  assign compressDataVec_hitReq_7_81 = _GEN_290;
  wire         _GEN_291 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h11;
  wire         compressDataVec_hitReq_8_17;
  assign compressDataVec_hitReq_8_17 = _GEN_291;
  wire         compressDataVec_hitReq_8_81;
  assign compressDataVec_hitReq_8_81 = _GEN_291;
  wire         _GEN_292 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h11;
  wire         compressDataVec_hitReq_9_17;
  assign compressDataVec_hitReq_9_17 = _GEN_292;
  wire         compressDataVec_hitReq_9_81;
  assign compressDataVec_hitReq_9_81 = _GEN_292;
  wire         _GEN_293 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h11;
  wire         compressDataVec_hitReq_10_17;
  assign compressDataVec_hitReq_10_17 = _GEN_293;
  wire         compressDataVec_hitReq_10_81;
  assign compressDataVec_hitReq_10_81 = _GEN_293;
  wire         _GEN_294 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h11;
  wire         compressDataVec_hitReq_11_17;
  assign compressDataVec_hitReq_11_17 = _GEN_294;
  wire         compressDataVec_hitReq_11_81;
  assign compressDataVec_hitReq_11_81 = _GEN_294;
  wire         _GEN_295 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h11;
  wire         compressDataVec_hitReq_12_17;
  assign compressDataVec_hitReq_12_17 = _GEN_295;
  wire         compressDataVec_hitReq_12_81;
  assign compressDataVec_hitReq_12_81 = _GEN_295;
  wire         _GEN_296 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h11;
  wire         compressDataVec_hitReq_13_17;
  assign compressDataVec_hitReq_13_17 = _GEN_296;
  wire         compressDataVec_hitReq_13_81;
  assign compressDataVec_hitReq_13_81 = _GEN_296;
  wire         _GEN_297 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h11;
  wire         compressDataVec_hitReq_14_17;
  assign compressDataVec_hitReq_14_17 = _GEN_297;
  wire         compressDataVec_hitReq_14_81;
  assign compressDataVec_hitReq_14_81 = _GEN_297;
  wire         _GEN_298 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h11;
  wire         compressDataVec_hitReq_15_17;
  assign compressDataVec_hitReq_15_17 = _GEN_298;
  wire         compressDataVec_hitReq_15_81;
  assign compressDataVec_hitReq_15_81 = _GEN_298;
  wire         compressDataVec_hitReq_16_17 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h11;
  wire         compressDataVec_hitReq_17_17 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h11;
  wire         compressDataVec_hitReq_18_17 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h11;
  wire         compressDataVec_hitReq_19_17 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h11;
  wire         compressDataVec_hitReq_20_17 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h11;
  wire         compressDataVec_hitReq_21_17 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h11;
  wire         compressDataVec_hitReq_22_17 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h11;
  wire         compressDataVec_hitReq_23_17 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h11;
  wire         compressDataVec_hitReq_24_17 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h11;
  wire         compressDataVec_hitReq_25_17 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h11;
  wire         compressDataVec_hitReq_26_17 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h11;
  wire         compressDataVec_hitReq_27_17 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h11;
  wire         compressDataVec_hitReq_28_17 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h11;
  wire         compressDataVec_hitReq_29_17 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h11;
  wire         compressDataVec_hitReq_30_17 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h11;
  wire         compressDataVec_hitReq_31_17 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h11;
  wire [7:0]   compressDataVec_selectReqData_17 =
    (compressDataVec_hitReq_0_17 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_17 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_17 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_17 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_17 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_17 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_17 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_17 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_17 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_17 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_17 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_17 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_17 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_17 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_17 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_17 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_17 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_17 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_17 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_17 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_17 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_17 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_17 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_17 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_17 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_17 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_17 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_17 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_17 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_17 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_17 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_17 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_17 = tailCount > 5'h11;
  wire         _GEN_299 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h12;
  wire         compressDataVec_hitReq_0_18;
  assign compressDataVec_hitReq_0_18 = _GEN_299;
  wire         compressDataVec_hitReq_0_82;
  assign compressDataVec_hitReq_0_82 = _GEN_299;
  wire         _GEN_300 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h12;
  wire         compressDataVec_hitReq_1_18;
  assign compressDataVec_hitReq_1_18 = _GEN_300;
  wire         compressDataVec_hitReq_1_82;
  assign compressDataVec_hitReq_1_82 = _GEN_300;
  wire         _GEN_301 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h12;
  wire         compressDataVec_hitReq_2_18;
  assign compressDataVec_hitReq_2_18 = _GEN_301;
  wire         compressDataVec_hitReq_2_82;
  assign compressDataVec_hitReq_2_82 = _GEN_301;
  wire         _GEN_302 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h12;
  wire         compressDataVec_hitReq_3_18;
  assign compressDataVec_hitReq_3_18 = _GEN_302;
  wire         compressDataVec_hitReq_3_82;
  assign compressDataVec_hitReq_3_82 = _GEN_302;
  wire         _GEN_303 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h12;
  wire         compressDataVec_hitReq_4_18;
  assign compressDataVec_hitReq_4_18 = _GEN_303;
  wire         compressDataVec_hitReq_4_82;
  assign compressDataVec_hitReq_4_82 = _GEN_303;
  wire         _GEN_304 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h12;
  wire         compressDataVec_hitReq_5_18;
  assign compressDataVec_hitReq_5_18 = _GEN_304;
  wire         compressDataVec_hitReq_5_82;
  assign compressDataVec_hitReq_5_82 = _GEN_304;
  wire         _GEN_305 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h12;
  wire         compressDataVec_hitReq_6_18;
  assign compressDataVec_hitReq_6_18 = _GEN_305;
  wire         compressDataVec_hitReq_6_82;
  assign compressDataVec_hitReq_6_82 = _GEN_305;
  wire         _GEN_306 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h12;
  wire         compressDataVec_hitReq_7_18;
  assign compressDataVec_hitReq_7_18 = _GEN_306;
  wire         compressDataVec_hitReq_7_82;
  assign compressDataVec_hitReq_7_82 = _GEN_306;
  wire         _GEN_307 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h12;
  wire         compressDataVec_hitReq_8_18;
  assign compressDataVec_hitReq_8_18 = _GEN_307;
  wire         compressDataVec_hitReq_8_82;
  assign compressDataVec_hitReq_8_82 = _GEN_307;
  wire         _GEN_308 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h12;
  wire         compressDataVec_hitReq_9_18;
  assign compressDataVec_hitReq_9_18 = _GEN_308;
  wire         compressDataVec_hitReq_9_82;
  assign compressDataVec_hitReq_9_82 = _GEN_308;
  wire         _GEN_309 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h12;
  wire         compressDataVec_hitReq_10_18;
  assign compressDataVec_hitReq_10_18 = _GEN_309;
  wire         compressDataVec_hitReq_10_82;
  assign compressDataVec_hitReq_10_82 = _GEN_309;
  wire         _GEN_310 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h12;
  wire         compressDataVec_hitReq_11_18;
  assign compressDataVec_hitReq_11_18 = _GEN_310;
  wire         compressDataVec_hitReq_11_82;
  assign compressDataVec_hitReq_11_82 = _GEN_310;
  wire         _GEN_311 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h12;
  wire         compressDataVec_hitReq_12_18;
  assign compressDataVec_hitReq_12_18 = _GEN_311;
  wire         compressDataVec_hitReq_12_82;
  assign compressDataVec_hitReq_12_82 = _GEN_311;
  wire         _GEN_312 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h12;
  wire         compressDataVec_hitReq_13_18;
  assign compressDataVec_hitReq_13_18 = _GEN_312;
  wire         compressDataVec_hitReq_13_82;
  assign compressDataVec_hitReq_13_82 = _GEN_312;
  wire         _GEN_313 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h12;
  wire         compressDataVec_hitReq_14_18;
  assign compressDataVec_hitReq_14_18 = _GEN_313;
  wire         compressDataVec_hitReq_14_82;
  assign compressDataVec_hitReq_14_82 = _GEN_313;
  wire         _GEN_314 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h12;
  wire         compressDataVec_hitReq_15_18;
  assign compressDataVec_hitReq_15_18 = _GEN_314;
  wire         compressDataVec_hitReq_15_82;
  assign compressDataVec_hitReq_15_82 = _GEN_314;
  wire         compressDataVec_hitReq_16_18 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h12;
  wire         compressDataVec_hitReq_17_18 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h12;
  wire         compressDataVec_hitReq_18_18 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h12;
  wire         compressDataVec_hitReq_19_18 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h12;
  wire         compressDataVec_hitReq_20_18 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h12;
  wire         compressDataVec_hitReq_21_18 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h12;
  wire         compressDataVec_hitReq_22_18 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h12;
  wire         compressDataVec_hitReq_23_18 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h12;
  wire         compressDataVec_hitReq_24_18 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h12;
  wire         compressDataVec_hitReq_25_18 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h12;
  wire         compressDataVec_hitReq_26_18 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h12;
  wire         compressDataVec_hitReq_27_18 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h12;
  wire         compressDataVec_hitReq_28_18 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h12;
  wire         compressDataVec_hitReq_29_18 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h12;
  wire         compressDataVec_hitReq_30_18 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h12;
  wire         compressDataVec_hitReq_31_18 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h12;
  wire [7:0]   compressDataVec_selectReqData_18 =
    (compressDataVec_hitReq_0_18 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_18 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_18 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_18 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_18 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_18 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_18 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_18 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_18 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_18 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_18 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_18 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_18 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_18 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_18 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_18 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_18 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_18 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_18 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_18 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_18 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_18 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_18 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_18 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_18 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_18 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_18 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_18 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_18 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_18 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_18 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_18 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_18 = tailCount > 5'h12;
  wire         _GEN_315 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h13;
  wire         compressDataVec_hitReq_0_19;
  assign compressDataVec_hitReq_0_19 = _GEN_315;
  wire         compressDataVec_hitReq_0_83;
  assign compressDataVec_hitReq_0_83 = _GEN_315;
  wire         _GEN_316 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h13;
  wire         compressDataVec_hitReq_1_19;
  assign compressDataVec_hitReq_1_19 = _GEN_316;
  wire         compressDataVec_hitReq_1_83;
  assign compressDataVec_hitReq_1_83 = _GEN_316;
  wire         _GEN_317 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h13;
  wire         compressDataVec_hitReq_2_19;
  assign compressDataVec_hitReq_2_19 = _GEN_317;
  wire         compressDataVec_hitReq_2_83;
  assign compressDataVec_hitReq_2_83 = _GEN_317;
  wire         _GEN_318 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h13;
  wire         compressDataVec_hitReq_3_19;
  assign compressDataVec_hitReq_3_19 = _GEN_318;
  wire         compressDataVec_hitReq_3_83;
  assign compressDataVec_hitReq_3_83 = _GEN_318;
  wire         _GEN_319 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h13;
  wire         compressDataVec_hitReq_4_19;
  assign compressDataVec_hitReq_4_19 = _GEN_319;
  wire         compressDataVec_hitReq_4_83;
  assign compressDataVec_hitReq_4_83 = _GEN_319;
  wire         _GEN_320 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h13;
  wire         compressDataVec_hitReq_5_19;
  assign compressDataVec_hitReq_5_19 = _GEN_320;
  wire         compressDataVec_hitReq_5_83;
  assign compressDataVec_hitReq_5_83 = _GEN_320;
  wire         _GEN_321 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h13;
  wire         compressDataVec_hitReq_6_19;
  assign compressDataVec_hitReq_6_19 = _GEN_321;
  wire         compressDataVec_hitReq_6_83;
  assign compressDataVec_hitReq_6_83 = _GEN_321;
  wire         _GEN_322 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h13;
  wire         compressDataVec_hitReq_7_19;
  assign compressDataVec_hitReq_7_19 = _GEN_322;
  wire         compressDataVec_hitReq_7_83;
  assign compressDataVec_hitReq_7_83 = _GEN_322;
  wire         _GEN_323 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h13;
  wire         compressDataVec_hitReq_8_19;
  assign compressDataVec_hitReq_8_19 = _GEN_323;
  wire         compressDataVec_hitReq_8_83;
  assign compressDataVec_hitReq_8_83 = _GEN_323;
  wire         _GEN_324 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h13;
  wire         compressDataVec_hitReq_9_19;
  assign compressDataVec_hitReq_9_19 = _GEN_324;
  wire         compressDataVec_hitReq_9_83;
  assign compressDataVec_hitReq_9_83 = _GEN_324;
  wire         _GEN_325 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h13;
  wire         compressDataVec_hitReq_10_19;
  assign compressDataVec_hitReq_10_19 = _GEN_325;
  wire         compressDataVec_hitReq_10_83;
  assign compressDataVec_hitReq_10_83 = _GEN_325;
  wire         _GEN_326 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h13;
  wire         compressDataVec_hitReq_11_19;
  assign compressDataVec_hitReq_11_19 = _GEN_326;
  wire         compressDataVec_hitReq_11_83;
  assign compressDataVec_hitReq_11_83 = _GEN_326;
  wire         _GEN_327 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h13;
  wire         compressDataVec_hitReq_12_19;
  assign compressDataVec_hitReq_12_19 = _GEN_327;
  wire         compressDataVec_hitReq_12_83;
  assign compressDataVec_hitReq_12_83 = _GEN_327;
  wire         _GEN_328 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h13;
  wire         compressDataVec_hitReq_13_19;
  assign compressDataVec_hitReq_13_19 = _GEN_328;
  wire         compressDataVec_hitReq_13_83;
  assign compressDataVec_hitReq_13_83 = _GEN_328;
  wire         _GEN_329 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h13;
  wire         compressDataVec_hitReq_14_19;
  assign compressDataVec_hitReq_14_19 = _GEN_329;
  wire         compressDataVec_hitReq_14_83;
  assign compressDataVec_hitReq_14_83 = _GEN_329;
  wire         _GEN_330 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h13;
  wire         compressDataVec_hitReq_15_19;
  assign compressDataVec_hitReq_15_19 = _GEN_330;
  wire         compressDataVec_hitReq_15_83;
  assign compressDataVec_hitReq_15_83 = _GEN_330;
  wire         compressDataVec_hitReq_16_19 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h13;
  wire         compressDataVec_hitReq_17_19 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h13;
  wire         compressDataVec_hitReq_18_19 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h13;
  wire         compressDataVec_hitReq_19_19 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h13;
  wire         compressDataVec_hitReq_20_19 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h13;
  wire         compressDataVec_hitReq_21_19 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h13;
  wire         compressDataVec_hitReq_22_19 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h13;
  wire         compressDataVec_hitReq_23_19 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h13;
  wire         compressDataVec_hitReq_24_19 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h13;
  wire         compressDataVec_hitReq_25_19 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h13;
  wire         compressDataVec_hitReq_26_19 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h13;
  wire         compressDataVec_hitReq_27_19 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h13;
  wire         compressDataVec_hitReq_28_19 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h13;
  wire         compressDataVec_hitReq_29_19 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h13;
  wire         compressDataVec_hitReq_30_19 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h13;
  wire         compressDataVec_hitReq_31_19 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h13;
  wire [7:0]   compressDataVec_selectReqData_19 =
    (compressDataVec_hitReq_0_19 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_19 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_19 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_19 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_19 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_19 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_19 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_19 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_19 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_19 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_19 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_19 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_19 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_19 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_19 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_19 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_19 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_19 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_19 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_19 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_19 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_19 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_19 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_19 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_19 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_19 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_19 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_19 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_19 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_19 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_19 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_19 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_19 = tailCount > 5'h13;
  wire         _GEN_331 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h14;
  wire         compressDataVec_hitReq_0_20;
  assign compressDataVec_hitReq_0_20 = _GEN_331;
  wire         compressDataVec_hitReq_0_84;
  assign compressDataVec_hitReq_0_84 = _GEN_331;
  wire         _GEN_332 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h14;
  wire         compressDataVec_hitReq_1_20;
  assign compressDataVec_hitReq_1_20 = _GEN_332;
  wire         compressDataVec_hitReq_1_84;
  assign compressDataVec_hitReq_1_84 = _GEN_332;
  wire         _GEN_333 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h14;
  wire         compressDataVec_hitReq_2_20;
  assign compressDataVec_hitReq_2_20 = _GEN_333;
  wire         compressDataVec_hitReq_2_84;
  assign compressDataVec_hitReq_2_84 = _GEN_333;
  wire         _GEN_334 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h14;
  wire         compressDataVec_hitReq_3_20;
  assign compressDataVec_hitReq_3_20 = _GEN_334;
  wire         compressDataVec_hitReq_3_84;
  assign compressDataVec_hitReq_3_84 = _GEN_334;
  wire         _GEN_335 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h14;
  wire         compressDataVec_hitReq_4_20;
  assign compressDataVec_hitReq_4_20 = _GEN_335;
  wire         compressDataVec_hitReq_4_84;
  assign compressDataVec_hitReq_4_84 = _GEN_335;
  wire         _GEN_336 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h14;
  wire         compressDataVec_hitReq_5_20;
  assign compressDataVec_hitReq_5_20 = _GEN_336;
  wire         compressDataVec_hitReq_5_84;
  assign compressDataVec_hitReq_5_84 = _GEN_336;
  wire         _GEN_337 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h14;
  wire         compressDataVec_hitReq_6_20;
  assign compressDataVec_hitReq_6_20 = _GEN_337;
  wire         compressDataVec_hitReq_6_84;
  assign compressDataVec_hitReq_6_84 = _GEN_337;
  wire         _GEN_338 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h14;
  wire         compressDataVec_hitReq_7_20;
  assign compressDataVec_hitReq_7_20 = _GEN_338;
  wire         compressDataVec_hitReq_7_84;
  assign compressDataVec_hitReq_7_84 = _GEN_338;
  wire         _GEN_339 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h14;
  wire         compressDataVec_hitReq_8_20;
  assign compressDataVec_hitReq_8_20 = _GEN_339;
  wire         compressDataVec_hitReq_8_84;
  assign compressDataVec_hitReq_8_84 = _GEN_339;
  wire         _GEN_340 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h14;
  wire         compressDataVec_hitReq_9_20;
  assign compressDataVec_hitReq_9_20 = _GEN_340;
  wire         compressDataVec_hitReq_9_84;
  assign compressDataVec_hitReq_9_84 = _GEN_340;
  wire         _GEN_341 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h14;
  wire         compressDataVec_hitReq_10_20;
  assign compressDataVec_hitReq_10_20 = _GEN_341;
  wire         compressDataVec_hitReq_10_84;
  assign compressDataVec_hitReq_10_84 = _GEN_341;
  wire         _GEN_342 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h14;
  wire         compressDataVec_hitReq_11_20;
  assign compressDataVec_hitReq_11_20 = _GEN_342;
  wire         compressDataVec_hitReq_11_84;
  assign compressDataVec_hitReq_11_84 = _GEN_342;
  wire         _GEN_343 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h14;
  wire         compressDataVec_hitReq_12_20;
  assign compressDataVec_hitReq_12_20 = _GEN_343;
  wire         compressDataVec_hitReq_12_84;
  assign compressDataVec_hitReq_12_84 = _GEN_343;
  wire         _GEN_344 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h14;
  wire         compressDataVec_hitReq_13_20;
  assign compressDataVec_hitReq_13_20 = _GEN_344;
  wire         compressDataVec_hitReq_13_84;
  assign compressDataVec_hitReq_13_84 = _GEN_344;
  wire         _GEN_345 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h14;
  wire         compressDataVec_hitReq_14_20;
  assign compressDataVec_hitReq_14_20 = _GEN_345;
  wire         compressDataVec_hitReq_14_84;
  assign compressDataVec_hitReq_14_84 = _GEN_345;
  wire         _GEN_346 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h14;
  wire         compressDataVec_hitReq_15_20;
  assign compressDataVec_hitReq_15_20 = _GEN_346;
  wire         compressDataVec_hitReq_15_84;
  assign compressDataVec_hitReq_15_84 = _GEN_346;
  wire         compressDataVec_hitReq_16_20 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h14;
  wire         compressDataVec_hitReq_17_20 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h14;
  wire         compressDataVec_hitReq_18_20 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h14;
  wire         compressDataVec_hitReq_19_20 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h14;
  wire         compressDataVec_hitReq_20_20 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h14;
  wire         compressDataVec_hitReq_21_20 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h14;
  wire         compressDataVec_hitReq_22_20 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h14;
  wire         compressDataVec_hitReq_23_20 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h14;
  wire         compressDataVec_hitReq_24_20 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h14;
  wire         compressDataVec_hitReq_25_20 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h14;
  wire         compressDataVec_hitReq_26_20 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h14;
  wire         compressDataVec_hitReq_27_20 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h14;
  wire         compressDataVec_hitReq_28_20 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h14;
  wire         compressDataVec_hitReq_29_20 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h14;
  wire         compressDataVec_hitReq_30_20 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h14;
  wire         compressDataVec_hitReq_31_20 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h14;
  wire [7:0]   compressDataVec_selectReqData_20 =
    (compressDataVec_hitReq_0_20 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_20 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_20 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_20 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_20 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_20 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_20 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_20 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_20 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_20 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_20 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_20 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_20 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_20 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_20 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_20 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_20 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_20 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_20 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_20 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_20 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_20 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_20 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_20 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_20 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_20 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_20 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_20 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_20 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_20 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_20 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_20 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_20 = tailCount > 5'h14;
  wire         _GEN_347 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h15;
  wire         compressDataVec_hitReq_0_21;
  assign compressDataVec_hitReq_0_21 = _GEN_347;
  wire         compressDataVec_hitReq_0_85;
  assign compressDataVec_hitReq_0_85 = _GEN_347;
  wire         _GEN_348 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h15;
  wire         compressDataVec_hitReq_1_21;
  assign compressDataVec_hitReq_1_21 = _GEN_348;
  wire         compressDataVec_hitReq_1_85;
  assign compressDataVec_hitReq_1_85 = _GEN_348;
  wire         _GEN_349 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h15;
  wire         compressDataVec_hitReq_2_21;
  assign compressDataVec_hitReq_2_21 = _GEN_349;
  wire         compressDataVec_hitReq_2_85;
  assign compressDataVec_hitReq_2_85 = _GEN_349;
  wire         _GEN_350 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h15;
  wire         compressDataVec_hitReq_3_21;
  assign compressDataVec_hitReq_3_21 = _GEN_350;
  wire         compressDataVec_hitReq_3_85;
  assign compressDataVec_hitReq_3_85 = _GEN_350;
  wire         _GEN_351 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h15;
  wire         compressDataVec_hitReq_4_21;
  assign compressDataVec_hitReq_4_21 = _GEN_351;
  wire         compressDataVec_hitReq_4_85;
  assign compressDataVec_hitReq_4_85 = _GEN_351;
  wire         _GEN_352 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h15;
  wire         compressDataVec_hitReq_5_21;
  assign compressDataVec_hitReq_5_21 = _GEN_352;
  wire         compressDataVec_hitReq_5_85;
  assign compressDataVec_hitReq_5_85 = _GEN_352;
  wire         _GEN_353 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h15;
  wire         compressDataVec_hitReq_6_21;
  assign compressDataVec_hitReq_6_21 = _GEN_353;
  wire         compressDataVec_hitReq_6_85;
  assign compressDataVec_hitReq_6_85 = _GEN_353;
  wire         _GEN_354 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h15;
  wire         compressDataVec_hitReq_7_21;
  assign compressDataVec_hitReq_7_21 = _GEN_354;
  wire         compressDataVec_hitReq_7_85;
  assign compressDataVec_hitReq_7_85 = _GEN_354;
  wire         _GEN_355 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h15;
  wire         compressDataVec_hitReq_8_21;
  assign compressDataVec_hitReq_8_21 = _GEN_355;
  wire         compressDataVec_hitReq_8_85;
  assign compressDataVec_hitReq_8_85 = _GEN_355;
  wire         _GEN_356 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h15;
  wire         compressDataVec_hitReq_9_21;
  assign compressDataVec_hitReq_9_21 = _GEN_356;
  wire         compressDataVec_hitReq_9_85;
  assign compressDataVec_hitReq_9_85 = _GEN_356;
  wire         _GEN_357 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h15;
  wire         compressDataVec_hitReq_10_21;
  assign compressDataVec_hitReq_10_21 = _GEN_357;
  wire         compressDataVec_hitReq_10_85;
  assign compressDataVec_hitReq_10_85 = _GEN_357;
  wire         _GEN_358 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h15;
  wire         compressDataVec_hitReq_11_21;
  assign compressDataVec_hitReq_11_21 = _GEN_358;
  wire         compressDataVec_hitReq_11_85;
  assign compressDataVec_hitReq_11_85 = _GEN_358;
  wire         _GEN_359 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h15;
  wire         compressDataVec_hitReq_12_21;
  assign compressDataVec_hitReq_12_21 = _GEN_359;
  wire         compressDataVec_hitReq_12_85;
  assign compressDataVec_hitReq_12_85 = _GEN_359;
  wire         _GEN_360 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h15;
  wire         compressDataVec_hitReq_13_21;
  assign compressDataVec_hitReq_13_21 = _GEN_360;
  wire         compressDataVec_hitReq_13_85;
  assign compressDataVec_hitReq_13_85 = _GEN_360;
  wire         _GEN_361 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h15;
  wire         compressDataVec_hitReq_14_21;
  assign compressDataVec_hitReq_14_21 = _GEN_361;
  wire         compressDataVec_hitReq_14_85;
  assign compressDataVec_hitReq_14_85 = _GEN_361;
  wire         _GEN_362 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h15;
  wire         compressDataVec_hitReq_15_21;
  assign compressDataVec_hitReq_15_21 = _GEN_362;
  wire         compressDataVec_hitReq_15_85;
  assign compressDataVec_hitReq_15_85 = _GEN_362;
  wire         compressDataVec_hitReq_16_21 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h15;
  wire         compressDataVec_hitReq_17_21 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h15;
  wire         compressDataVec_hitReq_18_21 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h15;
  wire         compressDataVec_hitReq_19_21 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h15;
  wire         compressDataVec_hitReq_20_21 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h15;
  wire         compressDataVec_hitReq_21_21 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h15;
  wire         compressDataVec_hitReq_22_21 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h15;
  wire         compressDataVec_hitReq_23_21 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h15;
  wire         compressDataVec_hitReq_24_21 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h15;
  wire         compressDataVec_hitReq_25_21 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h15;
  wire         compressDataVec_hitReq_26_21 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h15;
  wire         compressDataVec_hitReq_27_21 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h15;
  wire         compressDataVec_hitReq_28_21 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h15;
  wire         compressDataVec_hitReq_29_21 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h15;
  wire         compressDataVec_hitReq_30_21 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h15;
  wire         compressDataVec_hitReq_31_21 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h15;
  wire [7:0]   compressDataVec_selectReqData_21 =
    (compressDataVec_hitReq_0_21 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_21 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_21 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_21 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_21 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_21 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_21 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_21 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_21 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_21 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_21 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_21 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_21 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_21 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_21 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_21 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_21 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_21 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_21 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_21 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_21 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_21 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_21 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_21 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_21 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_21 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_21 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_21 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_21 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_21 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_21 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_21 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_21 = tailCount > 5'h15;
  wire         _GEN_363 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h16;
  wire         compressDataVec_hitReq_0_22;
  assign compressDataVec_hitReq_0_22 = _GEN_363;
  wire         compressDataVec_hitReq_0_86;
  assign compressDataVec_hitReq_0_86 = _GEN_363;
  wire         _GEN_364 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h16;
  wire         compressDataVec_hitReq_1_22;
  assign compressDataVec_hitReq_1_22 = _GEN_364;
  wire         compressDataVec_hitReq_1_86;
  assign compressDataVec_hitReq_1_86 = _GEN_364;
  wire         _GEN_365 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h16;
  wire         compressDataVec_hitReq_2_22;
  assign compressDataVec_hitReq_2_22 = _GEN_365;
  wire         compressDataVec_hitReq_2_86;
  assign compressDataVec_hitReq_2_86 = _GEN_365;
  wire         _GEN_366 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h16;
  wire         compressDataVec_hitReq_3_22;
  assign compressDataVec_hitReq_3_22 = _GEN_366;
  wire         compressDataVec_hitReq_3_86;
  assign compressDataVec_hitReq_3_86 = _GEN_366;
  wire         _GEN_367 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h16;
  wire         compressDataVec_hitReq_4_22;
  assign compressDataVec_hitReq_4_22 = _GEN_367;
  wire         compressDataVec_hitReq_4_86;
  assign compressDataVec_hitReq_4_86 = _GEN_367;
  wire         _GEN_368 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h16;
  wire         compressDataVec_hitReq_5_22;
  assign compressDataVec_hitReq_5_22 = _GEN_368;
  wire         compressDataVec_hitReq_5_86;
  assign compressDataVec_hitReq_5_86 = _GEN_368;
  wire         _GEN_369 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h16;
  wire         compressDataVec_hitReq_6_22;
  assign compressDataVec_hitReq_6_22 = _GEN_369;
  wire         compressDataVec_hitReq_6_86;
  assign compressDataVec_hitReq_6_86 = _GEN_369;
  wire         _GEN_370 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h16;
  wire         compressDataVec_hitReq_7_22;
  assign compressDataVec_hitReq_7_22 = _GEN_370;
  wire         compressDataVec_hitReq_7_86;
  assign compressDataVec_hitReq_7_86 = _GEN_370;
  wire         _GEN_371 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h16;
  wire         compressDataVec_hitReq_8_22;
  assign compressDataVec_hitReq_8_22 = _GEN_371;
  wire         compressDataVec_hitReq_8_86;
  assign compressDataVec_hitReq_8_86 = _GEN_371;
  wire         _GEN_372 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h16;
  wire         compressDataVec_hitReq_9_22;
  assign compressDataVec_hitReq_9_22 = _GEN_372;
  wire         compressDataVec_hitReq_9_86;
  assign compressDataVec_hitReq_9_86 = _GEN_372;
  wire         _GEN_373 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h16;
  wire         compressDataVec_hitReq_10_22;
  assign compressDataVec_hitReq_10_22 = _GEN_373;
  wire         compressDataVec_hitReq_10_86;
  assign compressDataVec_hitReq_10_86 = _GEN_373;
  wire         _GEN_374 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h16;
  wire         compressDataVec_hitReq_11_22;
  assign compressDataVec_hitReq_11_22 = _GEN_374;
  wire         compressDataVec_hitReq_11_86;
  assign compressDataVec_hitReq_11_86 = _GEN_374;
  wire         _GEN_375 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h16;
  wire         compressDataVec_hitReq_12_22;
  assign compressDataVec_hitReq_12_22 = _GEN_375;
  wire         compressDataVec_hitReq_12_86;
  assign compressDataVec_hitReq_12_86 = _GEN_375;
  wire         _GEN_376 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h16;
  wire         compressDataVec_hitReq_13_22;
  assign compressDataVec_hitReq_13_22 = _GEN_376;
  wire         compressDataVec_hitReq_13_86;
  assign compressDataVec_hitReq_13_86 = _GEN_376;
  wire         _GEN_377 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h16;
  wire         compressDataVec_hitReq_14_22;
  assign compressDataVec_hitReq_14_22 = _GEN_377;
  wire         compressDataVec_hitReq_14_86;
  assign compressDataVec_hitReq_14_86 = _GEN_377;
  wire         _GEN_378 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h16;
  wire         compressDataVec_hitReq_15_22;
  assign compressDataVec_hitReq_15_22 = _GEN_378;
  wire         compressDataVec_hitReq_15_86;
  assign compressDataVec_hitReq_15_86 = _GEN_378;
  wire         compressDataVec_hitReq_16_22 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h16;
  wire         compressDataVec_hitReq_17_22 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h16;
  wire         compressDataVec_hitReq_18_22 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h16;
  wire         compressDataVec_hitReq_19_22 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h16;
  wire         compressDataVec_hitReq_20_22 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h16;
  wire         compressDataVec_hitReq_21_22 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h16;
  wire         compressDataVec_hitReq_22_22 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h16;
  wire         compressDataVec_hitReq_23_22 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h16;
  wire         compressDataVec_hitReq_24_22 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h16;
  wire         compressDataVec_hitReq_25_22 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h16;
  wire         compressDataVec_hitReq_26_22 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h16;
  wire         compressDataVec_hitReq_27_22 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h16;
  wire         compressDataVec_hitReq_28_22 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h16;
  wire         compressDataVec_hitReq_29_22 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h16;
  wire         compressDataVec_hitReq_30_22 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h16;
  wire         compressDataVec_hitReq_31_22 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h16;
  wire [7:0]   compressDataVec_selectReqData_22 =
    (compressDataVec_hitReq_0_22 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_22 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_22 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_22 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_22 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_22 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_22 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_22 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_22 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_22 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_22 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_22 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_22 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_22 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_22 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_22 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_22 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_22 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_22 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_22 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_22 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_22 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_22 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_22 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_22 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_22 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_22 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_22 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_22 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_22 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_22 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_22 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_22 = tailCount > 5'h16;
  wire         _GEN_379 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h17;
  wire         compressDataVec_hitReq_0_23;
  assign compressDataVec_hitReq_0_23 = _GEN_379;
  wire         compressDataVec_hitReq_0_87;
  assign compressDataVec_hitReq_0_87 = _GEN_379;
  wire         _GEN_380 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h17;
  wire         compressDataVec_hitReq_1_23;
  assign compressDataVec_hitReq_1_23 = _GEN_380;
  wire         compressDataVec_hitReq_1_87;
  assign compressDataVec_hitReq_1_87 = _GEN_380;
  wire         _GEN_381 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h17;
  wire         compressDataVec_hitReq_2_23;
  assign compressDataVec_hitReq_2_23 = _GEN_381;
  wire         compressDataVec_hitReq_2_87;
  assign compressDataVec_hitReq_2_87 = _GEN_381;
  wire         _GEN_382 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h17;
  wire         compressDataVec_hitReq_3_23;
  assign compressDataVec_hitReq_3_23 = _GEN_382;
  wire         compressDataVec_hitReq_3_87;
  assign compressDataVec_hitReq_3_87 = _GEN_382;
  wire         _GEN_383 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h17;
  wire         compressDataVec_hitReq_4_23;
  assign compressDataVec_hitReq_4_23 = _GEN_383;
  wire         compressDataVec_hitReq_4_87;
  assign compressDataVec_hitReq_4_87 = _GEN_383;
  wire         _GEN_384 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h17;
  wire         compressDataVec_hitReq_5_23;
  assign compressDataVec_hitReq_5_23 = _GEN_384;
  wire         compressDataVec_hitReq_5_87;
  assign compressDataVec_hitReq_5_87 = _GEN_384;
  wire         _GEN_385 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h17;
  wire         compressDataVec_hitReq_6_23;
  assign compressDataVec_hitReq_6_23 = _GEN_385;
  wire         compressDataVec_hitReq_6_87;
  assign compressDataVec_hitReq_6_87 = _GEN_385;
  wire         _GEN_386 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h17;
  wire         compressDataVec_hitReq_7_23;
  assign compressDataVec_hitReq_7_23 = _GEN_386;
  wire         compressDataVec_hitReq_7_87;
  assign compressDataVec_hitReq_7_87 = _GEN_386;
  wire         _GEN_387 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h17;
  wire         compressDataVec_hitReq_8_23;
  assign compressDataVec_hitReq_8_23 = _GEN_387;
  wire         compressDataVec_hitReq_8_87;
  assign compressDataVec_hitReq_8_87 = _GEN_387;
  wire         _GEN_388 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h17;
  wire         compressDataVec_hitReq_9_23;
  assign compressDataVec_hitReq_9_23 = _GEN_388;
  wire         compressDataVec_hitReq_9_87;
  assign compressDataVec_hitReq_9_87 = _GEN_388;
  wire         _GEN_389 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h17;
  wire         compressDataVec_hitReq_10_23;
  assign compressDataVec_hitReq_10_23 = _GEN_389;
  wire         compressDataVec_hitReq_10_87;
  assign compressDataVec_hitReq_10_87 = _GEN_389;
  wire         _GEN_390 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h17;
  wire         compressDataVec_hitReq_11_23;
  assign compressDataVec_hitReq_11_23 = _GEN_390;
  wire         compressDataVec_hitReq_11_87;
  assign compressDataVec_hitReq_11_87 = _GEN_390;
  wire         _GEN_391 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h17;
  wire         compressDataVec_hitReq_12_23;
  assign compressDataVec_hitReq_12_23 = _GEN_391;
  wire         compressDataVec_hitReq_12_87;
  assign compressDataVec_hitReq_12_87 = _GEN_391;
  wire         _GEN_392 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h17;
  wire         compressDataVec_hitReq_13_23;
  assign compressDataVec_hitReq_13_23 = _GEN_392;
  wire         compressDataVec_hitReq_13_87;
  assign compressDataVec_hitReq_13_87 = _GEN_392;
  wire         _GEN_393 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h17;
  wire         compressDataVec_hitReq_14_23;
  assign compressDataVec_hitReq_14_23 = _GEN_393;
  wire         compressDataVec_hitReq_14_87;
  assign compressDataVec_hitReq_14_87 = _GEN_393;
  wire         _GEN_394 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h17;
  wire         compressDataVec_hitReq_15_23;
  assign compressDataVec_hitReq_15_23 = _GEN_394;
  wire         compressDataVec_hitReq_15_87;
  assign compressDataVec_hitReq_15_87 = _GEN_394;
  wire         compressDataVec_hitReq_16_23 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h17;
  wire         compressDataVec_hitReq_17_23 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h17;
  wire         compressDataVec_hitReq_18_23 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h17;
  wire         compressDataVec_hitReq_19_23 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h17;
  wire         compressDataVec_hitReq_20_23 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h17;
  wire         compressDataVec_hitReq_21_23 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h17;
  wire         compressDataVec_hitReq_22_23 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h17;
  wire         compressDataVec_hitReq_23_23 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h17;
  wire         compressDataVec_hitReq_24_23 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h17;
  wire         compressDataVec_hitReq_25_23 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h17;
  wire         compressDataVec_hitReq_26_23 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h17;
  wire         compressDataVec_hitReq_27_23 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h17;
  wire         compressDataVec_hitReq_28_23 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h17;
  wire         compressDataVec_hitReq_29_23 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h17;
  wire         compressDataVec_hitReq_30_23 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h17;
  wire         compressDataVec_hitReq_31_23 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h17;
  wire [7:0]   compressDataVec_selectReqData_23 =
    (compressDataVec_hitReq_0_23 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_23 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_23 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_23 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_23 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_23 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_23 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_23 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_23 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_23 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_23 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_23 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_23 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_23 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_23 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_23 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_23 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_23 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_23 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_23 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_23 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_23 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_23 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_23 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_23 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_23 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_23 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_23 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_23 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_23 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_23 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_23 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_23 = tailCount > 5'h17;
  wire         _GEN_395 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h18;
  wire         compressDataVec_hitReq_0_24;
  assign compressDataVec_hitReq_0_24 = _GEN_395;
  wire         compressDataVec_hitReq_0_88;
  assign compressDataVec_hitReq_0_88 = _GEN_395;
  wire         _GEN_396 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h18;
  wire         compressDataVec_hitReq_1_24;
  assign compressDataVec_hitReq_1_24 = _GEN_396;
  wire         compressDataVec_hitReq_1_88;
  assign compressDataVec_hitReq_1_88 = _GEN_396;
  wire         _GEN_397 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h18;
  wire         compressDataVec_hitReq_2_24;
  assign compressDataVec_hitReq_2_24 = _GEN_397;
  wire         compressDataVec_hitReq_2_88;
  assign compressDataVec_hitReq_2_88 = _GEN_397;
  wire         _GEN_398 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h18;
  wire         compressDataVec_hitReq_3_24;
  assign compressDataVec_hitReq_3_24 = _GEN_398;
  wire         compressDataVec_hitReq_3_88;
  assign compressDataVec_hitReq_3_88 = _GEN_398;
  wire         _GEN_399 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h18;
  wire         compressDataVec_hitReq_4_24;
  assign compressDataVec_hitReq_4_24 = _GEN_399;
  wire         compressDataVec_hitReq_4_88;
  assign compressDataVec_hitReq_4_88 = _GEN_399;
  wire         _GEN_400 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h18;
  wire         compressDataVec_hitReq_5_24;
  assign compressDataVec_hitReq_5_24 = _GEN_400;
  wire         compressDataVec_hitReq_5_88;
  assign compressDataVec_hitReq_5_88 = _GEN_400;
  wire         _GEN_401 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h18;
  wire         compressDataVec_hitReq_6_24;
  assign compressDataVec_hitReq_6_24 = _GEN_401;
  wire         compressDataVec_hitReq_6_88;
  assign compressDataVec_hitReq_6_88 = _GEN_401;
  wire         _GEN_402 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h18;
  wire         compressDataVec_hitReq_7_24;
  assign compressDataVec_hitReq_7_24 = _GEN_402;
  wire         compressDataVec_hitReq_7_88;
  assign compressDataVec_hitReq_7_88 = _GEN_402;
  wire         _GEN_403 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h18;
  wire         compressDataVec_hitReq_8_24;
  assign compressDataVec_hitReq_8_24 = _GEN_403;
  wire         compressDataVec_hitReq_8_88;
  assign compressDataVec_hitReq_8_88 = _GEN_403;
  wire         _GEN_404 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h18;
  wire         compressDataVec_hitReq_9_24;
  assign compressDataVec_hitReq_9_24 = _GEN_404;
  wire         compressDataVec_hitReq_9_88;
  assign compressDataVec_hitReq_9_88 = _GEN_404;
  wire         _GEN_405 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h18;
  wire         compressDataVec_hitReq_10_24;
  assign compressDataVec_hitReq_10_24 = _GEN_405;
  wire         compressDataVec_hitReq_10_88;
  assign compressDataVec_hitReq_10_88 = _GEN_405;
  wire         _GEN_406 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h18;
  wire         compressDataVec_hitReq_11_24;
  assign compressDataVec_hitReq_11_24 = _GEN_406;
  wire         compressDataVec_hitReq_11_88;
  assign compressDataVec_hitReq_11_88 = _GEN_406;
  wire         _GEN_407 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h18;
  wire         compressDataVec_hitReq_12_24;
  assign compressDataVec_hitReq_12_24 = _GEN_407;
  wire         compressDataVec_hitReq_12_88;
  assign compressDataVec_hitReq_12_88 = _GEN_407;
  wire         _GEN_408 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h18;
  wire         compressDataVec_hitReq_13_24;
  assign compressDataVec_hitReq_13_24 = _GEN_408;
  wire         compressDataVec_hitReq_13_88;
  assign compressDataVec_hitReq_13_88 = _GEN_408;
  wire         _GEN_409 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h18;
  wire         compressDataVec_hitReq_14_24;
  assign compressDataVec_hitReq_14_24 = _GEN_409;
  wire         compressDataVec_hitReq_14_88;
  assign compressDataVec_hitReq_14_88 = _GEN_409;
  wire         _GEN_410 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h18;
  wire         compressDataVec_hitReq_15_24;
  assign compressDataVec_hitReq_15_24 = _GEN_410;
  wire         compressDataVec_hitReq_15_88;
  assign compressDataVec_hitReq_15_88 = _GEN_410;
  wire         compressDataVec_hitReq_16_24 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h18;
  wire         compressDataVec_hitReq_17_24 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h18;
  wire         compressDataVec_hitReq_18_24 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h18;
  wire         compressDataVec_hitReq_19_24 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h18;
  wire         compressDataVec_hitReq_20_24 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h18;
  wire         compressDataVec_hitReq_21_24 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h18;
  wire         compressDataVec_hitReq_22_24 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h18;
  wire         compressDataVec_hitReq_23_24 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h18;
  wire         compressDataVec_hitReq_24_24 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h18;
  wire         compressDataVec_hitReq_25_24 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h18;
  wire         compressDataVec_hitReq_26_24 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h18;
  wire         compressDataVec_hitReq_27_24 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h18;
  wire         compressDataVec_hitReq_28_24 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h18;
  wire         compressDataVec_hitReq_29_24 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h18;
  wire         compressDataVec_hitReq_30_24 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h18;
  wire         compressDataVec_hitReq_31_24 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h18;
  wire [7:0]   compressDataVec_selectReqData_24 =
    (compressDataVec_hitReq_0_24 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_24 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_24 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_24 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_24 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_24 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_24 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_24 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_24 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_24 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_24 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_24 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_24 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_24 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_24 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_24 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_24 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_24 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_24 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_24 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_24 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_24 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_24 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_24 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_24 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_24 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_24 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_24 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_24 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_24 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_24 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_24 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_24 = tailCount > 5'h18;
  wire         _GEN_411 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h19;
  wire         compressDataVec_hitReq_0_25;
  assign compressDataVec_hitReq_0_25 = _GEN_411;
  wire         compressDataVec_hitReq_0_89;
  assign compressDataVec_hitReq_0_89 = _GEN_411;
  wire         _GEN_412 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h19;
  wire         compressDataVec_hitReq_1_25;
  assign compressDataVec_hitReq_1_25 = _GEN_412;
  wire         compressDataVec_hitReq_1_89;
  assign compressDataVec_hitReq_1_89 = _GEN_412;
  wire         _GEN_413 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h19;
  wire         compressDataVec_hitReq_2_25;
  assign compressDataVec_hitReq_2_25 = _GEN_413;
  wire         compressDataVec_hitReq_2_89;
  assign compressDataVec_hitReq_2_89 = _GEN_413;
  wire         _GEN_414 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h19;
  wire         compressDataVec_hitReq_3_25;
  assign compressDataVec_hitReq_3_25 = _GEN_414;
  wire         compressDataVec_hitReq_3_89;
  assign compressDataVec_hitReq_3_89 = _GEN_414;
  wire         _GEN_415 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h19;
  wire         compressDataVec_hitReq_4_25;
  assign compressDataVec_hitReq_4_25 = _GEN_415;
  wire         compressDataVec_hitReq_4_89;
  assign compressDataVec_hitReq_4_89 = _GEN_415;
  wire         _GEN_416 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h19;
  wire         compressDataVec_hitReq_5_25;
  assign compressDataVec_hitReq_5_25 = _GEN_416;
  wire         compressDataVec_hitReq_5_89;
  assign compressDataVec_hitReq_5_89 = _GEN_416;
  wire         _GEN_417 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h19;
  wire         compressDataVec_hitReq_6_25;
  assign compressDataVec_hitReq_6_25 = _GEN_417;
  wire         compressDataVec_hitReq_6_89;
  assign compressDataVec_hitReq_6_89 = _GEN_417;
  wire         _GEN_418 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h19;
  wire         compressDataVec_hitReq_7_25;
  assign compressDataVec_hitReq_7_25 = _GEN_418;
  wire         compressDataVec_hitReq_7_89;
  assign compressDataVec_hitReq_7_89 = _GEN_418;
  wire         _GEN_419 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h19;
  wire         compressDataVec_hitReq_8_25;
  assign compressDataVec_hitReq_8_25 = _GEN_419;
  wire         compressDataVec_hitReq_8_89;
  assign compressDataVec_hitReq_8_89 = _GEN_419;
  wire         _GEN_420 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h19;
  wire         compressDataVec_hitReq_9_25;
  assign compressDataVec_hitReq_9_25 = _GEN_420;
  wire         compressDataVec_hitReq_9_89;
  assign compressDataVec_hitReq_9_89 = _GEN_420;
  wire         _GEN_421 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h19;
  wire         compressDataVec_hitReq_10_25;
  assign compressDataVec_hitReq_10_25 = _GEN_421;
  wire         compressDataVec_hitReq_10_89;
  assign compressDataVec_hitReq_10_89 = _GEN_421;
  wire         _GEN_422 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h19;
  wire         compressDataVec_hitReq_11_25;
  assign compressDataVec_hitReq_11_25 = _GEN_422;
  wire         compressDataVec_hitReq_11_89;
  assign compressDataVec_hitReq_11_89 = _GEN_422;
  wire         _GEN_423 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h19;
  wire         compressDataVec_hitReq_12_25;
  assign compressDataVec_hitReq_12_25 = _GEN_423;
  wire         compressDataVec_hitReq_12_89;
  assign compressDataVec_hitReq_12_89 = _GEN_423;
  wire         _GEN_424 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h19;
  wire         compressDataVec_hitReq_13_25;
  assign compressDataVec_hitReq_13_25 = _GEN_424;
  wire         compressDataVec_hitReq_13_89;
  assign compressDataVec_hitReq_13_89 = _GEN_424;
  wire         _GEN_425 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h19;
  wire         compressDataVec_hitReq_14_25;
  assign compressDataVec_hitReq_14_25 = _GEN_425;
  wire         compressDataVec_hitReq_14_89;
  assign compressDataVec_hitReq_14_89 = _GEN_425;
  wire         _GEN_426 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h19;
  wire         compressDataVec_hitReq_15_25;
  assign compressDataVec_hitReq_15_25 = _GEN_426;
  wire         compressDataVec_hitReq_15_89;
  assign compressDataVec_hitReq_15_89 = _GEN_426;
  wire         compressDataVec_hitReq_16_25 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h19;
  wire         compressDataVec_hitReq_17_25 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h19;
  wire         compressDataVec_hitReq_18_25 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h19;
  wire         compressDataVec_hitReq_19_25 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h19;
  wire         compressDataVec_hitReq_20_25 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h19;
  wire         compressDataVec_hitReq_21_25 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h19;
  wire         compressDataVec_hitReq_22_25 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h19;
  wire         compressDataVec_hitReq_23_25 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h19;
  wire         compressDataVec_hitReq_24_25 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h19;
  wire         compressDataVec_hitReq_25_25 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h19;
  wire         compressDataVec_hitReq_26_25 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h19;
  wire         compressDataVec_hitReq_27_25 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h19;
  wire         compressDataVec_hitReq_28_25 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h19;
  wire         compressDataVec_hitReq_29_25 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h19;
  wire         compressDataVec_hitReq_30_25 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h19;
  wire         compressDataVec_hitReq_31_25 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h19;
  wire [7:0]   compressDataVec_selectReqData_25 =
    (compressDataVec_hitReq_0_25 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_25 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_25 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_25 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_25 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_25 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_25 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_25 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_25 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_25 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_25 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_25 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_25 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_25 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_25 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_25 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_25 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_25 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_25 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_25 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_25 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_25 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_25 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_25 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_25 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_25 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_25 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_25 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_25 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_25 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_25 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_25 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_25 = tailCount > 5'h19;
  wire         _GEN_427 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1A;
  wire         compressDataVec_hitReq_0_26;
  assign compressDataVec_hitReq_0_26 = _GEN_427;
  wire         compressDataVec_hitReq_0_90;
  assign compressDataVec_hitReq_0_90 = _GEN_427;
  wire         _GEN_428 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1A;
  wire         compressDataVec_hitReq_1_26;
  assign compressDataVec_hitReq_1_26 = _GEN_428;
  wire         compressDataVec_hitReq_1_90;
  assign compressDataVec_hitReq_1_90 = _GEN_428;
  wire         _GEN_429 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1A;
  wire         compressDataVec_hitReq_2_26;
  assign compressDataVec_hitReq_2_26 = _GEN_429;
  wire         compressDataVec_hitReq_2_90;
  assign compressDataVec_hitReq_2_90 = _GEN_429;
  wire         _GEN_430 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1A;
  wire         compressDataVec_hitReq_3_26;
  assign compressDataVec_hitReq_3_26 = _GEN_430;
  wire         compressDataVec_hitReq_3_90;
  assign compressDataVec_hitReq_3_90 = _GEN_430;
  wire         _GEN_431 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1A;
  wire         compressDataVec_hitReq_4_26;
  assign compressDataVec_hitReq_4_26 = _GEN_431;
  wire         compressDataVec_hitReq_4_90;
  assign compressDataVec_hitReq_4_90 = _GEN_431;
  wire         _GEN_432 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1A;
  wire         compressDataVec_hitReq_5_26;
  assign compressDataVec_hitReq_5_26 = _GEN_432;
  wire         compressDataVec_hitReq_5_90;
  assign compressDataVec_hitReq_5_90 = _GEN_432;
  wire         _GEN_433 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1A;
  wire         compressDataVec_hitReq_6_26;
  assign compressDataVec_hitReq_6_26 = _GEN_433;
  wire         compressDataVec_hitReq_6_90;
  assign compressDataVec_hitReq_6_90 = _GEN_433;
  wire         _GEN_434 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1A;
  wire         compressDataVec_hitReq_7_26;
  assign compressDataVec_hitReq_7_26 = _GEN_434;
  wire         compressDataVec_hitReq_7_90;
  assign compressDataVec_hitReq_7_90 = _GEN_434;
  wire         _GEN_435 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1A;
  wire         compressDataVec_hitReq_8_26;
  assign compressDataVec_hitReq_8_26 = _GEN_435;
  wire         compressDataVec_hitReq_8_90;
  assign compressDataVec_hitReq_8_90 = _GEN_435;
  wire         _GEN_436 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1A;
  wire         compressDataVec_hitReq_9_26;
  assign compressDataVec_hitReq_9_26 = _GEN_436;
  wire         compressDataVec_hitReq_9_90;
  assign compressDataVec_hitReq_9_90 = _GEN_436;
  wire         _GEN_437 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1A;
  wire         compressDataVec_hitReq_10_26;
  assign compressDataVec_hitReq_10_26 = _GEN_437;
  wire         compressDataVec_hitReq_10_90;
  assign compressDataVec_hitReq_10_90 = _GEN_437;
  wire         _GEN_438 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1A;
  wire         compressDataVec_hitReq_11_26;
  assign compressDataVec_hitReq_11_26 = _GEN_438;
  wire         compressDataVec_hitReq_11_90;
  assign compressDataVec_hitReq_11_90 = _GEN_438;
  wire         _GEN_439 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1A;
  wire         compressDataVec_hitReq_12_26;
  assign compressDataVec_hitReq_12_26 = _GEN_439;
  wire         compressDataVec_hitReq_12_90;
  assign compressDataVec_hitReq_12_90 = _GEN_439;
  wire         _GEN_440 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1A;
  wire         compressDataVec_hitReq_13_26;
  assign compressDataVec_hitReq_13_26 = _GEN_440;
  wire         compressDataVec_hitReq_13_90;
  assign compressDataVec_hitReq_13_90 = _GEN_440;
  wire         _GEN_441 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1A;
  wire         compressDataVec_hitReq_14_26;
  assign compressDataVec_hitReq_14_26 = _GEN_441;
  wire         compressDataVec_hitReq_14_90;
  assign compressDataVec_hitReq_14_90 = _GEN_441;
  wire         _GEN_442 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1A;
  wire         compressDataVec_hitReq_15_26;
  assign compressDataVec_hitReq_15_26 = _GEN_442;
  wire         compressDataVec_hitReq_15_90;
  assign compressDataVec_hitReq_15_90 = _GEN_442;
  wire         compressDataVec_hitReq_16_26 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1A;
  wire         compressDataVec_hitReq_17_26 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1A;
  wire         compressDataVec_hitReq_18_26 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1A;
  wire         compressDataVec_hitReq_19_26 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1A;
  wire         compressDataVec_hitReq_20_26 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1A;
  wire         compressDataVec_hitReq_21_26 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1A;
  wire         compressDataVec_hitReq_22_26 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1A;
  wire         compressDataVec_hitReq_23_26 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1A;
  wire         compressDataVec_hitReq_24_26 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1A;
  wire         compressDataVec_hitReq_25_26 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1A;
  wire         compressDataVec_hitReq_26_26 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1A;
  wire         compressDataVec_hitReq_27_26 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1A;
  wire         compressDataVec_hitReq_28_26 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1A;
  wire         compressDataVec_hitReq_29_26 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1A;
  wire         compressDataVec_hitReq_30_26 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1A;
  wire         compressDataVec_hitReq_31_26 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1A;
  wire [7:0]   compressDataVec_selectReqData_26 =
    (compressDataVec_hitReq_0_26 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_26 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_26 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_26 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_26 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_26 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_26 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_26 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_26 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_26 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_26 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_26 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_26 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_26 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_26 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_26 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_26 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_26 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_26 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_26 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_26 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_26 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_26 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_26 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_26 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_26 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_26 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_26 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_26 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_26 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_26 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_26 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_26 = tailCount > 5'h1A;
  wire         _GEN_443 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1B;
  wire         compressDataVec_hitReq_0_27;
  assign compressDataVec_hitReq_0_27 = _GEN_443;
  wire         compressDataVec_hitReq_0_91;
  assign compressDataVec_hitReq_0_91 = _GEN_443;
  wire         _GEN_444 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1B;
  wire         compressDataVec_hitReq_1_27;
  assign compressDataVec_hitReq_1_27 = _GEN_444;
  wire         compressDataVec_hitReq_1_91;
  assign compressDataVec_hitReq_1_91 = _GEN_444;
  wire         _GEN_445 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1B;
  wire         compressDataVec_hitReq_2_27;
  assign compressDataVec_hitReq_2_27 = _GEN_445;
  wire         compressDataVec_hitReq_2_91;
  assign compressDataVec_hitReq_2_91 = _GEN_445;
  wire         _GEN_446 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1B;
  wire         compressDataVec_hitReq_3_27;
  assign compressDataVec_hitReq_3_27 = _GEN_446;
  wire         compressDataVec_hitReq_3_91;
  assign compressDataVec_hitReq_3_91 = _GEN_446;
  wire         _GEN_447 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1B;
  wire         compressDataVec_hitReq_4_27;
  assign compressDataVec_hitReq_4_27 = _GEN_447;
  wire         compressDataVec_hitReq_4_91;
  assign compressDataVec_hitReq_4_91 = _GEN_447;
  wire         _GEN_448 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1B;
  wire         compressDataVec_hitReq_5_27;
  assign compressDataVec_hitReq_5_27 = _GEN_448;
  wire         compressDataVec_hitReq_5_91;
  assign compressDataVec_hitReq_5_91 = _GEN_448;
  wire         _GEN_449 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1B;
  wire         compressDataVec_hitReq_6_27;
  assign compressDataVec_hitReq_6_27 = _GEN_449;
  wire         compressDataVec_hitReq_6_91;
  assign compressDataVec_hitReq_6_91 = _GEN_449;
  wire         _GEN_450 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1B;
  wire         compressDataVec_hitReq_7_27;
  assign compressDataVec_hitReq_7_27 = _GEN_450;
  wire         compressDataVec_hitReq_7_91;
  assign compressDataVec_hitReq_7_91 = _GEN_450;
  wire         _GEN_451 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1B;
  wire         compressDataVec_hitReq_8_27;
  assign compressDataVec_hitReq_8_27 = _GEN_451;
  wire         compressDataVec_hitReq_8_91;
  assign compressDataVec_hitReq_8_91 = _GEN_451;
  wire         _GEN_452 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1B;
  wire         compressDataVec_hitReq_9_27;
  assign compressDataVec_hitReq_9_27 = _GEN_452;
  wire         compressDataVec_hitReq_9_91;
  assign compressDataVec_hitReq_9_91 = _GEN_452;
  wire         _GEN_453 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1B;
  wire         compressDataVec_hitReq_10_27;
  assign compressDataVec_hitReq_10_27 = _GEN_453;
  wire         compressDataVec_hitReq_10_91;
  assign compressDataVec_hitReq_10_91 = _GEN_453;
  wire         _GEN_454 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1B;
  wire         compressDataVec_hitReq_11_27;
  assign compressDataVec_hitReq_11_27 = _GEN_454;
  wire         compressDataVec_hitReq_11_91;
  assign compressDataVec_hitReq_11_91 = _GEN_454;
  wire         _GEN_455 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1B;
  wire         compressDataVec_hitReq_12_27;
  assign compressDataVec_hitReq_12_27 = _GEN_455;
  wire         compressDataVec_hitReq_12_91;
  assign compressDataVec_hitReq_12_91 = _GEN_455;
  wire         _GEN_456 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1B;
  wire         compressDataVec_hitReq_13_27;
  assign compressDataVec_hitReq_13_27 = _GEN_456;
  wire         compressDataVec_hitReq_13_91;
  assign compressDataVec_hitReq_13_91 = _GEN_456;
  wire         _GEN_457 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1B;
  wire         compressDataVec_hitReq_14_27;
  assign compressDataVec_hitReq_14_27 = _GEN_457;
  wire         compressDataVec_hitReq_14_91;
  assign compressDataVec_hitReq_14_91 = _GEN_457;
  wire         _GEN_458 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1B;
  wire         compressDataVec_hitReq_15_27;
  assign compressDataVec_hitReq_15_27 = _GEN_458;
  wire         compressDataVec_hitReq_15_91;
  assign compressDataVec_hitReq_15_91 = _GEN_458;
  wire         compressDataVec_hitReq_16_27 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1B;
  wire         compressDataVec_hitReq_17_27 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1B;
  wire         compressDataVec_hitReq_18_27 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1B;
  wire         compressDataVec_hitReq_19_27 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1B;
  wire         compressDataVec_hitReq_20_27 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1B;
  wire         compressDataVec_hitReq_21_27 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1B;
  wire         compressDataVec_hitReq_22_27 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1B;
  wire         compressDataVec_hitReq_23_27 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1B;
  wire         compressDataVec_hitReq_24_27 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1B;
  wire         compressDataVec_hitReq_25_27 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1B;
  wire         compressDataVec_hitReq_26_27 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1B;
  wire         compressDataVec_hitReq_27_27 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1B;
  wire         compressDataVec_hitReq_28_27 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1B;
  wire         compressDataVec_hitReq_29_27 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1B;
  wire         compressDataVec_hitReq_30_27 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1B;
  wire         compressDataVec_hitReq_31_27 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1B;
  wire [7:0]   compressDataVec_selectReqData_27 =
    (compressDataVec_hitReq_0_27 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_27 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_27 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_27 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_27 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_27 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_27 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_27 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_27 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_27 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_27 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_27 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_27 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_27 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_27 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_27 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_27 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_27 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_27 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_27 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_27 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_27 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_27 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_27 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_27 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_27 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_27 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_27 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_27 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_27 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_27 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_27 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_27 = tailCount > 5'h1B;
  wire         _GEN_459 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1C;
  wire         compressDataVec_hitReq_0_28;
  assign compressDataVec_hitReq_0_28 = _GEN_459;
  wire         compressDataVec_hitReq_0_92;
  assign compressDataVec_hitReq_0_92 = _GEN_459;
  wire         _GEN_460 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1C;
  wire         compressDataVec_hitReq_1_28;
  assign compressDataVec_hitReq_1_28 = _GEN_460;
  wire         compressDataVec_hitReq_1_92;
  assign compressDataVec_hitReq_1_92 = _GEN_460;
  wire         _GEN_461 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1C;
  wire         compressDataVec_hitReq_2_28;
  assign compressDataVec_hitReq_2_28 = _GEN_461;
  wire         compressDataVec_hitReq_2_92;
  assign compressDataVec_hitReq_2_92 = _GEN_461;
  wire         _GEN_462 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1C;
  wire         compressDataVec_hitReq_3_28;
  assign compressDataVec_hitReq_3_28 = _GEN_462;
  wire         compressDataVec_hitReq_3_92;
  assign compressDataVec_hitReq_3_92 = _GEN_462;
  wire         _GEN_463 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1C;
  wire         compressDataVec_hitReq_4_28;
  assign compressDataVec_hitReq_4_28 = _GEN_463;
  wire         compressDataVec_hitReq_4_92;
  assign compressDataVec_hitReq_4_92 = _GEN_463;
  wire         _GEN_464 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1C;
  wire         compressDataVec_hitReq_5_28;
  assign compressDataVec_hitReq_5_28 = _GEN_464;
  wire         compressDataVec_hitReq_5_92;
  assign compressDataVec_hitReq_5_92 = _GEN_464;
  wire         _GEN_465 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1C;
  wire         compressDataVec_hitReq_6_28;
  assign compressDataVec_hitReq_6_28 = _GEN_465;
  wire         compressDataVec_hitReq_6_92;
  assign compressDataVec_hitReq_6_92 = _GEN_465;
  wire         _GEN_466 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1C;
  wire         compressDataVec_hitReq_7_28;
  assign compressDataVec_hitReq_7_28 = _GEN_466;
  wire         compressDataVec_hitReq_7_92;
  assign compressDataVec_hitReq_7_92 = _GEN_466;
  wire         _GEN_467 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1C;
  wire         compressDataVec_hitReq_8_28;
  assign compressDataVec_hitReq_8_28 = _GEN_467;
  wire         compressDataVec_hitReq_8_92;
  assign compressDataVec_hitReq_8_92 = _GEN_467;
  wire         _GEN_468 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1C;
  wire         compressDataVec_hitReq_9_28;
  assign compressDataVec_hitReq_9_28 = _GEN_468;
  wire         compressDataVec_hitReq_9_92;
  assign compressDataVec_hitReq_9_92 = _GEN_468;
  wire         _GEN_469 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1C;
  wire         compressDataVec_hitReq_10_28;
  assign compressDataVec_hitReq_10_28 = _GEN_469;
  wire         compressDataVec_hitReq_10_92;
  assign compressDataVec_hitReq_10_92 = _GEN_469;
  wire         _GEN_470 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1C;
  wire         compressDataVec_hitReq_11_28;
  assign compressDataVec_hitReq_11_28 = _GEN_470;
  wire         compressDataVec_hitReq_11_92;
  assign compressDataVec_hitReq_11_92 = _GEN_470;
  wire         _GEN_471 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1C;
  wire         compressDataVec_hitReq_12_28;
  assign compressDataVec_hitReq_12_28 = _GEN_471;
  wire         compressDataVec_hitReq_12_92;
  assign compressDataVec_hitReq_12_92 = _GEN_471;
  wire         _GEN_472 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1C;
  wire         compressDataVec_hitReq_13_28;
  assign compressDataVec_hitReq_13_28 = _GEN_472;
  wire         compressDataVec_hitReq_13_92;
  assign compressDataVec_hitReq_13_92 = _GEN_472;
  wire         _GEN_473 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1C;
  wire         compressDataVec_hitReq_14_28;
  assign compressDataVec_hitReq_14_28 = _GEN_473;
  wire         compressDataVec_hitReq_14_92;
  assign compressDataVec_hitReq_14_92 = _GEN_473;
  wire         _GEN_474 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1C;
  wire         compressDataVec_hitReq_15_28;
  assign compressDataVec_hitReq_15_28 = _GEN_474;
  wire         compressDataVec_hitReq_15_92;
  assign compressDataVec_hitReq_15_92 = _GEN_474;
  wire         compressDataVec_hitReq_16_28 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1C;
  wire         compressDataVec_hitReq_17_28 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1C;
  wire         compressDataVec_hitReq_18_28 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1C;
  wire         compressDataVec_hitReq_19_28 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1C;
  wire         compressDataVec_hitReq_20_28 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1C;
  wire         compressDataVec_hitReq_21_28 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1C;
  wire         compressDataVec_hitReq_22_28 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1C;
  wire         compressDataVec_hitReq_23_28 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1C;
  wire         compressDataVec_hitReq_24_28 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1C;
  wire         compressDataVec_hitReq_25_28 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1C;
  wire         compressDataVec_hitReq_26_28 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1C;
  wire         compressDataVec_hitReq_27_28 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1C;
  wire         compressDataVec_hitReq_28_28 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1C;
  wire         compressDataVec_hitReq_29_28 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1C;
  wire         compressDataVec_hitReq_30_28 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1C;
  wire         compressDataVec_hitReq_31_28 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1C;
  wire [7:0]   compressDataVec_selectReqData_28 =
    (compressDataVec_hitReq_0_28 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_28 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_28 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_28 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_28 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_28 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_28 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_28 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_28 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_28 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_28 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_28 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_28 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_28 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_28 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_28 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_28 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_28 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_28 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_28 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_28 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_28 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_28 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_28 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_28 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_28 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_28 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_28 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_28 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_28 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_28 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_28 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_28 = tailCount > 5'h1C;
  wire         _GEN_475 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1D;
  wire         compressDataVec_hitReq_0_29;
  assign compressDataVec_hitReq_0_29 = _GEN_475;
  wire         compressDataVec_hitReq_0_93;
  assign compressDataVec_hitReq_0_93 = _GEN_475;
  wire         _GEN_476 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1D;
  wire         compressDataVec_hitReq_1_29;
  assign compressDataVec_hitReq_1_29 = _GEN_476;
  wire         compressDataVec_hitReq_1_93;
  assign compressDataVec_hitReq_1_93 = _GEN_476;
  wire         _GEN_477 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1D;
  wire         compressDataVec_hitReq_2_29;
  assign compressDataVec_hitReq_2_29 = _GEN_477;
  wire         compressDataVec_hitReq_2_93;
  assign compressDataVec_hitReq_2_93 = _GEN_477;
  wire         _GEN_478 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1D;
  wire         compressDataVec_hitReq_3_29;
  assign compressDataVec_hitReq_3_29 = _GEN_478;
  wire         compressDataVec_hitReq_3_93;
  assign compressDataVec_hitReq_3_93 = _GEN_478;
  wire         _GEN_479 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1D;
  wire         compressDataVec_hitReq_4_29;
  assign compressDataVec_hitReq_4_29 = _GEN_479;
  wire         compressDataVec_hitReq_4_93;
  assign compressDataVec_hitReq_4_93 = _GEN_479;
  wire         _GEN_480 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1D;
  wire         compressDataVec_hitReq_5_29;
  assign compressDataVec_hitReq_5_29 = _GEN_480;
  wire         compressDataVec_hitReq_5_93;
  assign compressDataVec_hitReq_5_93 = _GEN_480;
  wire         _GEN_481 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1D;
  wire         compressDataVec_hitReq_6_29;
  assign compressDataVec_hitReq_6_29 = _GEN_481;
  wire         compressDataVec_hitReq_6_93;
  assign compressDataVec_hitReq_6_93 = _GEN_481;
  wire         _GEN_482 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1D;
  wire         compressDataVec_hitReq_7_29;
  assign compressDataVec_hitReq_7_29 = _GEN_482;
  wire         compressDataVec_hitReq_7_93;
  assign compressDataVec_hitReq_7_93 = _GEN_482;
  wire         _GEN_483 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1D;
  wire         compressDataVec_hitReq_8_29;
  assign compressDataVec_hitReq_8_29 = _GEN_483;
  wire         compressDataVec_hitReq_8_93;
  assign compressDataVec_hitReq_8_93 = _GEN_483;
  wire         _GEN_484 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1D;
  wire         compressDataVec_hitReq_9_29;
  assign compressDataVec_hitReq_9_29 = _GEN_484;
  wire         compressDataVec_hitReq_9_93;
  assign compressDataVec_hitReq_9_93 = _GEN_484;
  wire         _GEN_485 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1D;
  wire         compressDataVec_hitReq_10_29;
  assign compressDataVec_hitReq_10_29 = _GEN_485;
  wire         compressDataVec_hitReq_10_93;
  assign compressDataVec_hitReq_10_93 = _GEN_485;
  wire         _GEN_486 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1D;
  wire         compressDataVec_hitReq_11_29;
  assign compressDataVec_hitReq_11_29 = _GEN_486;
  wire         compressDataVec_hitReq_11_93;
  assign compressDataVec_hitReq_11_93 = _GEN_486;
  wire         _GEN_487 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1D;
  wire         compressDataVec_hitReq_12_29;
  assign compressDataVec_hitReq_12_29 = _GEN_487;
  wire         compressDataVec_hitReq_12_93;
  assign compressDataVec_hitReq_12_93 = _GEN_487;
  wire         _GEN_488 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1D;
  wire         compressDataVec_hitReq_13_29;
  assign compressDataVec_hitReq_13_29 = _GEN_488;
  wire         compressDataVec_hitReq_13_93;
  assign compressDataVec_hitReq_13_93 = _GEN_488;
  wire         _GEN_489 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1D;
  wire         compressDataVec_hitReq_14_29;
  assign compressDataVec_hitReq_14_29 = _GEN_489;
  wire         compressDataVec_hitReq_14_93;
  assign compressDataVec_hitReq_14_93 = _GEN_489;
  wire         _GEN_490 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1D;
  wire         compressDataVec_hitReq_15_29;
  assign compressDataVec_hitReq_15_29 = _GEN_490;
  wire         compressDataVec_hitReq_15_93;
  assign compressDataVec_hitReq_15_93 = _GEN_490;
  wire         compressDataVec_hitReq_16_29 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1D;
  wire         compressDataVec_hitReq_17_29 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1D;
  wire         compressDataVec_hitReq_18_29 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1D;
  wire         compressDataVec_hitReq_19_29 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1D;
  wire         compressDataVec_hitReq_20_29 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1D;
  wire         compressDataVec_hitReq_21_29 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1D;
  wire         compressDataVec_hitReq_22_29 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1D;
  wire         compressDataVec_hitReq_23_29 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1D;
  wire         compressDataVec_hitReq_24_29 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1D;
  wire         compressDataVec_hitReq_25_29 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1D;
  wire         compressDataVec_hitReq_26_29 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1D;
  wire         compressDataVec_hitReq_27_29 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1D;
  wire         compressDataVec_hitReq_28_29 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1D;
  wire         compressDataVec_hitReq_29_29 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1D;
  wire         compressDataVec_hitReq_30_29 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1D;
  wire         compressDataVec_hitReq_31_29 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1D;
  wire [7:0]   compressDataVec_selectReqData_29 =
    (compressDataVec_hitReq_0_29 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_29 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_29 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_29 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_29 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_29 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_29 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_29 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_29 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_29 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_29 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_29 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_29 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_29 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_29 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_29 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_29 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_29 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_29 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_29 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_29 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_29 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_29 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_29 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_29 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_29 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_29 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_29 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_29 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_29 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_29 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_29 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_29 = tailCount > 5'h1D;
  wire         _GEN_491 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1E;
  wire         compressDataVec_hitReq_0_30;
  assign compressDataVec_hitReq_0_30 = _GEN_491;
  wire         compressDataVec_hitReq_0_94;
  assign compressDataVec_hitReq_0_94 = _GEN_491;
  wire         _GEN_492 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1E;
  wire         compressDataVec_hitReq_1_30;
  assign compressDataVec_hitReq_1_30 = _GEN_492;
  wire         compressDataVec_hitReq_1_94;
  assign compressDataVec_hitReq_1_94 = _GEN_492;
  wire         _GEN_493 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1E;
  wire         compressDataVec_hitReq_2_30;
  assign compressDataVec_hitReq_2_30 = _GEN_493;
  wire         compressDataVec_hitReq_2_94;
  assign compressDataVec_hitReq_2_94 = _GEN_493;
  wire         _GEN_494 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1E;
  wire         compressDataVec_hitReq_3_30;
  assign compressDataVec_hitReq_3_30 = _GEN_494;
  wire         compressDataVec_hitReq_3_94;
  assign compressDataVec_hitReq_3_94 = _GEN_494;
  wire         _GEN_495 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1E;
  wire         compressDataVec_hitReq_4_30;
  assign compressDataVec_hitReq_4_30 = _GEN_495;
  wire         compressDataVec_hitReq_4_94;
  assign compressDataVec_hitReq_4_94 = _GEN_495;
  wire         _GEN_496 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1E;
  wire         compressDataVec_hitReq_5_30;
  assign compressDataVec_hitReq_5_30 = _GEN_496;
  wire         compressDataVec_hitReq_5_94;
  assign compressDataVec_hitReq_5_94 = _GEN_496;
  wire         _GEN_497 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1E;
  wire         compressDataVec_hitReq_6_30;
  assign compressDataVec_hitReq_6_30 = _GEN_497;
  wire         compressDataVec_hitReq_6_94;
  assign compressDataVec_hitReq_6_94 = _GEN_497;
  wire         _GEN_498 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1E;
  wire         compressDataVec_hitReq_7_30;
  assign compressDataVec_hitReq_7_30 = _GEN_498;
  wire         compressDataVec_hitReq_7_94;
  assign compressDataVec_hitReq_7_94 = _GEN_498;
  wire         _GEN_499 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1E;
  wire         compressDataVec_hitReq_8_30;
  assign compressDataVec_hitReq_8_30 = _GEN_499;
  wire         compressDataVec_hitReq_8_94;
  assign compressDataVec_hitReq_8_94 = _GEN_499;
  wire         _GEN_500 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1E;
  wire         compressDataVec_hitReq_9_30;
  assign compressDataVec_hitReq_9_30 = _GEN_500;
  wire         compressDataVec_hitReq_9_94;
  assign compressDataVec_hitReq_9_94 = _GEN_500;
  wire         _GEN_501 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1E;
  wire         compressDataVec_hitReq_10_30;
  assign compressDataVec_hitReq_10_30 = _GEN_501;
  wire         compressDataVec_hitReq_10_94;
  assign compressDataVec_hitReq_10_94 = _GEN_501;
  wire         _GEN_502 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1E;
  wire         compressDataVec_hitReq_11_30;
  assign compressDataVec_hitReq_11_30 = _GEN_502;
  wire         compressDataVec_hitReq_11_94;
  assign compressDataVec_hitReq_11_94 = _GEN_502;
  wire         _GEN_503 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1E;
  wire         compressDataVec_hitReq_12_30;
  assign compressDataVec_hitReq_12_30 = _GEN_503;
  wire         compressDataVec_hitReq_12_94;
  assign compressDataVec_hitReq_12_94 = _GEN_503;
  wire         _GEN_504 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1E;
  wire         compressDataVec_hitReq_13_30;
  assign compressDataVec_hitReq_13_30 = _GEN_504;
  wire         compressDataVec_hitReq_13_94;
  assign compressDataVec_hitReq_13_94 = _GEN_504;
  wire         _GEN_505 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1E;
  wire         compressDataVec_hitReq_14_30;
  assign compressDataVec_hitReq_14_30 = _GEN_505;
  wire         compressDataVec_hitReq_14_94;
  assign compressDataVec_hitReq_14_94 = _GEN_505;
  wire         _GEN_506 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1E;
  wire         compressDataVec_hitReq_15_30;
  assign compressDataVec_hitReq_15_30 = _GEN_506;
  wire         compressDataVec_hitReq_15_94;
  assign compressDataVec_hitReq_15_94 = _GEN_506;
  wire         compressDataVec_hitReq_16_30 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1E;
  wire         compressDataVec_hitReq_17_30 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1E;
  wire         compressDataVec_hitReq_18_30 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1E;
  wire         compressDataVec_hitReq_19_30 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1E;
  wire         compressDataVec_hitReq_20_30 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1E;
  wire         compressDataVec_hitReq_21_30 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1E;
  wire         compressDataVec_hitReq_22_30 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1E;
  wire         compressDataVec_hitReq_23_30 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1E;
  wire         compressDataVec_hitReq_24_30 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1E;
  wire         compressDataVec_hitReq_25_30 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1E;
  wire         compressDataVec_hitReq_26_30 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1E;
  wire         compressDataVec_hitReq_27_30 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1E;
  wire         compressDataVec_hitReq_28_30 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1E;
  wire         compressDataVec_hitReq_29_30 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1E;
  wire         compressDataVec_hitReq_30_30 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1E;
  wire         compressDataVec_hitReq_31_30 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1E;
  wire [7:0]   compressDataVec_selectReqData_30 =
    (compressDataVec_hitReq_0_30 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_30 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_30 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_30 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_30 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_30 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_30 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_30 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_30 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_30 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_30 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_30 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_30 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_30 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_30 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_30 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_30 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_30 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_30 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_30 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_30 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_30 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_30 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_30 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_30 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_30 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_30 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_30 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_30 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_30 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_30 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_30 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_useTail_30 = &tailCount;
  wire         _GEN_507 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h1F;
  wire         compressDataVec_hitReq_0_31;
  assign compressDataVec_hitReq_0_31 = _GEN_507;
  wire         compressDataVec_hitReq_0_95;
  assign compressDataVec_hitReq_0_95 = _GEN_507;
  wire         _GEN_508 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h1F;
  wire         compressDataVec_hitReq_1_31;
  assign compressDataVec_hitReq_1_31 = _GEN_508;
  wire         compressDataVec_hitReq_1_95;
  assign compressDataVec_hitReq_1_95 = _GEN_508;
  wire         _GEN_509 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h1F;
  wire         compressDataVec_hitReq_2_31;
  assign compressDataVec_hitReq_2_31 = _GEN_509;
  wire         compressDataVec_hitReq_2_95;
  assign compressDataVec_hitReq_2_95 = _GEN_509;
  wire         _GEN_510 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h1F;
  wire         compressDataVec_hitReq_3_31;
  assign compressDataVec_hitReq_3_31 = _GEN_510;
  wire         compressDataVec_hitReq_3_95;
  assign compressDataVec_hitReq_3_95 = _GEN_510;
  wire         _GEN_511 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h1F;
  wire         compressDataVec_hitReq_4_31;
  assign compressDataVec_hitReq_4_31 = _GEN_511;
  wire         compressDataVec_hitReq_4_95;
  assign compressDataVec_hitReq_4_95 = _GEN_511;
  wire         _GEN_512 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h1F;
  wire         compressDataVec_hitReq_5_31;
  assign compressDataVec_hitReq_5_31 = _GEN_512;
  wire         compressDataVec_hitReq_5_95;
  assign compressDataVec_hitReq_5_95 = _GEN_512;
  wire         _GEN_513 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h1F;
  wire         compressDataVec_hitReq_6_31;
  assign compressDataVec_hitReq_6_31 = _GEN_513;
  wire         compressDataVec_hitReq_6_95;
  assign compressDataVec_hitReq_6_95 = _GEN_513;
  wire         _GEN_514 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h1F;
  wire         compressDataVec_hitReq_7_31;
  assign compressDataVec_hitReq_7_31 = _GEN_514;
  wire         compressDataVec_hitReq_7_95;
  assign compressDataVec_hitReq_7_95 = _GEN_514;
  wire         _GEN_515 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h1F;
  wire         compressDataVec_hitReq_8_31;
  assign compressDataVec_hitReq_8_31 = _GEN_515;
  wire         compressDataVec_hitReq_8_95;
  assign compressDataVec_hitReq_8_95 = _GEN_515;
  wire         _GEN_516 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h1F;
  wire         compressDataVec_hitReq_9_31;
  assign compressDataVec_hitReq_9_31 = _GEN_516;
  wire         compressDataVec_hitReq_9_95;
  assign compressDataVec_hitReq_9_95 = _GEN_516;
  wire         _GEN_517 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h1F;
  wire         compressDataVec_hitReq_10_31;
  assign compressDataVec_hitReq_10_31 = _GEN_517;
  wire         compressDataVec_hitReq_10_95;
  assign compressDataVec_hitReq_10_95 = _GEN_517;
  wire         _GEN_518 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h1F;
  wire         compressDataVec_hitReq_11_31;
  assign compressDataVec_hitReq_11_31 = _GEN_518;
  wire         compressDataVec_hitReq_11_95;
  assign compressDataVec_hitReq_11_95 = _GEN_518;
  wire         _GEN_519 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h1F;
  wire         compressDataVec_hitReq_12_31;
  assign compressDataVec_hitReq_12_31 = _GEN_519;
  wire         compressDataVec_hitReq_12_95;
  assign compressDataVec_hitReq_12_95 = _GEN_519;
  wire         _GEN_520 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h1F;
  wire         compressDataVec_hitReq_13_31;
  assign compressDataVec_hitReq_13_31 = _GEN_520;
  wire         compressDataVec_hitReq_13_95;
  assign compressDataVec_hitReq_13_95 = _GEN_520;
  wire         _GEN_521 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h1F;
  wire         compressDataVec_hitReq_14_31;
  assign compressDataVec_hitReq_14_31 = _GEN_521;
  wire         compressDataVec_hitReq_14_95;
  assign compressDataVec_hitReq_14_95 = _GEN_521;
  wire         _GEN_522 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h1F;
  wire         compressDataVec_hitReq_15_31;
  assign compressDataVec_hitReq_15_31 = _GEN_522;
  wire         compressDataVec_hitReq_15_95;
  assign compressDataVec_hitReq_15_95 = _GEN_522;
  wire         compressDataVec_hitReq_16_31 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h1F;
  wire         compressDataVec_hitReq_17_31 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h1F;
  wire         compressDataVec_hitReq_18_31 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h1F;
  wire         compressDataVec_hitReq_19_31 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h1F;
  wire         compressDataVec_hitReq_20_31 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h1F;
  wire         compressDataVec_hitReq_21_31 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h1F;
  wire         compressDataVec_hitReq_22_31 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h1F;
  wire         compressDataVec_hitReq_23_31 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h1F;
  wire         compressDataVec_hitReq_24_31 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h1F;
  wire         compressDataVec_hitReq_25_31 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h1F;
  wire         compressDataVec_hitReq_26_31 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h1F;
  wire         compressDataVec_hitReq_27_31 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h1F;
  wire         compressDataVec_hitReq_28_31 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h1F;
  wire         compressDataVec_hitReq_29_31 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h1F;
  wire         compressDataVec_hitReq_30_31 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h1F;
  wire         compressDataVec_hitReq_31_31 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h1F;
  wire [7:0]   compressDataVec_selectReqData_31 =
    (compressDataVec_hitReq_0_31 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_31 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_31 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_31 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_31 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_31 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_31 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_31 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_31 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_31 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_31 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_31 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_31 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_31 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_31 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_31 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_31 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_31 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_31 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_31 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_31 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_31 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_31 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_31 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_31 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_31 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_31 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_31 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_31 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_31 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_31 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_31 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_32 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h20;
  wire         compressDataVec_hitReq_1_32 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h20;
  wire         compressDataVec_hitReq_2_32 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h20;
  wire         compressDataVec_hitReq_3_32 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h20;
  wire         compressDataVec_hitReq_4_32 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h20;
  wire         compressDataVec_hitReq_5_32 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h20;
  wire         compressDataVec_hitReq_6_32 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h20;
  wire         compressDataVec_hitReq_7_32 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h20;
  wire         compressDataVec_hitReq_8_32 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h20;
  wire         compressDataVec_hitReq_9_32 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h20;
  wire         compressDataVec_hitReq_10_32 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h20;
  wire         compressDataVec_hitReq_11_32 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h20;
  wire         compressDataVec_hitReq_12_32 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h20;
  wire         compressDataVec_hitReq_13_32 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h20;
  wire         compressDataVec_hitReq_14_32 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h20;
  wire         compressDataVec_hitReq_15_32 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h20;
  wire         compressDataVec_hitReq_16_32 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h20;
  wire         compressDataVec_hitReq_17_32 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h20;
  wire         compressDataVec_hitReq_18_32 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h20;
  wire         compressDataVec_hitReq_19_32 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h20;
  wire         compressDataVec_hitReq_20_32 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h20;
  wire         compressDataVec_hitReq_21_32 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h20;
  wire         compressDataVec_hitReq_22_32 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h20;
  wire         compressDataVec_hitReq_23_32 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h20;
  wire         compressDataVec_hitReq_24_32 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h20;
  wire         compressDataVec_hitReq_25_32 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h20;
  wire         compressDataVec_hitReq_26_32 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h20;
  wire         compressDataVec_hitReq_27_32 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h20;
  wire         compressDataVec_hitReq_28_32 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h20;
  wire         compressDataVec_hitReq_29_32 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h20;
  wire         compressDataVec_hitReq_30_32 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h20;
  wire         compressDataVec_hitReq_31_32 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h20;
  wire [7:0]   compressDataVec_selectReqData_32 =
    (compressDataVec_hitReq_0_32 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_32 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_32 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_32 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_32 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_32 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_32 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_32 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_32 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_32 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_32 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_32 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_32 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_32 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_32 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_32 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_32 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_32 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_32 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_32 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_32 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_32 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_32 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_32 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_32 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_32 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_32 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_32 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_32 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_32 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_32 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_32 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_33 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h21;
  wire         compressDataVec_hitReq_1_33 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h21;
  wire         compressDataVec_hitReq_2_33 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h21;
  wire         compressDataVec_hitReq_3_33 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h21;
  wire         compressDataVec_hitReq_4_33 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h21;
  wire         compressDataVec_hitReq_5_33 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h21;
  wire         compressDataVec_hitReq_6_33 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h21;
  wire         compressDataVec_hitReq_7_33 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h21;
  wire         compressDataVec_hitReq_8_33 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h21;
  wire         compressDataVec_hitReq_9_33 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h21;
  wire         compressDataVec_hitReq_10_33 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h21;
  wire         compressDataVec_hitReq_11_33 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h21;
  wire         compressDataVec_hitReq_12_33 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h21;
  wire         compressDataVec_hitReq_13_33 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h21;
  wire         compressDataVec_hitReq_14_33 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h21;
  wire         compressDataVec_hitReq_15_33 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h21;
  wire         compressDataVec_hitReq_16_33 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h21;
  wire         compressDataVec_hitReq_17_33 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h21;
  wire         compressDataVec_hitReq_18_33 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h21;
  wire         compressDataVec_hitReq_19_33 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h21;
  wire         compressDataVec_hitReq_20_33 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h21;
  wire         compressDataVec_hitReq_21_33 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h21;
  wire         compressDataVec_hitReq_22_33 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h21;
  wire         compressDataVec_hitReq_23_33 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h21;
  wire         compressDataVec_hitReq_24_33 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h21;
  wire         compressDataVec_hitReq_25_33 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h21;
  wire         compressDataVec_hitReq_26_33 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h21;
  wire         compressDataVec_hitReq_27_33 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h21;
  wire         compressDataVec_hitReq_28_33 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h21;
  wire         compressDataVec_hitReq_29_33 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h21;
  wire         compressDataVec_hitReq_30_33 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h21;
  wire         compressDataVec_hitReq_31_33 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h21;
  wire [7:0]   compressDataVec_selectReqData_33 =
    (compressDataVec_hitReq_0_33 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_33 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_33 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_33 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_33 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_33 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_33 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_33 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_33 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_33 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_33 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_33 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_33 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_33 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_33 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_33 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_33 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_33 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_33 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_33 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_33 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_33 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_33 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_33 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_33 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_33 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_33 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_33 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_33 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_33 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_33 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_33 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_34 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h22;
  wire         compressDataVec_hitReq_1_34 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h22;
  wire         compressDataVec_hitReq_2_34 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h22;
  wire         compressDataVec_hitReq_3_34 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h22;
  wire         compressDataVec_hitReq_4_34 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h22;
  wire         compressDataVec_hitReq_5_34 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h22;
  wire         compressDataVec_hitReq_6_34 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h22;
  wire         compressDataVec_hitReq_7_34 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h22;
  wire         compressDataVec_hitReq_8_34 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h22;
  wire         compressDataVec_hitReq_9_34 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h22;
  wire         compressDataVec_hitReq_10_34 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h22;
  wire         compressDataVec_hitReq_11_34 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h22;
  wire         compressDataVec_hitReq_12_34 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h22;
  wire         compressDataVec_hitReq_13_34 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h22;
  wire         compressDataVec_hitReq_14_34 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h22;
  wire         compressDataVec_hitReq_15_34 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h22;
  wire         compressDataVec_hitReq_16_34 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h22;
  wire         compressDataVec_hitReq_17_34 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h22;
  wire         compressDataVec_hitReq_18_34 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h22;
  wire         compressDataVec_hitReq_19_34 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h22;
  wire         compressDataVec_hitReq_20_34 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h22;
  wire         compressDataVec_hitReq_21_34 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h22;
  wire         compressDataVec_hitReq_22_34 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h22;
  wire         compressDataVec_hitReq_23_34 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h22;
  wire         compressDataVec_hitReq_24_34 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h22;
  wire         compressDataVec_hitReq_25_34 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h22;
  wire         compressDataVec_hitReq_26_34 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h22;
  wire         compressDataVec_hitReq_27_34 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h22;
  wire         compressDataVec_hitReq_28_34 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h22;
  wire         compressDataVec_hitReq_29_34 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h22;
  wire         compressDataVec_hitReq_30_34 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h22;
  wire         compressDataVec_hitReq_31_34 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h22;
  wire [7:0]   compressDataVec_selectReqData_34 =
    (compressDataVec_hitReq_0_34 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_34 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_34 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_34 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_34 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_34 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_34 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_34 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_34 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_34 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_34 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_34 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_34 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_34 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_34 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_34 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_34 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_34 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_34 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_34 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_34 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_34 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_34 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_34 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_34 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_34 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_34 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_34 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_34 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_34 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_34 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_34 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_35 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h23;
  wire         compressDataVec_hitReq_1_35 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h23;
  wire         compressDataVec_hitReq_2_35 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h23;
  wire         compressDataVec_hitReq_3_35 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h23;
  wire         compressDataVec_hitReq_4_35 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h23;
  wire         compressDataVec_hitReq_5_35 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h23;
  wire         compressDataVec_hitReq_6_35 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h23;
  wire         compressDataVec_hitReq_7_35 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h23;
  wire         compressDataVec_hitReq_8_35 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h23;
  wire         compressDataVec_hitReq_9_35 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h23;
  wire         compressDataVec_hitReq_10_35 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h23;
  wire         compressDataVec_hitReq_11_35 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h23;
  wire         compressDataVec_hitReq_12_35 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h23;
  wire         compressDataVec_hitReq_13_35 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h23;
  wire         compressDataVec_hitReq_14_35 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h23;
  wire         compressDataVec_hitReq_15_35 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h23;
  wire         compressDataVec_hitReq_16_35 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h23;
  wire         compressDataVec_hitReq_17_35 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h23;
  wire         compressDataVec_hitReq_18_35 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h23;
  wire         compressDataVec_hitReq_19_35 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h23;
  wire         compressDataVec_hitReq_20_35 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h23;
  wire         compressDataVec_hitReq_21_35 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h23;
  wire         compressDataVec_hitReq_22_35 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h23;
  wire         compressDataVec_hitReq_23_35 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h23;
  wire         compressDataVec_hitReq_24_35 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h23;
  wire         compressDataVec_hitReq_25_35 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h23;
  wire         compressDataVec_hitReq_26_35 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h23;
  wire         compressDataVec_hitReq_27_35 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h23;
  wire         compressDataVec_hitReq_28_35 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h23;
  wire         compressDataVec_hitReq_29_35 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h23;
  wire         compressDataVec_hitReq_30_35 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h23;
  wire         compressDataVec_hitReq_31_35 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h23;
  wire [7:0]   compressDataVec_selectReqData_35 =
    (compressDataVec_hitReq_0_35 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_35 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_35 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_35 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_35 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_35 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_35 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_35 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_35 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_35 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_35 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_35 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_35 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_35 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_35 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_35 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_35 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_35 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_35 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_35 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_35 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_35 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_35 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_35 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_35 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_35 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_35 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_35 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_35 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_35 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_35 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_35 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_36 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h24;
  wire         compressDataVec_hitReq_1_36 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h24;
  wire         compressDataVec_hitReq_2_36 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h24;
  wire         compressDataVec_hitReq_3_36 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h24;
  wire         compressDataVec_hitReq_4_36 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h24;
  wire         compressDataVec_hitReq_5_36 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h24;
  wire         compressDataVec_hitReq_6_36 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h24;
  wire         compressDataVec_hitReq_7_36 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h24;
  wire         compressDataVec_hitReq_8_36 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h24;
  wire         compressDataVec_hitReq_9_36 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h24;
  wire         compressDataVec_hitReq_10_36 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h24;
  wire         compressDataVec_hitReq_11_36 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h24;
  wire         compressDataVec_hitReq_12_36 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h24;
  wire         compressDataVec_hitReq_13_36 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h24;
  wire         compressDataVec_hitReq_14_36 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h24;
  wire         compressDataVec_hitReq_15_36 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h24;
  wire         compressDataVec_hitReq_16_36 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h24;
  wire         compressDataVec_hitReq_17_36 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h24;
  wire         compressDataVec_hitReq_18_36 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h24;
  wire         compressDataVec_hitReq_19_36 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h24;
  wire         compressDataVec_hitReq_20_36 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h24;
  wire         compressDataVec_hitReq_21_36 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h24;
  wire         compressDataVec_hitReq_22_36 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h24;
  wire         compressDataVec_hitReq_23_36 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h24;
  wire         compressDataVec_hitReq_24_36 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h24;
  wire         compressDataVec_hitReq_25_36 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h24;
  wire         compressDataVec_hitReq_26_36 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h24;
  wire         compressDataVec_hitReq_27_36 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h24;
  wire         compressDataVec_hitReq_28_36 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h24;
  wire         compressDataVec_hitReq_29_36 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h24;
  wire         compressDataVec_hitReq_30_36 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h24;
  wire         compressDataVec_hitReq_31_36 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h24;
  wire [7:0]   compressDataVec_selectReqData_36 =
    (compressDataVec_hitReq_0_36 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_36 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_36 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_36 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_36 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_36 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_36 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_36 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_36 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_36 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_36 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_36 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_36 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_36 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_36 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_36 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_36 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_36 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_36 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_36 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_36 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_36 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_36 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_36 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_36 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_36 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_36 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_36 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_36 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_36 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_36 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_36 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_37 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h25;
  wire         compressDataVec_hitReq_1_37 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h25;
  wire         compressDataVec_hitReq_2_37 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h25;
  wire         compressDataVec_hitReq_3_37 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h25;
  wire         compressDataVec_hitReq_4_37 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h25;
  wire         compressDataVec_hitReq_5_37 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h25;
  wire         compressDataVec_hitReq_6_37 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h25;
  wire         compressDataVec_hitReq_7_37 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h25;
  wire         compressDataVec_hitReq_8_37 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h25;
  wire         compressDataVec_hitReq_9_37 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h25;
  wire         compressDataVec_hitReq_10_37 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h25;
  wire         compressDataVec_hitReq_11_37 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h25;
  wire         compressDataVec_hitReq_12_37 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h25;
  wire         compressDataVec_hitReq_13_37 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h25;
  wire         compressDataVec_hitReq_14_37 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h25;
  wire         compressDataVec_hitReq_15_37 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h25;
  wire         compressDataVec_hitReq_16_37 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h25;
  wire         compressDataVec_hitReq_17_37 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h25;
  wire         compressDataVec_hitReq_18_37 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h25;
  wire         compressDataVec_hitReq_19_37 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h25;
  wire         compressDataVec_hitReq_20_37 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h25;
  wire         compressDataVec_hitReq_21_37 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h25;
  wire         compressDataVec_hitReq_22_37 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h25;
  wire         compressDataVec_hitReq_23_37 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h25;
  wire         compressDataVec_hitReq_24_37 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h25;
  wire         compressDataVec_hitReq_25_37 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h25;
  wire         compressDataVec_hitReq_26_37 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h25;
  wire         compressDataVec_hitReq_27_37 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h25;
  wire         compressDataVec_hitReq_28_37 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h25;
  wire         compressDataVec_hitReq_29_37 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h25;
  wire         compressDataVec_hitReq_30_37 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h25;
  wire         compressDataVec_hitReq_31_37 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h25;
  wire [7:0]   compressDataVec_selectReqData_37 =
    (compressDataVec_hitReq_0_37 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_37 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_37 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_37 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_37 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_37 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_37 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_37 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_37 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_37 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_37 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_37 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_37 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_37 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_37 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_37 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_37 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_37 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_37 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_37 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_37 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_37 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_37 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_37 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_37 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_37 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_37 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_37 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_37 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_37 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_37 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_37 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_38 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h26;
  wire         compressDataVec_hitReq_1_38 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h26;
  wire         compressDataVec_hitReq_2_38 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h26;
  wire         compressDataVec_hitReq_3_38 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h26;
  wire         compressDataVec_hitReq_4_38 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h26;
  wire         compressDataVec_hitReq_5_38 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h26;
  wire         compressDataVec_hitReq_6_38 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h26;
  wire         compressDataVec_hitReq_7_38 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h26;
  wire         compressDataVec_hitReq_8_38 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h26;
  wire         compressDataVec_hitReq_9_38 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h26;
  wire         compressDataVec_hitReq_10_38 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h26;
  wire         compressDataVec_hitReq_11_38 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h26;
  wire         compressDataVec_hitReq_12_38 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h26;
  wire         compressDataVec_hitReq_13_38 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h26;
  wire         compressDataVec_hitReq_14_38 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h26;
  wire         compressDataVec_hitReq_15_38 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h26;
  wire         compressDataVec_hitReq_16_38 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h26;
  wire         compressDataVec_hitReq_17_38 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h26;
  wire         compressDataVec_hitReq_18_38 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h26;
  wire         compressDataVec_hitReq_19_38 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h26;
  wire         compressDataVec_hitReq_20_38 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h26;
  wire         compressDataVec_hitReq_21_38 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h26;
  wire         compressDataVec_hitReq_22_38 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h26;
  wire         compressDataVec_hitReq_23_38 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h26;
  wire         compressDataVec_hitReq_24_38 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h26;
  wire         compressDataVec_hitReq_25_38 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h26;
  wire         compressDataVec_hitReq_26_38 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h26;
  wire         compressDataVec_hitReq_27_38 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h26;
  wire         compressDataVec_hitReq_28_38 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h26;
  wire         compressDataVec_hitReq_29_38 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h26;
  wire         compressDataVec_hitReq_30_38 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h26;
  wire         compressDataVec_hitReq_31_38 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h26;
  wire [7:0]   compressDataVec_selectReqData_38 =
    (compressDataVec_hitReq_0_38 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_38 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_38 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_38 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_38 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_38 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_38 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_38 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_38 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_38 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_38 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_38 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_38 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_38 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_38 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_38 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_38 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_38 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_38 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_38 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_38 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_38 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_38 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_38 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_38 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_38 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_38 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_38 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_38 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_38 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_38 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_38 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_39 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h27;
  wire         compressDataVec_hitReq_1_39 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h27;
  wire         compressDataVec_hitReq_2_39 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h27;
  wire         compressDataVec_hitReq_3_39 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h27;
  wire         compressDataVec_hitReq_4_39 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h27;
  wire         compressDataVec_hitReq_5_39 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h27;
  wire         compressDataVec_hitReq_6_39 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h27;
  wire         compressDataVec_hitReq_7_39 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h27;
  wire         compressDataVec_hitReq_8_39 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h27;
  wire         compressDataVec_hitReq_9_39 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h27;
  wire         compressDataVec_hitReq_10_39 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h27;
  wire         compressDataVec_hitReq_11_39 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h27;
  wire         compressDataVec_hitReq_12_39 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h27;
  wire         compressDataVec_hitReq_13_39 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h27;
  wire         compressDataVec_hitReq_14_39 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h27;
  wire         compressDataVec_hitReq_15_39 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h27;
  wire         compressDataVec_hitReq_16_39 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h27;
  wire         compressDataVec_hitReq_17_39 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h27;
  wire         compressDataVec_hitReq_18_39 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h27;
  wire         compressDataVec_hitReq_19_39 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h27;
  wire         compressDataVec_hitReq_20_39 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h27;
  wire         compressDataVec_hitReq_21_39 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h27;
  wire         compressDataVec_hitReq_22_39 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h27;
  wire         compressDataVec_hitReq_23_39 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h27;
  wire         compressDataVec_hitReq_24_39 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h27;
  wire         compressDataVec_hitReq_25_39 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h27;
  wire         compressDataVec_hitReq_26_39 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h27;
  wire         compressDataVec_hitReq_27_39 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h27;
  wire         compressDataVec_hitReq_28_39 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h27;
  wire         compressDataVec_hitReq_29_39 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h27;
  wire         compressDataVec_hitReq_30_39 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h27;
  wire         compressDataVec_hitReq_31_39 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h27;
  wire [7:0]   compressDataVec_selectReqData_39 =
    (compressDataVec_hitReq_0_39 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_39 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_39 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_39 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_39 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_39 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_39 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_39 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_39 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_39 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_39 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_39 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_39 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_39 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_39 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_39 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_39 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_39 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_39 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_39 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_39 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_39 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_39 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_39 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_39 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_39 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_39 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_39 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_39 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_39 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_39 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_39 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_40 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h28;
  wire         compressDataVec_hitReq_1_40 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h28;
  wire         compressDataVec_hitReq_2_40 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h28;
  wire         compressDataVec_hitReq_3_40 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h28;
  wire         compressDataVec_hitReq_4_40 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h28;
  wire         compressDataVec_hitReq_5_40 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h28;
  wire         compressDataVec_hitReq_6_40 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h28;
  wire         compressDataVec_hitReq_7_40 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h28;
  wire         compressDataVec_hitReq_8_40 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h28;
  wire         compressDataVec_hitReq_9_40 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h28;
  wire         compressDataVec_hitReq_10_40 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h28;
  wire         compressDataVec_hitReq_11_40 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h28;
  wire         compressDataVec_hitReq_12_40 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h28;
  wire         compressDataVec_hitReq_13_40 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h28;
  wire         compressDataVec_hitReq_14_40 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h28;
  wire         compressDataVec_hitReq_15_40 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h28;
  wire         compressDataVec_hitReq_16_40 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h28;
  wire         compressDataVec_hitReq_17_40 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h28;
  wire         compressDataVec_hitReq_18_40 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h28;
  wire         compressDataVec_hitReq_19_40 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h28;
  wire         compressDataVec_hitReq_20_40 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h28;
  wire         compressDataVec_hitReq_21_40 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h28;
  wire         compressDataVec_hitReq_22_40 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h28;
  wire         compressDataVec_hitReq_23_40 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h28;
  wire         compressDataVec_hitReq_24_40 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h28;
  wire         compressDataVec_hitReq_25_40 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h28;
  wire         compressDataVec_hitReq_26_40 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h28;
  wire         compressDataVec_hitReq_27_40 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h28;
  wire         compressDataVec_hitReq_28_40 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h28;
  wire         compressDataVec_hitReq_29_40 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h28;
  wire         compressDataVec_hitReq_30_40 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h28;
  wire         compressDataVec_hitReq_31_40 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h28;
  wire [7:0]   compressDataVec_selectReqData_40 =
    (compressDataVec_hitReq_0_40 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_40 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_40 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_40 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_40 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_40 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_40 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_40 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_40 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_40 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_40 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_40 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_40 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_40 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_40 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_40 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_40 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_40 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_40 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_40 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_40 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_40 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_40 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_40 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_40 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_40 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_40 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_40 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_40 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_40 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_40 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_40 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_41 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h29;
  wire         compressDataVec_hitReq_1_41 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h29;
  wire         compressDataVec_hitReq_2_41 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h29;
  wire         compressDataVec_hitReq_3_41 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h29;
  wire         compressDataVec_hitReq_4_41 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h29;
  wire         compressDataVec_hitReq_5_41 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h29;
  wire         compressDataVec_hitReq_6_41 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h29;
  wire         compressDataVec_hitReq_7_41 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h29;
  wire         compressDataVec_hitReq_8_41 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h29;
  wire         compressDataVec_hitReq_9_41 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h29;
  wire         compressDataVec_hitReq_10_41 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h29;
  wire         compressDataVec_hitReq_11_41 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h29;
  wire         compressDataVec_hitReq_12_41 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h29;
  wire         compressDataVec_hitReq_13_41 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h29;
  wire         compressDataVec_hitReq_14_41 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h29;
  wire         compressDataVec_hitReq_15_41 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h29;
  wire         compressDataVec_hitReq_16_41 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h29;
  wire         compressDataVec_hitReq_17_41 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h29;
  wire         compressDataVec_hitReq_18_41 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h29;
  wire         compressDataVec_hitReq_19_41 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h29;
  wire         compressDataVec_hitReq_20_41 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h29;
  wire         compressDataVec_hitReq_21_41 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h29;
  wire         compressDataVec_hitReq_22_41 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h29;
  wire         compressDataVec_hitReq_23_41 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h29;
  wire         compressDataVec_hitReq_24_41 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h29;
  wire         compressDataVec_hitReq_25_41 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h29;
  wire         compressDataVec_hitReq_26_41 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h29;
  wire         compressDataVec_hitReq_27_41 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h29;
  wire         compressDataVec_hitReq_28_41 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h29;
  wire         compressDataVec_hitReq_29_41 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h29;
  wire         compressDataVec_hitReq_30_41 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h29;
  wire         compressDataVec_hitReq_31_41 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h29;
  wire [7:0]   compressDataVec_selectReqData_41 =
    (compressDataVec_hitReq_0_41 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_41 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_41 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_41 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_41 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_41 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_41 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_41 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_41 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_41 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_41 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_41 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_41 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_41 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_41 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_41 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_41 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_41 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_41 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_41 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_41 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_41 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_41 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_41 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_41 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_41 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_41 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_41 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_41 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_41 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_41 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_41 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_42 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2A;
  wire         compressDataVec_hitReq_1_42 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2A;
  wire         compressDataVec_hitReq_2_42 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2A;
  wire         compressDataVec_hitReq_3_42 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2A;
  wire         compressDataVec_hitReq_4_42 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2A;
  wire         compressDataVec_hitReq_5_42 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2A;
  wire         compressDataVec_hitReq_6_42 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2A;
  wire         compressDataVec_hitReq_7_42 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2A;
  wire         compressDataVec_hitReq_8_42 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2A;
  wire         compressDataVec_hitReq_9_42 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2A;
  wire         compressDataVec_hitReq_10_42 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2A;
  wire         compressDataVec_hitReq_11_42 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2A;
  wire         compressDataVec_hitReq_12_42 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2A;
  wire         compressDataVec_hitReq_13_42 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2A;
  wire         compressDataVec_hitReq_14_42 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2A;
  wire         compressDataVec_hitReq_15_42 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2A;
  wire         compressDataVec_hitReq_16_42 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2A;
  wire         compressDataVec_hitReq_17_42 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2A;
  wire         compressDataVec_hitReq_18_42 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2A;
  wire         compressDataVec_hitReq_19_42 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2A;
  wire         compressDataVec_hitReq_20_42 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2A;
  wire         compressDataVec_hitReq_21_42 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2A;
  wire         compressDataVec_hitReq_22_42 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2A;
  wire         compressDataVec_hitReq_23_42 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2A;
  wire         compressDataVec_hitReq_24_42 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2A;
  wire         compressDataVec_hitReq_25_42 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2A;
  wire         compressDataVec_hitReq_26_42 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2A;
  wire         compressDataVec_hitReq_27_42 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2A;
  wire         compressDataVec_hitReq_28_42 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2A;
  wire         compressDataVec_hitReq_29_42 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2A;
  wire         compressDataVec_hitReq_30_42 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2A;
  wire         compressDataVec_hitReq_31_42 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2A;
  wire [7:0]   compressDataVec_selectReqData_42 =
    (compressDataVec_hitReq_0_42 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_42 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_42 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_42 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_42 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_42 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_42 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_42 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_42 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_42 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_42 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_42 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_42 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_42 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_42 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_42 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_42 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_42 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_42 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_42 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_42 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_42 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_42 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_42 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_42 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_42 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_42 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_42 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_42 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_42 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_42 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_42 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_43 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2B;
  wire         compressDataVec_hitReq_1_43 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2B;
  wire         compressDataVec_hitReq_2_43 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2B;
  wire         compressDataVec_hitReq_3_43 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2B;
  wire         compressDataVec_hitReq_4_43 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2B;
  wire         compressDataVec_hitReq_5_43 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2B;
  wire         compressDataVec_hitReq_6_43 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2B;
  wire         compressDataVec_hitReq_7_43 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2B;
  wire         compressDataVec_hitReq_8_43 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2B;
  wire         compressDataVec_hitReq_9_43 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2B;
  wire         compressDataVec_hitReq_10_43 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2B;
  wire         compressDataVec_hitReq_11_43 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2B;
  wire         compressDataVec_hitReq_12_43 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2B;
  wire         compressDataVec_hitReq_13_43 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2B;
  wire         compressDataVec_hitReq_14_43 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2B;
  wire         compressDataVec_hitReq_15_43 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2B;
  wire         compressDataVec_hitReq_16_43 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2B;
  wire         compressDataVec_hitReq_17_43 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2B;
  wire         compressDataVec_hitReq_18_43 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2B;
  wire         compressDataVec_hitReq_19_43 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2B;
  wire         compressDataVec_hitReq_20_43 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2B;
  wire         compressDataVec_hitReq_21_43 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2B;
  wire         compressDataVec_hitReq_22_43 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2B;
  wire         compressDataVec_hitReq_23_43 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2B;
  wire         compressDataVec_hitReq_24_43 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2B;
  wire         compressDataVec_hitReq_25_43 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2B;
  wire         compressDataVec_hitReq_26_43 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2B;
  wire         compressDataVec_hitReq_27_43 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2B;
  wire         compressDataVec_hitReq_28_43 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2B;
  wire         compressDataVec_hitReq_29_43 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2B;
  wire         compressDataVec_hitReq_30_43 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2B;
  wire         compressDataVec_hitReq_31_43 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2B;
  wire [7:0]   compressDataVec_selectReqData_43 =
    (compressDataVec_hitReq_0_43 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_43 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_43 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_43 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_43 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_43 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_43 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_43 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_43 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_43 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_43 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_43 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_43 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_43 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_43 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_43 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_43 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_43 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_43 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_43 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_43 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_43 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_43 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_43 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_43 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_43 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_43 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_43 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_43 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_43 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_43 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_43 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_44 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2C;
  wire         compressDataVec_hitReq_1_44 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2C;
  wire         compressDataVec_hitReq_2_44 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2C;
  wire         compressDataVec_hitReq_3_44 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2C;
  wire         compressDataVec_hitReq_4_44 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2C;
  wire         compressDataVec_hitReq_5_44 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2C;
  wire         compressDataVec_hitReq_6_44 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2C;
  wire         compressDataVec_hitReq_7_44 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2C;
  wire         compressDataVec_hitReq_8_44 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2C;
  wire         compressDataVec_hitReq_9_44 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2C;
  wire         compressDataVec_hitReq_10_44 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2C;
  wire         compressDataVec_hitReq_11_44 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2C;
  wire         compressDataVec_hitReq_12_44 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2C;
  wire         compressDataVec_hitReq_13_44 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2C;
  wire         compressDataVec_hitReq_14_44 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2C;
  wire         compressDataVec_hitReq_15_44 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2C;
  wire         compressDataVec_hitReq_16_44 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2C;
  wire         compressDataVec_hitReq_17_44 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2C;
  wire         compressDataVec_hitReq_18_44 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2C;
  wire         compressDataVec_hitReq_19_44 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2C;
  wire         compressDataVec_hitReq_20_44 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2C;
  wire         compressDataVec_hitReq_21_44 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2C;
  wire         compressDataVec_hitReq_22_44 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2C;
  wire         compressDataVec_hitReq_23_44 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2C;
  wire         compressDataVec_hitReq_24_44 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2C;
  wire         compressDataVec_hitReq_25_44 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2C;
  wire         compressDataVec_hitReq_26_44 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2C;
  wire         compressDataVec_hitReq_27_44 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2C;
  wire         compressDataVec_hitReq_28_44 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2C;
  wire         compressDataVec_hitReq_29_44 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2C;
  wire         compressDataVec_hitReq_30_44 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2C;
  wire         compressDataVec_hitReq_31_44 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2C;
  wire [7:0]   compressDataVec_selectReqData_44 =
    (compressDataVec_hitReq_0_44 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_44 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_44 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_44 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_44 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_44 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_44 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_44 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_44 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_44 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_44 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_44 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_44 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_44 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_44 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_44 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_44 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_44 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_44 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_44 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_44 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_44 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_44 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_44 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_44 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_44 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_44 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_44 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_44 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_44 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_44 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_44 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_45 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2D;
  wire         compressDataVec_hitReq_1_45 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2D;
  wire         compressDataVec_hitReq_2_45 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2D;
  wire         compressDataVec_hitReq_3_45 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2D;
  wire         compressDataVec_hitReq_4_45 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2D;
  wire         compressDataVec_hitReq_5_45 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2D;
  wire         compressDataVec_hitReq_6_45 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2D;
  wire         compressDataVec_hitReq_7_45 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2D;
  wire         compressDataVec_hitReq_8_45 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2D;
  wire         compressDataVec_hitReq_9_45 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2D;
  wire         compressDataVec_hitReq_10_45 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2D;
  wire         compressDataVec_hitReq_11_45 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2D;
  wire         compressDataVec_hitReq_12_45 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2D;
  wire         compressDataVec_hitReq_13_45 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2D;
  wire         compressDataVec_hitReq_14_45 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2D;
  wire         compressDataVec_hitReq_15_45 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2D;
  wire         compressDataVec_hitReq_16_45 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2D;
  wire         compressDataVec_hitReq_17_45 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2D;
  wire         compressDataVec_hitReq_18_45 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2D;
  wire         compressDataVec_hitReq_19_45 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2D;
  wire         compressDataVec_hitReq_20_45 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2D;
  wire         compressDataVec_hitReq_21_45 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2D;
  wire         compressDataVec_hitReq_22_45 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2D;
  wire         compressDataVec_hitReq_23_45 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2D;
  wire         compressDataVec_hitReq_24_45 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2D;
  wire         compressDataVec_hitReq_25_45 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2D;
  wire         compressDataVec_hitReq_26_45 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2D;
  wire         compressDataVec_hitReq_27_45 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2D;
  wire         compressDataVec_hitReq_28_45 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2D;
  wire         compressDataVec_hitReq_29_45 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2D;
  wire         compressDataVec_hitReq_30_45 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2D;
  wire         compressDataVec_hitReq_31_45 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2D;
  wire [7:0]   compressDataVec_selectReqData_45 =
    (compressDataVec_hitReq_0_45 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_45 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_45 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_45 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_45 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_45 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_45 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_45 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_45 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_45 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_45 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_45 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_45 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_45 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_45 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_45 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_45 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_45 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_45 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_45 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_45 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_45 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_45 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_45 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_45 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_45 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_45 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_45 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_45 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_45 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_45 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_45 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_46 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2E;
  wire         compressDataVec_hitReq_1_46 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2E;
  wire         compressDataVec_hitReq_2_46 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2E;
  wire         compressDataVec_hitReq_3_46 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2E;
  wire         compressDataVec_hitReq_4_46 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2E;
  wire         compressDataVec_hitReq_5_46 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2E;
  wire         compressDataVec_hitReq_6_46 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2E;
  wire         compressDataVec_hitReq_7_46 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2E;
  wire         compressDataVec_hitReq_8_46 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2E;
  wire         compressDataVec_hitReq_9_46 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2E;
  wire         compressDataVec_hitReq_10_46 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2E;
  wire         compressDataVec_hitReq_11_46 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2E;
  wire         compressDataVec_hitReq_12_46 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2E;
  wire         compressDataVec_hitReq_13_46 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2E;
  wire         compressDataVec_hitReq_14_46 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2E;
  wire         compressDataVec_hitReq_15_46 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2E;
  wire         compressDataVec_hitReq_16_46 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2E;
  wire         compressDataVec_hitReq_17_46 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2E;
  wire         compressDataVec_hitReq_18_46 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2E;
  wire         compressDataVec_hitReq_19_46 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2E;
  wire         compressDataVec_hitReq_20_46 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2E;
  wire         compressDataVec_hitReq_21_46 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2E;
  wire         compressDataVec_hitReq_22_46 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2E;
  wire         compressDataVec_hitReq_23_46 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2E;
  wire         compressDataVec_hitReq_24_46 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2E;
  wire         compressDataVec_hitReq_25_46 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2E;
  wire         compressDataVec_hitReq_26_46 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2E;
  wire         compressDataVec_hitReq_27_46 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2E;
  wire         compressDataVec_hitReq_28_46 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2E;
  wire         compressDataVec_hitReq_29_46 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2E;
  wire         compressDataVec_hitReq_30_46 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2E;
  wire         compressDataVec_hitReq_31_46 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2E;
  wire [7:0]   compressDataVec_selectReqData_46 =
    (compressDataVec_hitReq_0_46 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_46 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_46 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_46 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_46 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_46 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_46 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_46 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_46 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_46 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_46 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_46 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_46 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_46 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_46 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_46 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_46 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_46 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_46 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_46 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_46 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_46 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_46 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_46 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_46 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_46 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_46 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_46 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_46 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_46 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_46 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_46 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_47 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h2F;
  wire         compressDataVec_hitReq_1_47 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h2F;
  wire         compressDataVec_hitReq_2_47 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h2F;
  wire         compressDataVec_hitReq_3_47 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h2F;
  wire         compressDataVec_hitReq_4_47 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h2F;
  wire         compressDataVec_hitReq_5_47 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h2F;
  wire         compressDataVec_hitReq_6_47 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h2F;
  wire         compressDataVec_hitReq_7_47 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h2F;
  wire         compressDataVec_hitReq_8_47 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h2F;
  wire         compressDataVec_hitReq_9_47 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h2F;
  wire         compressDataVec_hitReq_10_47 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h2F;
  wire         compressDataVec_hitReq_11_47 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h2F;
  wire         compressDataVec_hitReq_12_47 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h2F;
  wire         compressDataVec_hitReq_13_47 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h2F;
  wire         compressDataVec_hitReq_14_47 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h2F;
  wire         compressDataVec_hitReq_15_47 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h2F;
  wire         compressDataVec_hitReq_16_47 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h2F;
  wire         compressDataVec_hitReq_17_47 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h2F;
  wire         compressDataVec_hitReq_18_47 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h2F;
  wire         compressDataVec_hitReq_19_47 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h2F;
  wire         compressDataVec_hitReq_20_47 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h2F;
  wire         compressDataVec_hitReq_21_47 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h2F;
  wire         compressDataVec_hitReq_22_47 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h2F;
  wire         compressDataVec_hitReq_23_47 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h2F;
  wire         compressDataVec_hitReq_24_47 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h2F;
  wire         compressDataVec_hitReq_25_47 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h2F;
  wire         compressDataVec_hitReq_26_47 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h2F;
  wire         compressDataVec_hitReq_27_47 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h2F;
  wire         compressDataVec_hitReq_28_47 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h2F;
  wire         compressDataVec_hitReq_29_47 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h2F;
  wire         compressDataVec_hitReq_30_47 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h2F;
  wire         compressDataVec_hitReq_31_47 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h2F;
  wire [7:0]   compressDataVec_selectReqData_47 =
    (compressDataVec_hitReq_0_47 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_47 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_47 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_47 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_47 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_47 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_47 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_47 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_47 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_47 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_47 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_47 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_47 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_47 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_47 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_47 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_47 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_47 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_47 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_47 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_47 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_47 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_47 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_47 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_47 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_47 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_47 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_47 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_47 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_47 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_47 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_47 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_48 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h30;
  wire         compressDataVec_hitReq_1_48 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h30;
  wire         compressDataVec_hitReq_2_48 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h30;
  wire         compressDataVec_hitReq_3_48 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h30;
  wire         compressDataVec_hitReq_4_48 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h30;
  wire         compressDataVec_hitReq_5_48 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h30;
  wire         compressDataVec_hitReq_6_48 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h30;
  wire         compressDataVec_hitReq_7_48 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h30;
  wire         compressDataVec_hitReq_8_48 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h30;
  wire         compressDataVec_hitReq_9_48 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h30;
  wire         compressDataVec_hitReq_10_48 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h30;
  wire         compressDataVec_hitReq_11_48 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h30;
  wire         compressDataVec_hitReq_12_48 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h30;
  wire         compressDataVec_hitReq_13_48 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h30;
  wire         compressDataVec_hitReq_14_48 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h30;
  wire         compressDataVec_hitReq_15_48 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h30;
  wire         compressDataVec_hitReq_16_48 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h30;
  wire         compressDataVec_hitReq_17_48 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h30;
  wire         compressDataVec_hitReq_18_48 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h30;
  wire         compressDataVec_hitReq_19_48 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h30;
  wire         compressDataVec_hitReq_20_48 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h30;
  wire         compressDataVec_hitReq_21_48 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h30;
  wire         compressDataVec_hitReq_22_48 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h30;
  wire         compressDataVec_hitReq_23_48 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h30;
  wire         compressDataVec_hitReq_24_48 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h30;
  wire         compressDataVec_hitReq_25_48 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h30;
  wire         compressDataVec_hitReq_26_48 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h30;
  wire         compressDataVec_hitReq_27_48 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h30;
  wire         compressDataVec_hitReq_28_48 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h30;
  wire         compressDataVec_hitReq_29_48 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h30;
  wire         compressDataVec_hitReq_30_48 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h30;
  wire         compressDataVec_hitReq_31_48 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h30;
  wire [7:0]   compressDataVec_selectReqData_48 =
    (compressDataVec_hitReq_0_48 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_48 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_48 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_48 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_48 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_48 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_48 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_48 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_48 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_48 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_48 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_48 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_48 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_48 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_48 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_48 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_48 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_48 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_48 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_48 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_48 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_48 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_48 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_48 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_48 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_48 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_48 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_48 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_48 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_48 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_48 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_48 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_49 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h31;
  wire         compressDataVec_hitReq_1_49 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h31;
  wire         compressDataVec_hitReq_2_49 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h31;
  wire         compressDataVec_hitReq_3_49 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h31;
  wire         compressDataVec_hitReq_4_49 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h31;
  wire         compressDataVec_hitReq_5_49 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h31;
  wire         compressDataVec_hitReq_6_49 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h31;
  wire         compressDataVec_hitReq_7_49 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h31;
  wire         compressDataVec_hitReq_8_49 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h31;
  wire         compressDataVec_hitReq_9_49 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h31;
  wire         compressDataVec_hitReq_10_49 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h31;
  wire         compressDataVec_hitReq_11_49 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h31;
  wire         compressDataVec_hitReq_12_49 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h31;
  wire         compressDataVec_hitReq_13_49 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h31;
  wire         compressDataVec_hitReq_14_49 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h31;
  wire         compressDataVec_hitReq_15_49 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h31;
  wire         compressDataVec_hitReq_16_49 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h31;
  wire         compressDataVec_hitReq_17_49 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h31;
  wire         compressDataVec_hitReq_18_49 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h31;
  wire         compressDataVec_hitReq_19_49 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h31;
  wire         compressDataVec_hitReq_20_49 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h31;
  wire         compressDataVec_hitReq_21_49 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h31;
  wire         compressDataVec_hitReq_22_49 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h31;
  wire         compressDataVec_hitReq_23_49 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h31;
  wire         compressDataVec_hitReq_24_49 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h31;
  wire         compressDataVec_hitReq_25_49 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h31;
  wire         compressDataVec_hitReq_26_49 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h31;
  wire         compressDataVec_hitReq_27_49 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h31;
  wire         compressDataVec_hitReq_28_49 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h31;
  wire         compressDataVec_hitReq_29_49 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h31;
  wire         compressDataVec_hitReq_30_49 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h31;
  wire         compressDataVec_hitReq_31_49 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h31;
  wire [7:0]   compressDataVec_selectReqData_49 =
    (compressDataVec_hitReq_0_49 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_49 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_49 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_49 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_49 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_49 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_49 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_49 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_49 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_49 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_49 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_49 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_49 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_49 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_49 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_49 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_49 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_49 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_49 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_49 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_49 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_49 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_49 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_49 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_49 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_49 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_49 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_49 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_49 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_49 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_49 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_49 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_50 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h32;
  wire         compressDataVec_hitReq_1_50 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h32;
  wire         compressDataVec_hitReq_2_50 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h32;
  wire         compressDataVec_hitReq_3_50 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h32;
  wire         compressDataVec_hitReq_4_50 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h32;
  wire         compressDataVec_hitReq_5_50 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h32;
  wire         compressDataVec_hitReq_6_50 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h32;
  wire         compressDataVec_hitReq_7_50 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h32;
  wire         compressDataVec_hitReq_8_50 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h32;
  wire         compressDataVec_hitReq_9_50 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h32;
  wire         compressDataVec_hitReq_10_50 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h32;
  wire         compressDataVec_hitReq_11_50 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h32;
  wire         compressDataVec_hitReq_12_50 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h32;
  wire         compressDataVec_hitReq_13_50 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h32;
  wire         compressDataVec_hitReq_14_50 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h32;
  wire         compressDataVec_hitReq_15_50 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h32;
  wire         compressDataVec_hitReq_16_50 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h32;
  wire         compressDataVec_hitReq_17_50 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h32;
  wire         compressDataVec_hitReq_18_50 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h32;
  wire         compressDataVec_hitReq_19_50 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h32;
  wire         compressDataVec_hitReq_20_50 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h32;
  wire         compressDataVec_hitReq_21_50 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h32;
  wire         compressDataVec_hitReq_22_50 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h32;
  wire         compressDataVec_hitReq_23_50 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h32;
  wire         compressDataVec_hitReq_24_50 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h32;
  wire         compressDataVec_hitReq_25_50 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h32;
  wire         compressDataVec_hitReq_26_50 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h32;
  wire         compressDataVec_hitReq_27_50 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h32;
  wire         compressDataVec_hitReq_28_50 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h32;
  wire         compressDataVec_hitReq_29_50 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h32;
  wire         compressDataVec_hitReq_30_50 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h32;
  wire         compressDataVec_hitReq_31_50 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h32;
  wire [7:0]   compressDataVec_selectReqData_50 =
    (compressDataVec_hitReq_0_50 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_50 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_50 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_50 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_50 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_50 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_50 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_50 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_50 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_50 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_50 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_50 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_50 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_50 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_50 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_50 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_50 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_50 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_50 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_50 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_50 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_50 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_50 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_50 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_50 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_50 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_50 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_50 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_50 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_50 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_50 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_50 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_51 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h33;
  wire         compressDataVec_hitReq_1_51 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h33;
  wire         compressDataVec_hitReq_2_51 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h33;
  wire         compressDataVec_hitReq_3_51 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h33;
  wire         compressDataVec_hitReq_4_51 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h33;
  wire         compressDataVec_hitReq_5_51 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h33;
  wire         compressDataVec_hitReq_6_51 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h33;
  wire         compressDataVec_hitReq_7_51 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h33;
  wire         compressDataVec_hitReq_8_51 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h33;
  wire         compressDataVec_hitReq_9_51 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h33;
  wire         compressDataVec_hitReq_10_51 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h33;
  wire         compressDataVec_hitReq_11_51 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h33;
  wire         compressDataVec_hitReq_12_51 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h33;
  wire         compressDataVec_hitReq_13_51 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h33;
  wire         compressDataVec_hitReq_14_51 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h33;
  wire         compressDataVec_hitReq_15_51 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h33;
  wire         compressDataVec_hitReq_16_51 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h33;
  wire         compressDataVec_hitReq_17_51 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h33;
  wire         compressDataVec_hitReq_18_51 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h33;
  wire         compressDataVec_hitReq_19_51 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h33;
  wire         compressDataVec_hitReq_20_51 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h33;
  wire         compressDataVec_hitReq_21_51 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h33;
  wire         compressDataVec_hitReq_22_51 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h33;
  wire         compressDataVec_hitReq_23_51 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h33;
  wire         compressDataVec_hitReq_24_51 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h33;
  wire         compressDataVec_hitReq_25_51 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h33;
  wire         compressDataVec_hitReq_26_51 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h33;
  wire         compressDataVec_hitReq_27_51 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h33;
  wire         compressDataVec_hitReq_28_51 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h33;
  wire         compressDataVec_hitReq_29_51 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h33;
  wire         compressDataVec_hitReq_30_51 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h33;
  wire         compressDataVec_hitReq_31_51 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h33;
  wire [7:0]   compressDataVec_selectReqData_51 =
    (compressDataVec_hitReq_0_51 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_51 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_51 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_51 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_51 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_51 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_51 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_51 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_51 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_51 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_51 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_51 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_51 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_51 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_51 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_51 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_51 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_51 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_51 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_51 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_51 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_51 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_51 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_51 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_51 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_51 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_51 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_51 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_51 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_51 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_51 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_51 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_52 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h34;
  wire         compressDataVec_hitReq_1_52 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h34;
  wire         compressDataVec_hitReq_2_52 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h34;
  wire         compressDataVec_hitReq_3_52 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h34;
  wire         compressDataVec_hitReq_4_52 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h34;
  wire         compressDataVec_hitReq_5_52 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h34;
  wire         compressDataVec_hitReq_6_52 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h34;
  wire         compressDataVec_hitReq_7_52 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h34;
  wire         compressDataVec_hitReq_8_52 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h34;
  wire         compressDataVec_hitReq_9_52 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h34;
  wire         compressDataVec_hitReq_10_52 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h34;
  wire         compressDataVec_hitReq_11_52 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h34;
  wire         compressDataVec_hitReq_12_52 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h34;
  wire         compressDataVec_hitReq_13_52 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h34;
  wire         compressDataVec_hitReq_14_52 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h34;
  wire         compressDataVec_hitReq_15_52 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h34;
  wire         compressDataVec_hitReq_16_52 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h34;
  wire         compressDataVec_hitReq_17_52 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h34;
  wire         compressDataVec_hitReq_18_52 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h34;
  wire         compressDataVec_hitReq_19_52 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h34;
  wire         compressDataVec_hitReq_20_52 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h34;
  wire         compressDataVec_hitReq_21_52 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h34;
  wire         compressDataVec_hitReq_22_52 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h34;
  wire         compressDataVec_hitReq_23_52 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h34;
  wire         compressDataVec_hitReq_24_52 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h34;
  wire         compressDataVec_hitReq_25_52 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h34;
  wire         compressDataVec_hitReq_26_52 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h34;
  wire         compressDataVec_hitReq_27_52 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h34;
  wire         compressDataVec_hitReq_28_52 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h34;
  wire         compressDataVec_hitReq_29_52 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h34;
  wire         compressDataVec_hitReq_30_52 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h34;
  wire         compressDataVec_hitReq_31_52 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h34;
  wire [7:0]   compressDataVec_selectReqData_52 =
    (compressDataVec_hitReq_0_52 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_52 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_52 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_52 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_52 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_52 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_52 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_52 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_52 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_52 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_52 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_52 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_52 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_52 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_52 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_52 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_52 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_52 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_52 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_52 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_52 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_52 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_52 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_52 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_52 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_52 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_52 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_52 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_52 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_52 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_52 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_52 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_53 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h35;
  wire         compressDataVec_hitReq_1_53 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h35;
  wire         compressDataVec_hitReq_2_53 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h35;
  wire         compressDataVec_hitReq_3_53 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h35;
  wire         compressDataVec_hitReq_4_53 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h35;
  wire         compressDataVec_hitReq_5_53 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h35;
  wire         compressDataVec_hitReq_6_53 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h35;
  wire         compressDataVec_hitReq_7_53 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h35;
  wire         compressDataVec_hitReq_8_53 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h35;
  wire         compressDataVec_hitReq_9_53 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h35;
  wire         compressDataVec_hitReq_10_53 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h35;
  wire         compressDataVec_hitReq_11_53 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h35;
  wire         compressDataVec_hitReq_12_53 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h35;
  wire         compressDataVec_hitReq_13_53 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h35;
  wire         compressDataVec_hitReq_14_53 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h35;
  wire         compressDataVec_hitReq_15_53 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h35;
  wire         compressDataVec_hitReq_16_53 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h35;
  wire         compressDataVec_hitReq_17_53 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h35;
  wire         compressDataVec_hitReq_18_53 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h35;
  wire         compressDataVec_hitReq_19_53 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h35;
  wire         compressDataVec_hitReq_20_53 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h35;
  wire         compressDataVec_hitReq_21_53 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h35;
  wire         compressDataVec_hitReq_22_53 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h35;
  wire         compressDataVec_hitReq_23_53 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h35;
  wire         compressDataVec_hitReq_24_53 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h35;
  wire         compressDataVec_hitReq_25_53 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h35;
  wire         compressDataVec_hitReq_26_53 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h35;
  wire         compressDataVec_hitReq_27_53 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h35;
  wire         compressDataVec_hitReq_28_53 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h35;
  wire         compressDataVec_hitReq_29_53 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h35;
  wire         compressDataVec_hitReq_30_53 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h35;
  wire         compressDataVec_hitReq_31_53 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h35;
  wire [7:0]   compressDataVec_selectReqData_53 =
    (compressDataVec_hitReq_0_53 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_53 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_53 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_53 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_53 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_53 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_53 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_53 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_53 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_53 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_53 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_53 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_53 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_53 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_53 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_53 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_53 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_53 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_53 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_53 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_53 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_53 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_53 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_53 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_53 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_53 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_53 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_53 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_53 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_53 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_53 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_53 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_54 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h36;
  wire         compressDataVec_hitReq_1_54 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h36;
  wire         compressDataVec_hitReq_2_54 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h36;
  wire         compressDataVec_hitReq_3_54 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h36;
  wire         compressDataVec_hitReq_4_54 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h36;
  wire         compressDataVec_hitReq_5_54 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h36;
  wire         compressDataVec_hitReq_6_54 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h36;
  wire         compressDataVec_hitReq_7_54 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h36;
  wire         compressDataVec_hitReq_8_54 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h36;
  wire         compressDataVec_hitReq_9_54 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h36;
  wire         compressDataVec_hitReq_10_54 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h36;
  wire         compressDataVec_hitReq_11_54 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h36;
  wire         compressDataVec_hitReq_12_54 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h36;
  wire         compressDataVec_hitReq_13_54 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h36;
  wire         compressDataVec_hitReq_14_54 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h36;
  wire         compressDataVec_hitReq_15_54 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h36;
  wire         compressDataVec_hitReq_16_54 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h36;
  wire         compressDataVec_hitReq_17_54 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h36;
  wire         compressDataVec_hitReq_18_54 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h36;
  wire         compressDataVec_hitReq_19_54 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h36;
  wire         compressDataVec_hitReq_20_54 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h36;
  wire         compressDataVec_hitReq_21_54 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h36;
  wire         compressDataVec_hitReq_22_54 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h36;
  wire         compressDataVec_hitReq_23_54 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h36;
  wire         compressDataVec_hitReq_24_54 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h36;
  wire         compressDataVec_hitReq_25_54 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h36;
  wire         compressDataVec_hitReq_26_54 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h36;
  wire         compressDataVec_hitReq_27_54 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h36;
  wire         compressDataVec_hitReq_28_54 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h36;
  wire         compressDataVec_hitReq_29_54 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h36;
  wire         compressDataVec_hitReq_30_54 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h36;
  wire         compressDataVec_hitReq_31_54 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h36;
  wire [7:0]   compressDataVec_selectReqData_54 =
    (compressDataVec_hitReq_0_54 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_54 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_54 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_54 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_54 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_54 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_54 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_54 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_54 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_54 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_54 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_54 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_54 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_54 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_54 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_54 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_54 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_54 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_54 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_54 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_54 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_54 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_54 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_54 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_54 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_54 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_54 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_54 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_54 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_54 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_54 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_54 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_55 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h37;
  wire         compressDataVec_hitReq_1_55 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h37;
  wire         compressDataVec_hitReq_2_55 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h37;
  wire         compressDataVec_hitReq_3_55 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h37;
  wire         compressDataVec_hitReq_4_55 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h37;
  wire         compressDataVec_hitReq_5_55 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h37;
  wire         compressDataVec_hitReq_6_55 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h37;
  wire         compressDataVec_hitReq_7_55 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h37;
  wire         compressDataVec_hitReq_8_55 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h37;
  wire         compressDataVec_hitReq_9_55 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h37;
  wire         compressDataVec_hitReq_10_55 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h37;
  wire         compressDataVec_hitReq_11_55 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h37;
  wire         compressDataVec_hitReq_12_55 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h37;
  wire         compressDataVec_hitReq_13_55 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h37;
  wire         compressDataVec_hitReq_14_55 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h37;
  wire         compressDataVec_hitReq_15_55 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h37;
  wire         compressDataVec_hitReq_16_55 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h37;
  wire         compressDataVec_hitReq_17_55 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h37;
  wire         compressDataVec_hitReq_18_55 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h37;
  wire         compressDataVec_hitReq_19_55 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h37;
  wire         compressDataVec_hitReq_20_55 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h37;
  wire         compressDataVec_hitReq_21_55 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h37;
  wire         compressDataVec_hitReq_22_55 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h37;
  wire         compressDataVec_hitReq_23_55 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h37;
  wire         compressDataVec_hitReq_24_55 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h37;
  wire         compressDataVec_hitReq_25_55 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h37;
  wire         compressDataVec_hitReq_26_55 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h37;
  wire         compressDataVec_hitReq_27_55 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h37;
  wire         compressDataVec_hitReq_28_55 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h37;
  wire         compressDataVec_hitReq_29_55 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h37;
  wire         compressDataVec_hitReq_30_55 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h37;
  wire         compressDataVec_hitReq_31_55 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h37;
  wire [7:0]   compressDataVec_selectReqData_55 =
    (compressDataVec_hitReq_0_55 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_55 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_55 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_55 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_55 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_55 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_55 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_55 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_55 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_55 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_55 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_55 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_55 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_55 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_55 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_55 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_55 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_55 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_55 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_55 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_55 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_55 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_55 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_55 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_55 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_55 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_55 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_55 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_55 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_55 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_55 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_55 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_56 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h38;
  wire         compressDataVec_hitReq_1_56 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h38;
  wire         compressDataVec_hitReq_2_56 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h38;
  wire         compressDataVec_hitReq_3_56 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h38;
  wire         compressDataVec_hitReq_4_56 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h38;
  wire         compressDataVec_hitReq_5_56 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h38;
  wire         compressDataVec_hitReq_6_56 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h38;
  wire         compressDataVec_hitReq_7_56 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h38;
  wire         compressDataVec_hitReq_8_56 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h38;
  wire         compressDataVec_hitReq_9_56 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h38;
  wire         compressDataVec_hitReq_10_56 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h38;
  wire         compressDataVec_hitReq_11_56 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h38;
  wire         compressDataVec_hitReq_12_56 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h38;
  wire         compressDataVec_hitReq_13_56 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h38;
  wire         compressDataVec_hitReq_14_56 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h38;
  wire         compressDataVec_hitReq_15_56 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h38;
  wire         compressDataVec_hitReq_16_56 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h38;
  wire         compressDataVec_hitReq_17_56 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h38;
  wire         compressDataVec_hitReq_18_56 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h38;
  wire         compressDataVec_hitReq_19_56 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h38;
  wire         compressDataVec_hitReq_20_56 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h38;
  wire         compressDataVec_hitReq_21_56 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h38;
  wire         compressDataVec_hitReq_22_56 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h38;
  wire         compressDataVec_hitReq_23_56 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h38;
  wire         compressDataVec_hitReq_24_56 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h38;
  wire         compressDataVec_hitReq_25_56 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h38;
  wire         compressDataVec_hitReq_26_56 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h38;
  wire         compressDataVec_hitReq_27_56 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h38;
  wire         compressDataVec_hitReq_28_56 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h38;
  wire         compressDataVec_hitReq_29_56 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h38;
  wire         compressDataVec_hitReq_30_56 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h38;
  wire         compressDataVec_hitReq_31_56 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h38;
  wire [7:0]   compressDataVec_selectReqData_56 =
    (compressDataVec_hitReq_0_56 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_56 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_56 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_56 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_56 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_56 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_56 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_56 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_56 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_56 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_56 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_56 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_56 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_56 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_56 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_56 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_56 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_56 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_56 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_56 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_56 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_56 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_56 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_56 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_56 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_56 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_56 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_56 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_56 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_56 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_56 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_56 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_57 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h39;
  wire         compressDataVec_hitReq_1_57 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h39;
  wire         compressDataVec_hitReq_2_57 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h39;
  wire         compressDataVec_hitReq_3_57 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h39;
  wire         compressDataVec_hitReq_4_57 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h39;
  wire         compressDataVec_hitReq_5_57 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h39;
  wire         compressDataVec_hitReq_6_57 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h39;
  wire         compressDataVec_hitReq_7_57 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h39;
  wire         compressDataVec_hitReq_8_57 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h39;
  wire         compressDataVec_hitReq_9_57 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h39;
  wire         compressDataVec_hitReq_10_57 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h39;
  wire         compressDataVec_hitReq_11_57 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h39;
  wire         compressDataVec_hitReq_12_57 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h39;
  wire         compressDataVec_hitReq_13_57 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h39;
  wire         compressDataVec_hitReq_14_57 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h39;
  wire         compressDataVec_hitReq_15_57 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h39;
  wire         compressDataVec_hitReq_16_57 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h39;
  wire         compressDataVec_hitReq_17_57 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h39;
  wire         compressDataVec_hitReq_18_57 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h39;
  wire         compressDataVec_hitReq_19_57 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h39;
  wire         compressDataVec_hitReq_20_57 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h39;
  wire         compressDataVec_hitReq_21_57 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h39;
  wire         compressDataVec_hitReq_22_57 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h39;
  wire         compressDataVec_hitReq_23_57 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h39;
  wire         compressDataVec_hitReq_24_57 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h39;
  wire         compressDataVec_hitReq_25_57 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h39;
  wire         compressDataVec_hitReq_26_57 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h39;
  wire         compressDataVec_hitReq_27_57 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h39;
  wire         compressDataVec_hitReq_28_57 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h39;
  wire         compressDataVec_hitReq_29_57 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h39;
  wire         compressDataVec_hitReq_30_57 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h39;
  wire         compressDataVec_hitReq_31_57 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h39;
  wire [7:0]   compressDataVec_selectReqData_57 =
    (compressDataVec_hitReq_0_57 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_57 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_57 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_57 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_57 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_57 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_57 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_57 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_57 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_57 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_57 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_57 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_57 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_57 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_57 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_57 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_57 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_57 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_57 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_57 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_57 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_57 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_57 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_57 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_57 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_57 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_57 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_57 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_57 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_57 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_57 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_57 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_58 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3A;
  wire         compressDataVec_hitReq_1_58 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3A;
  wire         compressDataVec_hitReq_2_58 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3A;
  wire         compressDataVec_hitReq_3_58 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3A;
  wire         compressDataVec_hitReq_4_58 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3A;
  wire         compressDataVec_hitReq_5_58 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3A;
  wire         compressDataVec_hitReq_6_58 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3A;
  wire         compressDataVec_hitReq_7_58 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3A;
  wire         compressDataVec_hitReq_8_58 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3A;
  wire         compressDataVec_hitReq_9_58 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3A;
  wire         compressDataVec_hitReq_10_58 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3A;
  wire         compressDataVec_hitReq_11_58 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3A;
  wire         compressDataVec_hitReq_12_58 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3A;
  wire         compressDataVec_hitReq_13_58 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3A;
  wire         compressDataVec_hitReq_14_58 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3A;
  wire         compressDataVec_hitReq_15_58 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3A;
  wire         compressDataVec_hitReq_16_58 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3A;
  wire         compressDataVec_hitReq_17_58 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3A;
  wire         compressDataVec_hitReq_18_58 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3A;
  wire         compressDataVec_hitReq_19_58 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3A;
  wire         compressDataVec_hitReq_20_58 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3A;
  wire         compressDataVec_hitReq_21_58 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3A;
  wire         compressDataVec_hitReq_22_58 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3A;
  wire         compressDataVec_hitReq_23_58 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3A;
  wire         compressDataVec_hitReq_24_58 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3A;
  wire         compressDataVec_hitReq_25_58 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3A;
  wire         compressDataVec_hitReq_26_58 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3A;
  wire         compressDataVec_hitReq_27_58 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3A;
  wire         compressDataVec_hitReq_28_58 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3A;
  wire         compressDataVec_hitReq_29_58 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3A;
  wire         compressDataVec_hitReq_30_58 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3A;
  wire         compressDataVec_hitReq_31_58 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3A;
  wire [7:0]   compressDataVec_selectReqData_58 =
    (compressDataVec_hitReq_0_58 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_58 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_58 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_58 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_58 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_58 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_58 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_58 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_58 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_58 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_58 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_58 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_58 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_58 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_58 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_58 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_58 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_58 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_58 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_58 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_58 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_58 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_58 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_58 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_58 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_58 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_58 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_58 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_58 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_58 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_58 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_58 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_59 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3B;
  wire         compressDataVec_hitReq_1_59 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3B;
  wire         compressDataVec_hitReq_2_59 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3B;
  wire         compressDataVec_hitReq_3_59 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3B;
  wire         compressDataVec_hitReq_4_59 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3B;
  wire         compressDataVec_hitReq_5_59 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3B;
  wire         compressDataVec_hitReq_6_59 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3B;
  wire         compressDataVec_hitReq_7_59 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3B;
  wire         compressDataVec_hitReq_8_59 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3B;
  wire         compressDataVec_hitReq_9_59 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3B;
  wire         compressDataVec_hitReq_10_59 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3B;
  wire         compressDataVec_hitReq_11_59 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3B;
  wire         compressDataVec_hitReq_12_59 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3B;
  wire         compressDataVec_hitReq_13_59 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3B;
  wire         compressDataVec_hitReq_14_59 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3B;
  wire         compressDataVec_hitReq_15_59 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3B;
  wire         compressDataVec_hitReq_16_59 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3B;
  wire         compressDataVec_hitReq_17_59 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3B;
  wire         compressDataVec_hitReq_18_59 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3B;
  wire         compressDataVec_hitReq_19_59 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3B;
  wire         compressDataVec_hitReq_20_59 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3B;
  wire         compressDataVec_hitReq_21_59 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3B;
  wire         compressDataVec_hitReq_22_59 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3B;
  wire         compressDataVec_hitReq_23_59 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3B;
  wire         compressDataVec_hitReq_24_59 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3B;
  wire         compressDataVec_hitReq_25_59 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3B;
  wire         compressDataVec_hitReq_26_59 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3B;
  wire         compressDataVec_hitReq_27_59 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3B;
  wire         compressDataVec_hitReq_28_59 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3B;
  wire         compressDataVec_hitReq_29_59 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3B;
  wire         compressDataVec_hitReq_30_59 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3B;
  wire         compressDataVec_hitReq_31_59 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3B;
  wire [7:0]   compressDataVec_selectReqData_59 =
    (compressDataVec_hitReq_0_59 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_59 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_59 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_59 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_59 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_59 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_59 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_59 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_59 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_59 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_59 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_59 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_59 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_59 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_59 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_59 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_59 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_59 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_59 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_59 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_59 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_59 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_59 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_59 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_59 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_59 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_59 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_59 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_59 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_59 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_59 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_59 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_60 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3C;
  wire         compressDataVec_hitReq_1_60 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3C;
  wire         compressDataVec_hitReq_2_60 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3C;
  wire         compressDataVec_hitReq_3_60 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3C;
  wire         compressDataVec_hitReq_4_60 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3C;
  wire         compressDataVec_hitReq_5_60 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3C;
  wire         compressDataVec_hitReq_6_60 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3C;
  wire         compressDataVec_hitReq_7_60 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3C;
  wire         compressDataVec_hitReq_8_60 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3C;
  wire         compressDataVec_hitReq_9_60 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3C;
  wire         compressDataVec_hitReq_10_60 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3C;
  wire         compressDataVec_hitReq_11_60 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3C;
  wire         compressDataVec_hitReq_12_60 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3C;
  wire         compressDataVec_hitReq_13_60 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3C;
  wire         compressDataVec_hitReq_14_60 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3C;
  wire         compressDataVec_hitReq_15_60 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3C;
  wire         compressDataVec_hitReq_16_60 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3C;
  wire         compressDataVec_hitReq_17_60 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3C;
  wire         compressDataVec_hitReq_18_60 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3C;
  wire         compressDataVec_hitReq_19_60 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3C;
  wire         compressDataVec_hitReq_20_60 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3C;
  wire         compressDataVec_hitReq_21_60 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3C;
  wire         compressDataVec_hitReq_22_60 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3C;
  wire         compressDataVec_hitReq_23_60 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3C;
  wire         compressDataVec_hitReq_24_60 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3C;
  wire         compressDataVec_hitReq_25_60 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3C;
  wire         compressDataVec_hitReq_26_60 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3C;
  wire         compressDataVec_hitReq_27_60 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3C;
  wire         compressDataVec_hitReq_28_60 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3C;
  wire         compressDataVec_hitReq_29_60 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3C;
  wire         compressDataVec_hitReq_30_60 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3C;
  wire         compressDataVec_hitReq_31_60 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3C;
  wire [7:0]   compressDataVec_selectReqData_60 =
    (compressDataVec_hitReq_0_60 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_60 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_60 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_60 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_60 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_60 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_60 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_60 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_60 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_60 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_60 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_60 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_60 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_60 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_60 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_60 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_60 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_60 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_60 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_60 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_60 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_60 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_60 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_60 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_60 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_60 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_60 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_60 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_60 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_60 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_60 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_60 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_61 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3D;
  wire         compressDataVec_hitReq_1_61 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3D;
  wire         compressDataVec_hitReq_2_61 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3D;
  wire         compressDataVec_hitReq_3_61 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3D;
  wire         compressDataVec_hitReq_4_61 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3D;
  wire         compressDataVec_hitReq_5_61 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3D;
  wire         compressDataVec_hitReq_6_61 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3D;
  wire         compressDataVec_hitReq_7_61 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3D;
  wire         compressDataVec_hitReq_8_61 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3D;
  wire         compressDataVec_hitReq_9_61 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3D;
  wire         compressDataVec_hitReq_10_61 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3D;
  wire         compressDataVec_hitReq_11_61 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3D;
  wire         compressDataVec_hitReq_12_61 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3D;
  wire         compressDataVec_hitReq_13_61 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3D;
  wire         compressDataVec_hitReq_14_61 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3D;
  wire         compressDataVec_hitReq_15_61 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3D;
  wire         compressDataVec_hitReq_16_61 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3D;
  wire         compressDataVec_hitReq_17_61 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3D;
  wire         compressDataVec_hitReq_18_61 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3D;
  wire         compressDataVec_hitReq_19_61 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3D;
  wire         compressDataVec_hitReq_20_61 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3D;
  wire         compressDataVec_hitReq_21_61 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3D;
  wire         compressDataVec_hitReq_22_61 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3D;
  wire         compressDataVec_hitReq_23_61 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3D;
  wire         compressDataVec_hitReq_24_61 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3D;
  wire         compressDataVec_hitReq_25_61 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3D;
  wire         compressDataVec_hitReq_26_61 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3D;
  wire         compressDataVec_hitReq_27_61 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3D;
  wire         compressDataVec_hitReq_28_61 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3D;
  wire         compressDataVec_hitReq_29_61 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3D;
  wire         compressDataVec_hitReq_30_61 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3D;
  wire         compressDataVec_hitReq_31_61 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3D;
  wire [7:0]   compressDataVec_selectReqData_61 =
    (compressDataVec_hitReq_0_61 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_61 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_61 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_61 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_61 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_61 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_61 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_61 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_61 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_61 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_61 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_61 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_61 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_61 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_61 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_61 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_61 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_61 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_61 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_61 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_61 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_61 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_61 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_61 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_61 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_61 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_61 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_61 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_61 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_61 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_61 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_61 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_62 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3E;
  wire         compressDataVec_hitReq_1_62 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3E;
  wire         compressDataVec_hitReq_2_62 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3E;
  wire         compressDataVec_hitReq_3_62 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3E;
  wire         compressDataVec_hitReq_4_62 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3E;
  wire         compressDataVec_hitReq_5_62 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3E;
  wire         compressDataVec_hitReq_6_62 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3E;
  wire         compressDataVec_hitReq_7_62 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3E;
  wire         compressDataVec_hitReq_8_62 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3E;
  wire         compressDataVec_hitReq_9_62 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3E;
  wire         compressDataVec_hitReq_10_62 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3E;
  wire         compressDataVec_hitReq_11_62 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3E;
  wire         compressDataVec_hitReq_12_62 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3E;
  wire         compressDataVec_hitReq_13_62 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3E;
  wire         compressDataVec_hitReq_14_62 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3E;
  wire         compressDataVec_hitReq_15_62 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3E;
  wire         compressDataVec_hitReq_16_62 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3E;
  wire         compressDataVec_hitReq_17_62 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3E;
  wire         compressDataVec_hitReq_18_62 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3E;
  wire         compressDataVec_hitReq_19_62 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3E;
  wire         compressDataVec_hitReq_20_62 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3E;
  wire         compressDataVec_hitReq_21_62 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3E;
  wire         compressDataVec_hitReq_22_62 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3E;
  wire         compressDataVec_hitReq_23_62 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3E;
  wire         compressDataVec_hitReq_24_62 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3E;
  wire         compressDataVec_hitReq_25_62 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3E;
  wire         compressDataVec_hitReq_26_62 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3E;
  wire         compressDataVec_hitReq_27_62 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3E;
  wire         compressDataVec_hitReq_28_62 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3E;
  wire         compressDataVec_hitReq_29_62 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3E;
  wire         compressDataVec_hitReq_30_62 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3E;
  wire         compressDataVec_hitReq_31_62 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3E;
  wire [7:0]   compressDataVec_selectReqData_62 =
    (compressDataVec_hitReq_0_62 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_62 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_62 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_62 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_62 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_62 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_62 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_62 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_62 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_62 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_62 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_62 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_62 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_62 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_62 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_62 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_62 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_62 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_62 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_62 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_62 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_62 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_62 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_62 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_62 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_62 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_62 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_62 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_62 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_62 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_62 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_62 ? source2Pipe[255:248] : 8'h0);
  wire         compressDataVec_hitReq_0_63 = compressMaskVecPipe_0 & compressVecPipe_0 == 10'h3F;
  wire         compressDataVec_hitReq_1_63 = compressMaskVecPipe_1 & compressVecPipe_1 == 10'h3F;
  wire         compressDataVec_hitReq_2_63 = compressMaskVecPipe_2 & compressVecPipe_2 == 10'h3F;
  wire         compressDataVec_hitReq_3_63 = compressMaskVecPipe_3 & compressVecPipe_3 == 10'h3F;
  wire         compressDataVec_hitReq_4_63 = compressMaskVecPipe_4 & compressVecPipe_4 == 10'h3F;
  wire         compressDataVec_hitReq_5_63 = compressMaskVecPipe_5 & compressVecPipe_5 == 10'h3F;
  wire         compressDataVec_hitReq_6_63 = compressMaskVecPipe_6 & compressVecPipe_6 == 10'h3F;
  wire         compressDataVec_hitReq_7_63 = compressMaskVecPipe_7 & compressVecPipe_7 == 10'h3F;
  wire         compressDataVec_hitReq_8_63 = compressMaskVecPipe_8 & compressVecPipe_8 == 10'h3F;
  wire         compressDataVec_hitReq_9_63 = compressMaskVecPipe_9 & compressVecPipe_9 == 10'h3F;
  wire         compressDataVec_hitReq_10_63 = compressMaskVecPipe_10 & compressVecPipe_10 == 10'h3F;
  wire         compressDataVec_hitReq_11_63 = compressMaskVecPipe_11 & compressVecPipe_11 == 10'h3F;
  wire         compressDataVec_hitReq_12_63 = compressMaskVecPipe_12 & compressVecPipe_12 == 10'h3F;
  wire         compressDataVec_hitReq_13_63 = compressMaskVecPipe_13 & compressVecPipe_13 == 10'h3F;
  wire         compressDataVec_hitReq_14_63 = compressMaskVecPipe_14 & compressVecPipe_14 == 10'h3F;
  wire         compressDataVec_hitReq_15_63 = compressMaskVecPipe_15 & compressVecPipe_15 == 10'h3F;
  wire         compressDataVec_hitReq_16_63 = compressMaskVecPipe_16 & compressVecPipe_16 == 10'h3F;
  wire         compressDataVec_hitReq_17_63 = compressMaskVecPipe_17 & compressVecPipe_17 == 10'h3F;
  wire         compressDataVec_hitReq_18_63 = compressMaskVecPipe_18 & compressVecPipe_18 == 10'h3F;
  wire         compressDataVec_hitReq_19_63 = compressMaskVecPipe_19 & compressVecPipe_19 == 10'h3F;
  wire         compressDataVec_hitReq_20_63 = compressMaskVecPipe_20 & compressVecPipe_20 == 10'h3F;
  wire         compressDataVec_hitReq_21_63 = compressMaskVecPipe_21 & compressVecPipe_21 == 10'h3F;
  wire         compressDataVec_hitReq_22_63 = compressMaskVecPipe_22 & compressVecPipe_22 == 10'h3F;
  wire         compressDataVec_hitReq_23_63 = compressMaskVecPipe_23 & compressVecPipe_23 == 10'h3F;
  wire         compressDataVec_hitReq_24_63 = compressMaskVecPipe_24 & compressVecPipe_24 == 10'h3F;
  wire         compressDataVec_hitReq_25_63 = compressMaskVecPipe_25 & compressVecPipe_25 == 10'h3F;
  wire         compressDataVec_hitReq_26_63 = compressMaskVecPipe_26 & compressVecPipe_26 == 10'h3F;
  wire         compressDataVec_hitReq_27_63 = compressMaskVecPipe_27 & compressVecPipe_27 == 10'h3F;
  wire         compressDataVec_hitReq_28_63 = compressMaskVecPipe_28 & compressVecPipe_28 == 10'h3F;
  wire         compressDataVec_hitReq_29_63 = compressMaskVecPipe_29 & compressVecPipe_29 == 10'h3F;
  wire         compressDataVec_hitReq_30_63 = compressMaskVecPipe_30 & compressVecPipe_30 == 10'h3F;
  wire         compressDataVec_hitReq_31_63 = compressMaskVecPipe_31 & compressVecPipe_31 == 10'h3F;
  wire [7:0]   compressDataVec_selectReqData_63 =
    (compressDataVec_hitReq_0_63 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_63 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_63 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_63 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_63 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_63 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_63 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_63 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_63 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_63 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_63 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_63 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_63 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_63 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_63 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_63 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_63 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_63 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_63 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_63 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_63 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_63 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_63 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_63 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_63 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_63 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_63 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_63 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_63 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_63 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_63 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_63 ? source2Pipe[255:248] : 8'h0);
  wire [15:0]  compressDataVec_lo_lo_lo_lo_lo = {compressDataVec_useTail_1 ? compressDataReg[15:8] : compressDataVec_selectReqData_1, compressDataVec_useTail ? compressDataReg[7:0] : compressDataVec_selectReqData};
  wire [15:0]  compressDataVec_lo_lo_lo_lo_hi = {compressDataVec_useTail_3 ? compressDataReg[31:24] : compressDataVec_selectReqData_3, compressDataVec_useTail_2 ? compressDataReg[23:16] : compressDataVec_selectReqData_2};
  wire [31:0]  compressDataVec_lo_lo_lo_lo = {compressDataVec_lo_lo_lo_lo_hi, compressDataVec_lo_lo_lo_lo_lo};
  wire [15:0]  compressDataVec_lo_lo_lo_hi_lo = {compressDataVec_useTail_5 ? compressDataReg[47:40] : compressDataVec_selectReqData_5, compressDataVec_useTail_4 ? compressDataReg[39:32] : compressDataVec_selectReqData_4};
  wire [15:0]  compressDataVec_lo_lo_lo_hi_hi = {compressDataVec_useTail_7 ? compressDataReg[63:56] : compressDataVec_selectReqData_7, compressDataVec_useTail_6 ? compressDataReg[55:48] : compressDataVec_selectReqData_6};
  wire [31:0]  compressDataVec_lo_lo_lo_hi = {compressDataVec_lo_lo_lo_hi_hi, compressDataVec_lo_lo_lo_hi_lo};
  wire [63:0]  compressDataVec_lo_lo_lo = {compressDataVec_lo_lo_lo_hi, compressDataVec_lo_lo_lo_lo};
  wire [15:0]  compressDataVec_lo_lo_hi_lo_lo = {compressDataVec_useTail_9 ? compressDataReg[79:72] : compressDataVec_selectReqData_9, compressDataVec_useTail_8 ? compressDataReg[71:64] : compressDataVec_selectReqData_8};
  wire [15:0]  compressDataVec_lo_lo_hi_lo_hi = {compressDataVec_useTail_11 ? compressDataReg[95:88] : compressDataVec_selectReqData_11, compressDataVec_useTail_10 ? compressDataReg[87:80] : compressDataVec_selectReqData_10};
  wire [31:0]  compressDataVec_lo_lo_hi_lo = {compressDataVec_lo_lo_hi_lo_hi, compressDataVec_lo_lo_hi_lo_lo};
  wire [15:0]  compressDataVec_lo_lo_hi_hi_lo = {compressDataVec_useTail_13 ? compressDataReg[111:104] : compressDataVec_selectReqData_13, compressDataVec_useTail_12 ? compressDataReg[103:96] : compressDataVec_selectReqData_12};
  wire [15:0]  compressDataVec_lo_lo_hi_hi_hi = {compressDataVec_useTail_15 ? compressDataReg[127:120] : compressDataVec_selectReqData_15, compressDataVec_useTail_14 ? compressDataReg[119:112] : compressDataVec_selectReqData_14};
  wire [31:0]  compressDataVec_lo_lo_hi_hi = {compressDataVec_lo_lo_hi_hi_hi, compressDataVec_lo_lo_hi_hi_lo};
  wire [63:0]  compressDataVec_lo_lo_hi = {compressDataVec_lo_lo_hi_hi, compressDataVec_lo_lo_hi_lo};
  wire [127:0] compressDataVec_lo_lo = {compressDataVec_lo_lo_hi, compressDataVec_lo_lo_lo};
  wire [15:0]  compressDataVec_lo_hi_lo_lo_lo = {compressDataVec_useTail_17 ? compressDataReg[143:136] : compressDataVec_selectReqData_17, compressDataVec_useTail_16 ? compressDataReg[135:128] : compressDataVec_selectReqData_16};
  wire [15:0]  compressDataVec_lo_hi_lo_lo_hi = {compressDataVec_useTail_19 ? compressDataReg[159:152] : compressDataVec_selectReqData_19, compressDataVec_useTail_18 ? compressDataReg[151:144] : compressDataVec_selectReqData_18};
  wire [31:0]  compressDataVec_lo_hi_lo_lo = {compressDataVec_lo_hi_lo_lo_hi, compressDataVec_lo_hi_lo_lo_lo};
  wire [15:0]  compressDataVec_lo_hi_lo_hi_lo = {compressDataVec_useTail_21 ? compressDataReg[175:168] : compressDataVec_selectReqData_21, compressDataVec_useTail_20 ? compressDataReg[167:160] : compressDataVec_selectReqData_20};
  wire [15:0]  compressDataVec_lo_hi_lo_hi_hi = {compressDataVec_useTail_23 ? compressDataReg[191:184] : compressDataVec_selectReqData_23, compressDataVec_useTail_22 ? compressDataReg[183:176] : compressDataVec_selectReqData_22};
  wire [31:0]  compressDataVec_lo_hi_lo_hi = {compressDataVec_lo_hi_lo_hi_hi, compressDataVec_lo_hi_lo_hi_lo};
  wire [63:0]  compressDataVec_lo_hi_lo = {compressDataVec_lo_hi_lo_hi, compressDataVec_lo_hi_lo_lo};
  wire [15:0]  compressDataVec_lo_hi_hi_lo_lo = {compressDataVec_useTail_25 ? compressDataReg[207:200] : compressDataVec_selectReqData_25, compressDataVec_useTail_24 ? compressDataReg[199:192] : compressDataVec_selectReqData_24};
  wire [15:0]  compressDataVec_lo_hi_hi_lo_hi = {compressDataVec_useTail_27 ? compressDataReg[223:216] : compressDataVec_selectReqData_27, compressDataVec_useTail_26 ? compressDataReg[215:208] : compressDataVec_selectReqData_26};
  wire [31:0]  compressDataVec_lo_hi_hi_lo = {compressDataVec_lo_hi_hi_lo_hi, compressDataVec_lo_hi_hi_lo_lo};
  wire [15:0]  compressDataVec_lo_hi_hi_hi_lo = {compressDataVec_useTail_29 ? compressDataReg[239:232] : compressDataVec_selectReqData_29, compressDataVec_useTail_28 ? compressDataReg[231:224] : compressDataVec_selectReqData_28};
  wire [15:0]  compressDataVec_lo_hi_hi_hi_hi = {compressDataVec_selectReqData_31, compressDataVec_useTail_30 ? compressDataReg[247:240] : compressDataVec_selectReqData_30};
  wire [31:0]  compressDataVec_lo_hi_hi_hi = {compressDataVec_lo_hi_hi_hi_hi, compressDataVec_lo_hi_hi_hi_lo};
  wire [63:0]  compressDataVec_lo_hi_hi = {compressDataVec_lo_hi_hi_hi, compressDataVec_lo_hi_hi_lo};
  wire [127:0] compressDataVec_lo_hi = {compressDataVec_lo_hi_hi, compressDataVec_lo_hi_lo};
  wire [255:0] compressDataVec_lo = {compressDataVec_lo_hi, compressDataVec_lo_lo};
  wire [15:0]  compressDataVec_hi_lo_lo_lo_lo = {compressDataVec_selectReqData_33, compressDataVec_selectReqData_32};
  wire [15:0]  compressDataVec_hi_lo_lo_lo_hi = {compressDataVec_selectReqData_35, compressDataVec_selectReqData_34};
  wire [31:0]  compressDataVec_hi_lo_lo_lo = {compressDataVec_hi_lo_lo_lo_hi, compressDataVec_hi_lo_lo_lo_lo};
  wire [15:0]  compressDataVec_hi_lo_lo_hi_lo = {compressDataVec_selectReqData_37, compressDataVec_selectReqData_36};
  wire [15:0]  compressDataVec_hi_lo_lo_hi_hi = {compressDataVec_selectReqData_39, compressDataVec_selectReqData_38};
  wire [31:0]  compressDataVec_hi_lo_lo_hi = {compressDataVec_hi_lo_lo_hi_hi, compressDataVec_hi_lo_lo_hi_lo};
  wire [63:0]  compressDataVec_hi_lo_lo = {compressDataVec_hi_lo_lo_hi, compressDataVec_hi_lo_lo_lo};
  wire [15:0]  compressDataVec_hi_lo_hi_lo_lo = {compressDataVec_selectReqData_41, compressDataVec_selectReqData_40};
  wire [15:0]  compressDataVec_hi_lo_hi_lo_hi = {compressDataVec_selectReqData_43, compressDataVec_selectReqData_42};
  wire [31:0]  compressDataVec_hi_lo_hi_lo = {compressDataVec_hi_lo_hi_lo_hi, compressDataVec_hi_lo_hi_lo_lo};
  wire [15:0]  compressDataVec_hi_lo_hi_hi_lo = {compressDataVec_selectReqData_45, compressDataVec_selectReqData_44};
  wire [15:0]  compressDataVec_hi_lo_hi_hi_hi = {compressDataVec_selectReqData_47, compressDataVec_selectReqData_46};
  wire [31:0]  compressDataVec_hi_lo_hi_hi = {compressDataVec_hi_lo_hi_hi_hi, compressDataVec_hi_lo_hi_hi_lo};
  wire [63:0]  compressDataVec_hi_lo_hi = {compressDataVec_hi_lo_hi_hi, compressDataVec_hi_lo_hi_lo};
  wire [127:0] compressDataVec_hi_lo = {compressDataVec_hi_lo_hi, compressDataVec_hi_lo_lo};
  wire [15:0]  compressDataVec_hi_hi_lo_lo_lo = {compressDataVec_selectReqData_49, compressDataVec_selectReqData_48};
  wire [15:0]  compressDataVec_hi_hi_lo_lo_hi = {compressDataVec_selectReqData_51, compressDataVec_selectReqData_50};
  wire [31:0]  compressDataVec_hi_hi_lo_lo = {compressDataVec_hi_hi_lo_lo_hi, compressDataVec_hi_hi_lo_lo_lo};
  wire [15:0]  compressDataVec_hi_hi_lo_hi_lo = {compressDataVec_selectReqData_53, compressDataVec_selectReqData_52};
  wire [15:0]  compressDataVec_hi_hi_lo_hi_hi = {compressDataVec_selectReqData_55, compressDataVec_selectReqData_54};
  wire [31:0]  compressDataVec_hi_hi_lo_hi = {compressDataVec_hi_hi_lo_hi_hi, compressDataVec_hi_hi_lo_hi_lo};
  wire [63:0]  compressDataVec_hi_hi_lo = {compressDataVec_hi_hi_lo_hi, compressDataVec_hi_hi_lo_lo};
  wire [15:0]  compressDataVec_hi_hi_hi_lo_lo = {compressDataVec_selectReqData_57, compressDataVec_selectReqData_56};
  wire [15:0]  compressDataVec_hi_hi_hi_lo_hi = {compressDataVec_selectReqData_59, compressDataVec_selectReqData_58};
  wire [31:0]  compressDataVec_hi_hi_hi_lo = {compressDataVec_hi_hi_hi_lo_hi, compressDataVec_hi_hi_hi_lo_lo};
  wire [15:0]  compressDataVec_hi_hi_hi_hi_lo = {compressDataVec_selectReqData_61, compressDataVec_selectReqData_60};
  wire [15:0]  compressDataVec_hi_hi_hi_hi_hi = {compressDataVec_selectReqData_63, compressDataVec_selectReqData_62};
  wire [31:0]  compressDataVec_hi_hi_hi_hi = {compressDataVec_hi_hi_hi_hi_hi, compressDataVec_hi_hi_hi_hi_lo};
  wire [63:0]  compressDataVec_hi_hi_hi = {compressDataVec_hi_hi_hi_hi, compressDataVec_hi_hi_hi_lo};
  wire [127:0] compressDataVec_hi_hi = {compressDataVec_hi_hi_hi, compressDataVec_hi_hi_lo};
  wire [255:0] compressDataVec_hi = {compressDataVec_hi_hi, compressDataVec_hi_lo};
  wire [511:0] compressDataVec_0 = {compressDataVec_hi, compressDataVec_lo};
  wire [15:0]  compressDataVec_selectReqData_64 =
    (compressDataVec_hitReq_0_64 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_64 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_64 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_64 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_64 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_64 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_64 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_64 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_64 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_64 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_64 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_64 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_64 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_64 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_64 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_64 ? source2Pipe[255:240] : 16'h0);
  wire         compressDataVec_useTail_32;
  assign compressDataVec_useTail_32 = |tailCount;
  wire [15:0]  compressDataVec_selectReqData_65 =
    (compressDataVec_hitReq_0_65 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_65 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_65 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_65 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_65 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_65 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_65 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_65 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_65 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_65 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_65 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_65 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_65 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_65 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_65 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_65 ? source2Pipe[255:240] : 16'h0);
  wire         compressDataVec_useTail_33;
  assign compressDataVec_useTail_33 = |(tailCount[4:1]);
  wire [15:0]  compressDataVec_selectReqData_66 =
    (compressDataVec_hitReq_0_66 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_66 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_66 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_66 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_66 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_66 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_66 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_66 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_66 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_66 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_66 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_66 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_66 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_66 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_66 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_66 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_67 =
    (compressDataVec_hitReq_0_67 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_67 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_67 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_67 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_67 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_67 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_67 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_67 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_67 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_67 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_67 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_67 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_67 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_67 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_67 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_67 ? source2Pipe[255:240] : 16'h0);
  wire         compressDataVec_useTail_35;
  assign compressDataVec_useTail_35 = |(tailCount[4:2]);
  wire [15:0]  compressDataVec_selectReqData_68 =
    (compressDataVec_hitReq_0_68 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_68 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_68 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_68 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_68 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_68 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_68 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_68 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_68 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_68 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_68 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_68 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_68 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_68 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_68 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_68 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_69 =
    (compressDataVec_hitReq_0_69 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_69 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_69 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_69 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_69 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_69 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_69 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_69 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_69 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_69 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_69 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_69 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_69 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_69 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_69 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_69 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_70 =
    (compressDataVec_hitReq_0_70 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_70 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_70 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_70 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_70 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_70 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_70 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_70 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_70 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_70 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_70 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_70 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_70 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_70 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_70 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_70 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_71 =
    (compressDataVec_hitReq_0_71 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_71 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_71 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_71 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_71 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_71 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_71 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_71 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_71 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_71 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_71 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_71 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_71 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_71 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_71 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_71 ? source2Pipe[255:240] : 16'h0);
  wire         compressDataVec_useTail_39;
  assign compressDataVec_useTail_39 = |(tailCount[4:3]);
  wire [15:0]  compressDataVec_selectReqData_72 =
    (compressDataVec_hitReq_0_72 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_72 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_72 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_72 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_72 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_72 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_72 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_72 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_72 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_72 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_72 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_72 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_72 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_72 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_72 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_72 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_73 =
    (compressDataVec_hitReq_0_73 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_73 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_73 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_73 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_73 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_73 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_73 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_73 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_73 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_73 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_73 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_73 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_73 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_73 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_73 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_73 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_74 =
    (compressDataVec_hitReq_0_74 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_74 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_74 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_74 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_74 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_74 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_74 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_74 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_74 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_74 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_74 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_74 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_74 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_74 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_74 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_74 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_75 =
    (compressDataVec_hitReq_0_75 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_75 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_75 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_75 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_75 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_75 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_75 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_75 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_75 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_75 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_75 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_75 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_75 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_75 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_75 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_75 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_76 =
    (compressDataVec_hitReq_0_76 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_76 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_76 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_76 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_76 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_76 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_76 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_76 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_76 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_76 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_76 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_76 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_76 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_76 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_76 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_76 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_77 =
    (compressDataVec_hitReq_0_77 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_77 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_77 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_77 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_77 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_77 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_77 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_77 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_77 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_77 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_77 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_77 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_77 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_77 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_77 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_77 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_78 =
    (compressDataVec_hitReq_0_78 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_78 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_78 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_78 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_78 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_78 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_78 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_78 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_78 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_78 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_78 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_78 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_78 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_78 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_78 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_78 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_79 =
    (compressDataVec_hitReq_0_79 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_79 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_79 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_79 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_79 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_79 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_79 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_79 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_79 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_79 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_79 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_79 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_79 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_79 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_79 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_79 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_80 =
    (compressDataVec_hitReq_0_80 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_80 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_80 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_80 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_80 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_80 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_80 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_80 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_80 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_80 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_80 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_80 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_80 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_80 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_80 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_80 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_81 =
    (compressDataVec_hitReq_0_81 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_81 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_81 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_81 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_81 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_81 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_81 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_81 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_81 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_81 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_81 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_81 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_81 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_81 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_81 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_81 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_82 =
    (compressDataVec_hitReq_0_82 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_82 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_82 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_82 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_82 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_82 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_82 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_82 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_82 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_82 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_82 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_82 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_82 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_82 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_82 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_82 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_83 =
    (compressDataVec_hitReq_0_83 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_83 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_83 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_83 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_83 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_83 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_83 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_83 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_83 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_83 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_83 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_83 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_83 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_83 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_83 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_83 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_84 =
    (compressDataVec_hitReq_0_84 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_84 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_84 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_84 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_84 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_84 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_84 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_84 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_84 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_84 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_84 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_84 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_84 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_84 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_84 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_84 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_85 =
    (compressDataVec_hitReq_0_85 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_85 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_85 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_85 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_85 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_85 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_85 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_85 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_85 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_85 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_85 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_85 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_85 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_85 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_85 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_85 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_86 =
    (compressDataVec_hitReq_0_86 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_86 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_86 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_86 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_86 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_86 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_86 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_86 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_86 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_86 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_86 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_86 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_86 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_86 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_86 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_86 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_87 =
    (compressDataVec_hitReq_0_87 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_87 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_87 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_87 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_87 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_87 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_87 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_87 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_87 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_87 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_87 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_87 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_87 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_87 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_87 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_87 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_88 =
    (compressDataVec_hitReq_0_88 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_88 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_88 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_88 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_88 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_88 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_88 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_88 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_88 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_88 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_88 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_88 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_88 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_88 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_88 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_88 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_89 =
    (compressDataVec_hitReq_0_89 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_89 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_89 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_89 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_89 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_89 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_89 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_89 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_89 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_89 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_89 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_89 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_89 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_89 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_89 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_89 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_90 =
    (compressDataVec_hitReq_0_90 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_90 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_90 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_90 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_90 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_90 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_90 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_90 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_90 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_90 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_90 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_90 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_90 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_90 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_90 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_90 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_91 =
    (compressDataVec_hitReq_0_91 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_91 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_91 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_91 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_91 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_91 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_91 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_91 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_91 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_91 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_91 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_91 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_91 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_91 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_91 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_91 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_92 =
    (compressDataVec_hitReq_0_92 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_92 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_92 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_92 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_92 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_92 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_92 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_92 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_92 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_92 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_92 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_92 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_92 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_92 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_92 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_92 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_93 =
    (compressDataVec_hitReq_0_93 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_93 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_93 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_93 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_93 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_93 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_93 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_93 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_93 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_93 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_93 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_93 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_93 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_93 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_93 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_93 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_94 =
    (compressDataVec_hitReq_0_94 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_94 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_94 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_94 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_94 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_94 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_94 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_94 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_94 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_94 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_94 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_94 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_94 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_94 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_94 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_94 ? source2Pipe[255:240] : 16'h0);
  wire [15:0]  compressDataVec_selectReqData_95 =
    (compressDataVec_hitReq_0_95 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_95 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_95 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_95 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_95 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_95 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_95 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_95 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_95 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_95 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_95 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_95 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_95 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_95 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_95 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_95 ? source2Pipe[255:240] : 16'h0);
  wire [31:0]  compressDataVec_lo_lo_lo_lo_1 = {compressDataVec_useTail_33 ? compressDataReg[31:16] : compressDataVec_selectReqData_65, compressDataVec_useTail_32 ? compressDataReg[15:0] : compressDataVec_selectReqData_64};
  wire [31:0]  compressDataVec_lo_lo_lo_hi_1 = {compressDataVec_useTail_35 ? compressDataReg[63:48] : compressDataVec_selectReqData_67, compressDataVec_useTail_34 ? compressDataReg[47:32] : compressDataVec_selectReqData_66};
  wire [63:0]  compressDataVec_lo_lo_lo_1 = {compressDataVec_lo_lo_lo_hi_1, compressDataVec_lo_lo_lo_lo_1};
  wire [31:0]  compressDataVec_lo_lo_hi_lo_1 = {compressDataVec_useTail_37 ? compressDataReg[95:80] : compressDataVec_selectReqData_69, compressDataVec_useTail_36 ? compressDataReg[79:64] : compressDataVec_selectReqData_68};
  wire [31:0]  compressDataVec_lo_lo_hi_hi_1 = {compressDataVec_useTail_39 ? compressDataReg[127:112] : compressDataVec_selectReqData_71, compressDataVec_useTail_38 ? compressDataReg[111:96] : compressDataVec_selectReqData_70};
  wire [63:0]  compressDataVec_lo_lo_hi_1 = {compressDataVec_lo_lo_hi_hi_1, compressDataVec_lo_lo_hi_lo_1};
  wire [127:0] compressDataVec_lo_lo_1 = {compressDataVec_lo_lo_hi_1, compressDataVec_lo_lo_lo_1};
  wire [31:0]  compressDataVec_lo_hi_lo_lo_1 = {compressDataVec_useTail_41 ? compressDataReg[159:144] : compressDataVec_selectReqData_73, compressDataVec_useTail_40 ? compressDataReg[143:128] : compressDataVec_selectReqData_72};
  wire [31:0]  compressDataVec_lo_hi_lo_hi_1 = {compressDataVec_useTail_43 ? compressDataReg[191:176] : compressDataVec_selectReqData_75, compressDataVec_useTail_42 ? compressDataReg[175:160] : compressDataVec_selectReqData_74};
  wire [63:0]  compressDataVec_lo_hi_lo_1 = {compressDataVec_lo_hi_lo_hi_1, compressDataVec_lo_hi_lo_lo_1};
  wire [31:0]  compressDataVec_lo_hi_hi_lo_1 = {compressDataVec_useTail_45 ? compressDataReg[223:208] : compressDataVec_selectReqData_77, compressDataVec_useTail_44 ? compressDataReg[207:192] : compressDataVec_selectReqData_76};
  wire [31:0]  compressDataVec_lo_hi_hi_hi_1 = {compressDataVec_useTail_47 ? compressDataReg[255:240] : compressDataVec_selectReqData_79, compressDataVec_useTail_46 ? compressDataReg[239:224] : compressDataVec_selectReqData_78};
  wire [63:0]  compressDataVec_lo_hi_hi_1 = {compressDataVec_lo_hi_hi_hi_1, compressDataVec_lo_hi_hi_lo_1};
  wire [127:0] compressDataVec_lo_hi_1 = {compressDataVec_lo_hi_hi_1, compressDataVec_lo_hi_lo_1};
  wire [255:0] compressDataVec_lo_1 = {compressDataVec_lo_hi_1, compressDataVec_lo_lo_1};
  wire [31:0]  compressDataVec_hi_lo_lo_lo_1 = {compressDataVec_selectReqData_81, compressDataVec_selectReqData_80};
  wire [31:0]  compressDataVec_hi_lo_lo_hi_1 = {compressDataVec_selectReqData_83, compressDataVec_selectReqData_82};
  wire [63:0]  compressDataVec_hi_lo_lo_1 = {compressDataVec_hi_lo_lo_hi_1, compressDataVec_hi_lo_lo_lo_1};
  wire [31:0]  compressDataVec_hi_lo_hi_lo_1 = {compressDataVec_selectReqData_85, compressDataVec_selectReqData_84};
  wire [31:0]  compressDataVec_hi_lo_hi_hi_1 = {compressDataVec_selectReqData_87, compressDataVec_selectReqData_86};
  wire [63:0]  compressDataVec_hi_lo_hi_1 = {compressDataVec_hi_lo_hi_hi_1, compressDataVec_hi_lo_hi_lo_1};
  wire [127:0] compressDataVec_hi_lo_1 = {compressDataVec_hi_lo_hi_1, compressDataVec_hi_lo_lo_1};
  wire [31:0]  compressDataVec_hi_hi_lo_lo_1 = {compressDataVec_selectReqData_89, compressDataVec_selectReqData_88};
  wire [31:0]  compressDataVec_hi_hi_lo_hi_1 = {compressDataVec_selectReqData_91, compressDataVec_selectReqData_90};
  wire [63:0]  compressDataVec_hi_hi_lo_1 = {compressDataVec_hi_hi_lo_hi_1, compressDataVec_hi_hi_lo_lo_1};
  wire [31:0]  compressDataVec_hi_hi_hi_lo_1 = {compressDataVec_selectReqData_93, compressDataVec_selectReqData_92};
  wire [31:0]  compressDataVec_hi_hi_hi_hi_1 = {compressDataVec_selectReqData_95, compressDataVec_selectReqData_94};
  wire [63:0]  compressDataVec_hi_hi_hi_1 = {compressDataVec_hi_hi_hi_hi_1, compressDataVec_hi_hi_hi_lo_1};
  wire [127:0] compressDataVec_hi_hi_1 = {compressDataVec_hi_hi_hi_1, compressDataVec_hi_hi_lo_1};
  wire [255:0] compressDataVec_hi_1 = {compressDataVec_hi_hi_1, compressDataVec_hi_lo_1};
  wire [511:0] compressDataVec_1 = {compressDataVec_hi_1, compressDataVec_lo_1};
  wire [31:0]  compressDataVec_selectReqData_96 =
    (compressDataVec_hitReq_0_96 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_96 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_96 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_96 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_96 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_96 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_96 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_96 ? source2Pipe[255:224] : 32'h0);
  wire         compressDataVec_useTail_48;
  assign compressDataVec_useTail_48 = |tailCount;
  wire [31:0]  compressDataVec_selectReqData_97 =
    (compressDataVec_hitReq_0_97 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_97 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_97 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_97 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_97 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_97 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_97 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_97 ? source2Pipe[255:224] : 32'h0);
  wire         compressDataVec_useTail_49;
  assign compressDataVec_useTail_49 = |(tailCount[4:1]);
  wire [31:0]  compressDataVec_selectReqData_98 =
    (compressDataVec_hitReq_0_98 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_98 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_98 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_98 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_98 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_98 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_98 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_98 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_99 =
    (compressDataVec_hitReq_0_99 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_99 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_99 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_99 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_99 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_99 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_99 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_99 ? source2Pipe[255:224] : 32'h0);
  wire         compressDataVec_useTail_51;
  assign compressDataVec_useTail_51 = |(tailCount[4:2]);
  wire [31:0]  compressDataVec_selectReqData_100 =
    (compressDataVec_hitReq_0_100 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_100 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_100 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_100 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_100 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_100 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_100 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_100 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_101 =
    (compressDataVec_hitReq_0_101 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_101 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_101 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_101 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_101 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_101 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_101 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_101 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_102 =
    (compressDataVec_hitReq_0_102 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_102 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_102 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_102 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_102 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_102 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_102 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_102 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_103 =
    (compressDataVec_hitReq_0_103 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_103 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_103 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_103 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_103 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_103 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_103 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_103 ? source2Pipe[255:224] : 32'h0);
  wire         compressDataVec_useTail_55;
  assign compressDataVec_useTail_55 = |(tailCount[4:3]);
  wire [31:0]  compressDataVec_selectReqData_104 =
    (compressDataVec_hitReq_0_104 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_104 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_104 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_104 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_104 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_104 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_104 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_104 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_105 =
    (compressDataVec_hitReq_0_105 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_105 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_105 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_105 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_105 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_105 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_105 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_105 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_106 =
    (compressDataVec_hitReq_0_106 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_106 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_106 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_106 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_106 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_106 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_106 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_106 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_107 =
    (compressDataVec_hitReq_0_107 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_107 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_107 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_107 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_107 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_107 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_107 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_107 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_108 =
    (compressDataVec_hitReq_0_108 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_108 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_108 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_108 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_108 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_108 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_108 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_108 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_109 =
    (compressDataVec_hitReq_0_109 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_109 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_109 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_109 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_109 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_109 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_109 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_109 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_110 =
    (compressDataVec_hitReq_0_110 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_110 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_110 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_110 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_110 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_110 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_110 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_110 ? source2Pipe[255:224] : 32'h0);
  wire [31:0]  compressDataVec_selectReqData_111 =
    (compressDataVec_hitReq_0_111 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_111 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_111 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_111 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_111 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_111 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_111 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_111 ? source2Pipe[255:224] : 32'h0);
  wire [63:0]  compressDataVec_lo_lo_lo_2 = {compressDataVec_useTail_49 ? compressDataReg[63:32] : compressDataVec_selectReqData_97, compressDataVec_useTail_48 ? compressDataReg[31:0] : compressDataVec_selectReqData_96};
  wire [63:0]  compressDataVec_lo_lo_hi_2 = {compressDataVec_useTail_51 ? compressDataReg[127:96] : compressDataVec_selectReqData_99, compressDataVec_useTail_50 ? compressDataReg[95:64] : compressDataVec_selectReqData_98};
  wire [127:0] compressDataVec_lo_lo_2 = {compressDataVec_lo_lo_hi_2, compressDataVec_lo_lo_lo_2};
  wire [63:0]  compressDataVec_lo_hi_lo_2 = {compressDataVec_useTail_53 ? compressDataReg[191:160] : compressDataVec_selectReqData_101, compressDataVec_useTail_52 ? compressDataReg[159:128] : compressDataVec_selectReqData_100};
  wire [63:0]  compressDataVec_lo_hi_hi_2 = {compressDataVec_useTail_55 ? compressDataReg[255:224] : compressDataVec_selectReqData_103, compressDataVec_useTail_54 ? compressDataReg[223:192] : compressDataVec_selectReqData_102};
  wire [127:0] compressDataVec_lo_hi_2 = {compressDataVec_lo_hi_hi_2, compressDataVec_lo_hi_lo_2};
  wire [255:0] compressDataVec_lo_2 = {compressDataVec_lo_hi_2, compressDataVec_lo_lo_2};
  wire [63:0]  compressDataVec_hi_lo_lo_2 = {compressDataVec_selectReqData_105, compressDataVec_selectReqData_104};
  wire [63:0]  compressDataVec_hi_lo_hi_2 = {compressDataVec_selectReqData_107, compressDataVec_selectReqData_106};
  wire [127:0] compressDataVec_hi_lo_2 = {compressDataVec_hi_lo_hi_2, compressDataVec_hi_lo_lo_2};
  wire [63:0]  compressDataVec_hi_hi_lo_2 = {compressDataVec_selectReqData_109, compressDataVec_selectReqData_108};
  wire [63:0]  compressDataVec_hi_hi_hi_2 = {compressDataVec_selectReqData_111, compressDataVec_selectReqData_110};
  wire [127:0] compressDataVec_hi_hi_2 = {compressDataVec_hi_hi_hi_2, compressDataVec_hi_hi_lo_2};
  wire [255:0] compressDataVec_hi_2 = {compressDataVec_hi_hi_2, compressDataVec_hi_lo_2};
  wire [511:0] compressDataVec_2 = {compressDataVec_hi_2, compressDataVec_lo_2};
  wire [511:0] compressResult = (eew1H[0] ? compressDataVec_0 : 512'h0) | (eew1H[1] ? compressDataVec_1 : 512'h0) | (eew1H[2] ? compressDataVec_2 : 512'h0);
  wire         lastCompressEnq = stage2Valid & lastCompressPipe;
  wire [255:0] splitCompressResult_0 = compressResult[255:0];
  wire [255:0] splitCompressResult_1 = compressResult[511:256];
  wire         compressTailMask_elementValid;
  assign compressTailMask_elementValid = |tailCountForMask;
  wire         compressTailMask_elementValid_1;
  assign compressTailMask_elementValid_1 = |(tailCountForMask[4:1]);
  wire         _GEN_523 = tailCountForMask > 5'h2;
  wire         compressTailMask_elementValid_2;
  assign compressTailMask_elementValid_2 = _GEN_523;
  wire         compressTailMask_elementValid_34;
  assign compressTailMask_elementValid_34 = _GEN_523;
  wire         compressTailMask_elementValid_50;
  assign compressTailMask_elementValid_50 = _GEN_523;
  wire         compressTailMask_elementValid_3;
  assign compressTailMask_elementValid_3 = |(tailCountForMask[4:2]);
  wire         _GEN_524 = tailCountForMask > 5'h4;
  wire         compressTailMask_elementValid_4;
  assign compressTailMask_elementValid_4 = _GEN_524;
  wire         compressTailMask_elementValid_36;
  assign compressTailMask_elementValid_36 = _GEN_524;
  wire         compressTailMask_elementValid_52;
  assign compressTailMask_elementValid_52 = _GEN_524;
  wire         _GEN_525 = tailCountForMask > 5'h5;
  wire         compressTailMask_elementValid_5;
  assign compressTailMask_elementValid_5 = _GEN_525;
  wire         compressTailMask_elementValid_37;
  assign compressTailMask_elementValid_37 = _GEN_525;
  wire         compressTailMask_elementValid_53;
  assign compressTailMask_elementValid_53 = _GEN_525;
  wire         _GEN_526 = tailCountForMask > 5'h6;
  wire         compressTailMask_elementValid_6;
  assign compressTailMask_elementValid_6 = _GEN_526;
  wire         compressTailMask_elementValid_38;
  assign compressTailMask_elementValid_38 = _GEN_526;
  wire         compressTailMask_elementValid_54;
  assign compressTailMask_elementValid_54 = _GEN_526;
  wire         compressTailMask_elementValid_7;
  assign compressTailMask_elementValid_7 = |(tailCountForMask[4:3]);
  wire         _GEN_527 = tailCountForMask > 5'h8;
  wire         compressTailMask_elementValid_8;
  assign compressTailMask_elementValid_8 = _GEN_527;
  wire         compressTailMask_elementValid_40;
  assign compressTailMask_elementValid_40 = _GEN_527;
  wire         _GEN_528 = tailCountForMask > 5'h9;
  wire         compressTailMask_elementValid_9;
  assign compressTailMask_elementValid_9 = _GEN_528;
  wire         compressTailMask_elementValid_41;
  assign compressTailMask_elementValid_41 = _GEN_528;
  wire         _GEN_529 = tailCountForMask > 5'hA;
  wire         compressTailMask_elementValid_10;
  assign compressTailMask_elementValid_10 = _GEN_529;
  wire         compressTailMask_elementValid_42;
  assign compressTailMask_elementValid_42 = _GEN_529;
  wire         _GEN_530 = tailCountForMask > 5'hB;
  wire         compressTailMask_elementValid_11;
  assign compressTailMask_elementValid_11 = _GEN_530;
  wire         compressTailMask_elementValid_43;
  assign compressTailMask_elementValid_43 = _GEN_530;
  wire         _GEN_531 = tailCountForMask > 5'hC;
  wire         compressTailMask_elementValid_12;
  assign compressTailMask_elementValid_12 = _GEN_531;
  wire         compressTailMask_elementValid_44;
  assign compressTailMask_elementValid_44 = _GEN_531;
  wire         _GEN_532 = tailCountForMask > 5'hD;
  wire         compressTailMask_elementValid_13;
  assign compressTailMask_elementValid_13 = _GEN_532;
  wire         compressTailMask_elementValid_45;
  assign compressTailMask_elementValid_45 = _GEN_532;
  wire         _GEN_533 = tailCountForMask > 5'hE;
  wire         compressTailMask_elementValid_14;
  assign compressTailMask_elementValid_14 = _GEN_533;
  wire         compressTailMask_elementValid_46;
  assign compressTailMask_elementValid_46 = _GEN_533;
  wire         compressTailMask_elementValid_15 = tailCountForMask[4];
  wire         compressTailMask_elementValid_47 = tailCountForMask[4];
  wire         compressTailMask_elementValid_16 = tailCountForMask > 5'h10;
  wire         compressTailMask_elementValid_17 = tailCountForMask > 5'h11;
  wire         compressTailMask_elementValid_18 = tailCountForMask > 5'h12;
  wire         compressTailMask_elementValid_19 = tailCountForMask > 5'h13;
  wire         compressTailMask_elementValid_20 = tailCountForMask > 5'h14;
  wire         compressTailMask_elementValid_21 = tailCountForMask > 5'h15;
  wire         compressTailMask_elementValid_22 = tailCountForMask > 5'h16;
  wire         compressTailMask_elementValid_23 = tailCountForMask > 5'h17;
  wire         compressTailMask_elementValid_24 = tailCountForMask > 5'h18;
  wire         compressTailMask_elementValid_25 = tailCountForMask > 5'h19;
  wire         compressTailMask_elementValid_26 = tailCountForMask > 5'h1A;
  wire         compressTailMask_elementValid_27 = tailCountForMask > 5'h1B;
  wire         compressTailMask_elementValid_28 = tailCountForMask > 5'h1C;
  wire         compressTailMask_elementValid_29 = tailCountForMask > 5'h1D;
  wire         compressTailMask_elementValid_30 = &tailCountForMask;
  wire [1:0]   compressTailMask_lo_lo_lo_lo = {compressTailMask_elementValid_1, compressTailMask_elementValid};
  wire [1:0]   compressTailMask_lo_lo_lo_hi = {compressTailMask_elementValid_3, compressTailMask_elementValid_2};
  wire [3:0]   compressTailMask_lo_lo_lo = {compressTailMask_lo_lo_lo_hi, compressTailMask_lo_lo_lo_lo};
  wire [1:0]   compressTailMask_lo_lo_hi_lo = {compressTailMask_elementValid_5, compressTailMask_elementValid_4};
  wire [1:0]   compressTailMask_lo_lo_hi_hi = {compressTailMask_elementValid_7, compressTailMask_elementValid_6};
  wire [3:0]   compressTailMask_lo_lo_hi = {compressTailMask_lo_lo_hi_hi, compressTailMask_lo_lo_hi_lo};
  wire [7:0]   compressTailMask_lo_lo = {compressTailMask_lo_lo_hi, compressTailMask_lo_lo_lo};
  wire [1:0]   compressTailMask_lo_hi_lo_lo = {compressTailMask_elementValid_9, compressTailMask_elementValid_8};
  wire [1:0]   compressTailMask_lo_hi_lo_hi = {compressTailMask_elementValid_11, compressTailMask_elementValid_10};
  wire [3:0]   compressTailMask_lo_hi_lo = {compressTailMask_lo_hi_lo_hi, compressTailMask_lo_hi_lo_lo};
  wire [1:0]   compressTailMask_lo_hi_hi_lo = {compressTailMask_elementValid_13, compressTailMask_elementValid_12};
  wire [1:0]   compressTailMask_lo_hi_hi_hi = {compressTailMask_elementValid_15, compressTailMask_elementValid_14};
  wire [3:0]   compressTailMask_lo_hi_hi = {compressTailMask_lo_hi_hi_hi, compressTailMask_lo_hi_hi_lo};
  wire [7:0]   compressTailMask_lo_hi = {compressTailMask_lo_hi_hi, compressTailMask_lo_hi_lo};
  wire [15:0]  compressTailMask_lo = {compressTailMask_lo_hi, compressTailMask_lo_lo};
  wire [1:0]   compressTailMask_hi_lo_lo_lo = {compressTailMask_elementValid_17, compressTailMask_elementValid_16};
  wire [1:0]   compressTailMask_hi_lo_lo_hi = {compressTailMask_elementValid_19, compressTailMask_elementValid_18};
  wire [3:0]   compressTailMask_hi_lo_lo = {compressTailMask_hi_lo_lo_hi, compressTailMask_hi_lo_lo_lo};
  wire [1:0]   compressTailMask_hi_lo_hi_lo = {compressTailMask_elementValid_21, compressTailMask_elementValid_20};
  wire [1:0]   compressTailMask_hi_lo_hi_hi = {compressTailMask_elementValid_23, compressTailMask_elementValid_22};
  wire [3:0]   compressTailMask_hi_lo_hi = {compressTailMask_hi_lo_hi_hi, compressTailMask_hi_lo_hi_lo};
  wire [7:0]   compressTailMask_hi_lo = {compressTailMask_hi_lo_hi, compressTailMask_hi_lo_lo};
  wire [1:0]   compressTailMask_hi_hi_lo_lo = {compressTailMask_elementValid_25, compressTailMask_elementValid_24};
  wire [1:0]   compressTailMask_hi_hi_lo_hi = {compressTailMask_elementValid_27, compressTailMask_elementValid_26};
  wire [3:0]   compressTailMask_hi_hi_lo = {compressTailMask_hi_hi_lo_hi, compressTailMask_hi_hi_lo_lo};
  wire [1:0]   compressTailMask_hi_hi_hi_lo = {compressTailMask_elementValid_29, compressTailMask_elementValid_28};
  wire [1:0]   compressTailMask_hi_hi_hi_hi = {1'h0, compressTailMask_elementValid_30};
  wire [3:0]   compressTailMask_hi_hi_hi = {compressTailMask_hi_hi_hi_hi, compressTailMask_hi_hi_hi_lo};
  wire [7:0]   compressTailMask_hi_hi = {compressTailMask_hi_hi_hi, compressTailMask_hi_hi_lo};
  wire [15:0]  compressTailMask_hi = {compressTailMask_hi_hi, compressTailMask_hi_lo};
  wire         compressTailMask_elementValid_32;
  assign compressTailMask_elementValid_32 = |tailCountForMask;
  wire [1:0]   compressTailMask_elementMask = {2{compressTailMask_elementValid_32}};
  wire         compressTailMask_elementValid_33;
  assign compressTailMask_elementValid_33 = |(tailCountForMask[4:1]);
  wire [1:0]   compressTailMask_elementMask_1 = {2{compressTailMask_elementValid_33}};
  wire [1:0]   compressTailMask_elementMask_2 = {2{compressTailMask_elementValid_34}};
  wire         compressTailMask_elementValid_35;
  assign compressTailMask_elementValid_35 = |(tailCountForMask[4:2]);
  wire [1:0]   compressTailMask_elementMask_3 = {2{compressTailMask_elementValid_35}};
  wire [1:0]   compressTailMask_elementMask_4 = {2{compressTailMask_elementValid_36}};
  wire [1:0]   compressTailMask_elementMask_5 = {2{compressTailMask_elementValid_37}};
  wire [1:0]   compressTailMask_elementMask_6 = {2{compressTailMask_elementValid_38}};
  wire         compressTailMask_elementValid_39;
  assign compressTailMask_elementValid_39 = |(tailCountForMask[4:3]);
  wire [1:0]   compressTailMask_elementMask_7 = {2{compressTailMask_elementValid_39}};
  wire [1:0]   compressTailMask_elementMask_8 = {2{compressTailMask_elementValid_40}};
  wire [1:0]   compressTailMask_elementMask_9 = {2{compressTailMask_elementValid_41}};
  wire [1:0]   compressTailMask_elementMask_10 = {2{compressTailMask_elementValid_42}};
  wire [1:0]   compressTailMask_elementMask_11 = {2{compressTailMask_elementValid_43}};
  wire [1:0]   compressTailMask_elementMask_12 = {2{compressTailMask_elementValid_44}};
  wire [1:0]   compressTailMask_elementMask_13 = {2{compressTailMask_elementValid_45}};
  wire [1:0]   compressTailMask_elementMask_14 = {2{compressTailMask_elementValid_46}};
  wire [1:0]   compressTailMask_elementMask_15 = {2{compressTailMask_elementValid_47}};
  wire [3:0]   compressTailMask_lo_lo_lo_1 = {compressTailMask_elementMask_1, compressTailMask_elementMask};
  wire [3:0]   compressTailMask_lo_lo_hi_1 = {compressTailMask_elementMask_3, compressTailMask_elementMask_2};
  wire [7:0]   compressTailMask_lo_lo_1 = {compressTailMask_lo_lo_hi_1, compressTailMask_lo_lo_lo_1};
  wire [3:0]   compressTailMask_lo_hi_lo_1 = {compressTailMask_elementMask_5, compressTailMask_elementMask_4};
  wire [3:0]   compressTailMask_lo_hi_hi_1 = {compressTailMask_elementMask_7, compressTailMask_elementMask_6};
  wire [7:0]   compressTailMask_lo_hi_1 = {compressTailMask_lo_hi_hi_1, compressTailMask_lo_hi_lo_1};
  wire [15:0]  compressTailMask_lo_1 = {compressTailMask_lo_hi_1, compressTailMask_lo_lo_1};
  wire [3:0]   compressTailMask_hi_lo_lo_1 = {compressTailMask_elementMask_9, compressTailMask_elementMask_8};
  wire [3:0]   compressTailMask_hi_lo_hi_1 = {compressTailMask_elementMask_11, compressTailMask_elementMask_10};
  wire [7:0]   compressTailMask_hi_lo_1 = {compressTailMask_hi_lo_hi_1, compressTailMask_hi_lo_lo_1};
  wire [3:0]   compressTailMask_hi_hi_lo_1 = {compressTailMask_elementMask_13, compressTailMask_elementMask_12};
  wire [3:0]   compressTailMask_hi_hi_hi_1 = {compressTailMask_elementMask_15, compressTailMask_elementMask_14};
  wire [7:0]   compressTailMask_hi_hi_1 = {compressTailMask_hi_hi_hi_1, compressTailMask_hi_hi_lo_1};
  wire [15:0]  compressTailMask_hi_1 = {compressTailMask_hi_hi_1, compressTailMask_hi_lo_1};
  wire         compressTailMask_elementValid_48;
  assign compressTailMask_elementValid_48 = |tailCountForMask;
  wire [3:0]   compressTailMask_elementMask_16 = {4{compressTailMask_elementValid_48}};
  wire         compressTailMask_elementValid_49;
  assign compressTailMask_elementValid_49 = |(tailCountForMask[4:1]);
  wire [3:0]   compressTailMask_elementMask_17 = {4{compressTailMask_elementValid_49}};
  wire [3:0]   compressTailMask_elementMask_18 = {4{compressTailMask_elementValid_50}};
  wire         compressTailMask_elementValid_51;
  assign compressTailMask_elementValid_51 = |(tailCountForMask[4:2]);
  wire [3:0]   compressTailMask_elementMask_19 = {4{compressTailMask_elementValid_51}};
  wire [3:0]   compressTailMask_elementMask_20 = {4{compressTailMask_elementValid_52}};
  wire [3:0]   compressTailMask_elementMask_21 = {4{compressTailMask_elementValid_53}};
  wire [3:0]   compressTailMask_elementMask_22 = {4{compressTailMask_elementValid_54}};
  wire         compressTailMask_elementValid_55;
  assign compressTailMask_elementValid_55 = |(tailCountForMask[4:3]);
  wire [3:0]   compressTailMask_elementMask_23 = {4{compressTailMask_elementValid_55}};
  wire [7:0]   compressTailMask_lo_lo_2 = {compressTailMask_elementMask_17, compressTailMask_elementMask_16};
  wire [7:0]   compressTailMask_lo_hi_2 = {compressTailMask_elementMask_19, compressTailMask_elementMask_18};
  wire [15:0]  compressTailMask_lo_2 = {compressTailMask_lo_hi_2, compressTailMask_lo_lo_2};
  wire [7:0]   compressTailMask_hi_lo_2 = {compressTailMask_elementMask_21, compressTailMask_elementMask_20};
  wire [7:0]   compressTailMask_hi_hi_2 = {compressTailMask_elementMask_23, compressTailMask_elementMask_22};
  wire [15:0]  compressTailMask_hi_2 = {compressTailMask_hi_hi_2, compressTailMask_hi_lo_2};
  wire [31:0]  compressTailMask = (eew1H[0] ? {compressTailMask_hi, compressTailMask_lo} : 32'h0) | (eew1H[1] ? {compressTailMask_hi_1, compressTailMask_lo_1} : 32'h0) | (eew1H[2] ? {compressTailMask_hi_2, compressTailMask_lo_2} : 32'h0);
  wire [31:0]  compressMask = compressTailValid ? compressTailMask : 32'hFFFFFFFF;
  reg  [7:0]   validInputPipe;
  reg  [31:0]  readFromScalarPipe;
  wire [3:0]   mvMask = {2'h0, {1'h0, eew1H[0]} | {2{eew1H[1]}}} | {4{eew1H[2]}};
  wire [7:0]   ffoMask_lo_lo = {{4{validInputPipe[1]}}, {4{validInputPipe[0]}}};
  wire [7:0]   ffoMask_lo_hi = {{4{validInputPipe[3]}}, {4{validInputPipe[2]}}};
  wire [15:0]  ffoMask_lo = {ffoMask_lo_hi, ffoMask_lo_lo};
  wire [7:0]   ffoMask_hi_lo = {{4{validInputPipe[5]}}, {4{validInputPipe[4]}}};
  wire [7:0]   ffoMask_hi_hi = {{4{validInputPipe[7]}}, {4{validInputPipe[6]}}};
  wire [15:0]  ffoMask_hi = {ffoMask_hi_hi, ffoMask_hi_lo};
  wire [31:0]  ffoMask = {ffoMask_hi, ffoMask_lo};
  wire [7:0]   outWire_ffoOutput;
  wire [63:0]  ffoData_lo_lo = {outWire_ffoOutput[1] ? in_1_bits_pipeData[63:32] : in_1_bits_source2[63:32], outWire_ffoOutput[0] ? in_1_bits_pipeData[31:0] : in_1_bits_source2[31:0]};
  wire [63:0]  ffoData_lo_hi = {outWire_ffoOutput[3] ? in_1_bits_pipeData[127:96] : in_1_bits_source2[127:96], outWire_ffoOutput[2] ? in_1_bits_pipeData[95:64] : in_1_bits_source2[95:64]};
  wire [127:0] ffoData_lo = {ffoData_lo_hi, ffoData_lo_lo};
  wire [63:0]  ffoData_hi_lo = {outWire_ffoOutput[5] ? in_1_bits_pipeData[191:160] : in_1_bits_source2[191:160], outWire_ffoOutput[4] ? in_1_bits_pipeData[159:128] : in_1_bits_source2[159:128]};
  wire [63:0]  ffoData_hi_hi = {outWire_ffoOutput[7] ? in_1_bits_pipeData[255:224] : in_1_bits_source2[255:224], outWire_ffoOutput[6] ? in_1_bits_pipeData[223:192] : in_1_bits_source2[223:192]};
  wire [127:0] ffoData_hi = {ffoData_hi_hi, ffoData_hi_lo};
  wire [255:0] ffoData = {ffoData_hi, ffoData_lo};
  wire [255:0] _GEN_534 = (compress ? compressResult[255:0] : 256'h0) | (viota ? viotaResult : 256'h0);
  wire [255:0] outWire_data = {_GEN_534[255:32], _GEN_534[31:0] | (mv ? readFromScalarPipe : 32'h0)} | (ffoType ? ffoData : 256'h0);
  wire [31:0]  _outWire_mask_T_4 = (compress ? compressMask : 32'h0) | (viota ? viotaMask : 32'h0);
  wire [31:0]  outWire_mask = {_outWire_mask_T_4[31:4], _outWire_mask_T_4[3:0] | (mv ? mvMask : 4'h0)} | (ffoType ? ffoMask : 32'h0);
  wire         outWire_compressValid = (compressTailValid | compressDeqValidPipe & stage2Valid) & ~writeRD;
  wire [5:0]   outWire_groupCounter = compress ? compressWriteGroupCount : groupCounterPipe;
  wire [6:0]   _completedLeftOr_T_2 = in_1_bits_ffoInput[6:0] | {in_1_bits_ffoInput[5:0], 1'h0};
  wire [6:0]   _GEN_535 = {_completedLeftOr_T_2[4:0], 2'h0};
  wire [6:0]   _firstLane_T_5 = _completedLeftOr_T_2 | _GEN_535;
  wire [7:0]   firstLane = {~(_firstLane_T_5 | {_firstLane_T_5[2:0], 4'h0}), 1'h1} & in_1_bits_ffoInput;
  wire [3:0]   firstLaneIndex_hi = firstLane[7:4];
  wire [3:0]   firstLaneIndex_lo = firstLane[3:0];
  wire [3:0]   _firstLaneIndex_T_1 = firstLaneIndex_hi | firstLaneIndex_lo;
  wire [1:0]   firstLaneIndex_hi_1 = _firstLaneIndex_T_1[3:2];
  wire [1:0]   firstLaneIndex_lo_1 = _firstLaneIndex_T_1[1:0];
  wire [2:0]   firstLaneIndex = {|firstLaneIndex_hi, |firstLaneIndex_hi_1, firstLaneIndex_hi_1[1] | firstLaneIndex_lo_1[1]};
  wire [31:0]  source1SigExtend = (eew1H[0] ? {{24{in_1_bits_source1[7]}}, in_1_bits_source1[7:0]} : 32'h0) | (eew1H[1] ? {{16{in_1_bits_source1[15]}}, in_1_bits_source1[15:0]} : 32'h0) | (eew1H[2] ? in_1_bits_source1 : 32'h0);
  wire [6:0]   _completedLeftOr_T_5 = _completedLeftOr_T_2 | _GEN_535;
  wire [7:0]   completedLeftOr = {_completedLeftOr_T_5 | {_completedLeftOr_T_5[2:0], 4'h0}, 1'h0};
  reg  [7:0]   ffoOutPipe;
  assign outWire_ffoOutput = ffoOutPipe;
  reg  [255:0] view__out_REG_data;
  reg  [31:0]  view__out_REG_mask;
  reg  [5:0]   view__out_REG_groupCounter;
  reg  [7:0]   view__out_REG_ffoOutput;
  reg          view__out_REG_compressValid;
  always @(posedge clock) begin
    if (reset) begin
      in_1_valid <= 1'h0;
      in_1_bits_maskType <= 1'h0;
      in_1_bits_eew <= 2'h0;
      in_1_bits_uop <= 3'h0;
      in_1_bits_readFromScalar <= 32'h0;
      in_1_bits_source1 <= 32'h0;
      in_1_bits_mask <= 32'h0;
      in_1_bits_source2 <= 256'h0;
      in_1_bits_pipeData <= 256'h0;
      in_1_bits_groupCounter <= 6'h0;
      in_1_bits_ffoInput <= 8'h0;
      in_1_bits_validInput <= 8'h0;
      in_1_bits_lastCompress <= 1'h0;
      compressInit <= 10'h0;
      ffoIndex <= 32'h0;
      ffoValid <= 1'h0;
      compressVecPipe_0 <= 10'h0;
      compressVecPipe_1 <= 10'h0;
      compressVecPipe_2 <= 10'h0;
      compressVecPipe_3 <= 10'h0;
      compressVecPipe_4 <= 10'h0;
      compressVecPipe_5 <= 10'h0;
      compressVecPipe_6 <= 10'h0;
      compressVecPipe_7 <= 10'h0;
      compressVecPipe_8 <= 10'h0;
      compressVecPipe_9 <= 10'h0;
      compressVecPipe_10 <= 10'h0;
      compressVecPipe_11 <= 10'h0;
      compressVecPipe_12 <= 10'h0;
      compressVecPipe_13 <= 10'h0;
      compressVecPipe_14 <= 10'h0;
      compressVecPipe_15 <= 10'h0;
      compressVecPipe_16 <= 10'h0;
      compressVecPipe_17 <= 10'h0;
      compressVecPipe_18 <= 10'h0;
      compressVecPipe_19 <= 10'h0;
      compressVecPipe_20 <= 10'h0;
      compressVecPipe_21 <= 10'h0;
      compressVecPipe_22 <= 10'h0;
      compressVecPipe_23 <= 10'h0;
      compressVecPipe_24 <= 10'h0;
      compressVecPipe_25 <= 10'h0;
      compressVecPipe_26 <= 10'h0;
      compressVecPipe_27 <= 10'h0;
      compressVecPipe_28 <= 10'h0;
      compressVecPipe_29 <= 10'h0;
      compressVecPipe_30 <= 10'h0;
      compressVecPipe_31 <= 10'h0;
      compressMaskVecPipe_0 <= 1'h0;
      compressMaskVecPipe_1 <= 1'h0;
      compressMaskVecPipe_2 <= 1'h0;
      compressMaskVecPipe_3 <= 1'h0;
      compressMaskVecPipe_4 <= 1'h0;
      compressMaskVecPipe_5 <= 1'h0;
      compressMaskVecPipe_6 <= 1'h0;
      compressMaskVecPipe_7 <= 1'h0;
      compressMaskVecPipe_8 <= 1'h0;
      compressMaskVecPipe_9 <= 1'h0;
      compressMaskVecPipe_10 <= 1'h0;
      compressMaskVecPipe_11 <= 1'h0;
      compressMaskVecPipe_12 <= 1'h0;
      compressMaskVecPipe_13 <= 1'h0;
      compressMaskVecPipe_14 <= 1'h0;
      compressMaskVecPipe_15 <= 1'h0;
      compressMaskVecPipe_16 <= 1'h0;
      compressMaskVecPipe_17 <= 1'h0;
      compressMaskVecPipe_18 <= 1'h0;
      compressMaskVecPipe_19 <= 1'h0;
      compressMaskVecPipe_20 <= 1'h0;
      compressMaskVecPipe_21 <= 1'h0;
      compressMaskVecPipe_22 <= 1'h0;
      compressMaskVecPipe_23 <= 1'h0;
      compressMaskVecPipe_24 <= 1'h0;
      compressMaskVecPipe_25 <= 1'h0;
      compressMaskVecPipe_26 <= 1'h0;
      compressMaskVecPipe_27 <= 1'h0;
      compressMaskVecPipe_28 <= 1'h0;
      compressMaskVecPipe_29 <= 1'h0;
      compressMaskVecPipe_30 <= 1'h0;
      compressMaskVecPipe_31 <= 1'h0;
      maskPipe <= 32'h0;
      source2Pipe <= 256'h0;
      lastCompressPipe <= 1'h0;
      stage2Valid <= 1'h0;
      newInstructionPipe <= 1'h0;
      compressInitPipe <= 10'h0;
      compressDeqValidPipe <= 1'h0;
      groupCounterPipe <= 6'h0;
      compressDataReg <= 256'h0;
      compressTailValid <= 1'h0;
      compressWriteGroupCount <= 6'h0;
      validInputPipe <= 8'h0;
      readFromScalarPipe <= 32'h0;
      ffoOutPipe <= 8'h0;
      view__out_REG_data <= 256'h0;
      view__out_REG_mask <= 32'h0;
      view__out_REG_groupCounter <= 6'h0;
      view__out_REG_ffoOutput <= 8'h0;
      view__out_REG_compressValid <= 1'h0;
    end
    else begin
      automatic logic _GEN_536;
      automatic logic _GEN_537;
      _GEN_536 = newInstruction & ffoInstruction;
      _GEN_537 = in_1_valid & (|in_1_bits_ffoInput) & ffoType;
      in_1_valid <= in_valid;
      in_1_bits_maskType <= in_bits_maskType;
      in_1_bits_eew <= in_bits_eew;
      in_1_bits_uop <= in_bits_uop;
      in_1_bits_readFromScalar <= in_bits_readFromScalar;
      in_1_bits_source1 <= in_bits_source1;
      in_1_bits_mask <= in_bits_mask;
      in_1_bits_source2 <= in_bits_source2;
      in_1_bits_pipeData <= in_bits_pipeData;
      in_1_bits_groupCounter <= in_bits_groupCounter;
      in_1_bits_ffoInput <= in_bits_ffoInput;
      in_1_bits_validInput <= in_bits_validInput;
      in_1_bits_lastCompress <= in_bits_lastCompress;
      if (in_1_valid) begin
        compressInit <= viota ? compressCount : {5'h0, compressCountSelect};
        compressVecPipe_0 <= compressVec_0;
        compressVecPipe_1 <= compressVec_1;
        compressVecPipe_2 <= compressVec_2;
        compressVecPipe_3 <= compressVec_3;
        compressVecPipe_4 <= compressVec_4;
        compressVecPipe_5 <= compressVec_5;
        compressVecPipe_6 <= compressVec_6;
        compressVecPipe_7 <= compressVec_7;
        compressVecPipe_8 <= compressVec_8;
        compressVecPipe_9 <= compressVec_9;
        compressVecPipe_10 <= compressVec_10;
        compressVecPipe_11 <= compressVec_11;
        compressVecPipe_12 <= compressVec_12;
        compressVecPipe_13 <= compressVec_13;
        compressVecPipe_14 <= compressVec_14;
        compressVecPipe_15 <= compressVec_15;
        compressVecPipe_16 <= compressVec_16;
        compressVecPipe_17 <= compressVec_17;
        compressVecPipe_18 <= compressVec_18;
        compressVecPipe_19 <= compressVec_19;
        compressVecPipe_20 <= compressVec_20;
        compressVecPipe_21 <= compressVec_21;
        compressVecPipe_22 <= compressVec_22;
        compressVecPipe_23 <= compressVec_23;
        compressVecPipe_24 <= compressVec_24;
        compressVecPipe_25 <= compressVec_25;
        compressVecPipe_26 <= compressVec_26;
        compressVecPipe_27 <= compressVec_27;
        compressVecPipe_28 <= compressVec_28;
        compressVecPipe_29 <= compressVec_29;
        compressVecPipe_30 <= compressVec_30;
        compressVecPipe_31 <= compressVec_31;
        compressMaskVecPipe_0 <= compressMaskVec_0;
        compressMaskVecPipe_1 <= compressMaskVec_1;
        compressMaskVecPipe_2 <= compressMaskVec_2;
        compressMaskVecPipe_3 <= compressMaskVec_3;
        compressMaskVecPipe_4 <= compressMaskVec_4;
        compressMaskVecPipe_5 <= compressMaskVec_5;
        compressMaskVecPipe_6 <= compressMaskVec_6;
        compressMaskVecPipe_7 <= compressMaskVec_7;
        compressMaskVecPipe_8 <= compressMaskVec_8;
        compressMaskVecPipe_9 <= compressMaskVec_9;
        compressMaskVecPipe_10 <= compressMaskVec_10;
        compressMaskVecPipe_11 <= compressMaskVec_11;
        compressMaskVecPipe_12 <= compressMaskVec_12;
        compressMaskVecPipe_13 <= compressMaskVec_13;
        compressMaskVecPipe_14 <= compressMaskVec_14;
        compressMaskVecPipe_15 <= compressMaskVec_15;
        compressMaskVecPipe_16 <= compressMaskVec_16;
        compressMaskVecPipe_17 <= compressMaskVec_17;
        compressMaskVecPipe_18 <= compressMaskVec_18;
        compressMaskVecPipe_19 <= compressMaskVec_19;
        compressMaskVecPipe_20 <= compressMaskVec_20;
        compressMaskVecPipe_21 <= compressMaskVec_21;
        compressMaskVecPipe_22 <= compressMaskVec_22;
        compressMaskVecPipe_23 <= compressMaskVec_23;
        compressMaskVecPipe_24 <= compressMaskVec_24;
        compressMaskVecPipe_25 <= compressMaskVec_25;
        compressMaskVecPipe_26 <= compressMaskVec_26;
        compressMaskVecPipe_27 <= compressMaskVec_27;
        compressMaskVecPipe_28 <= compressMaskVec_28;
        compressMaskVecPipe_29 <= compressMaskVec_29;
        compressMaskVecPipe_30 <= compressMaskVec_30;
        compressMaskVecPipe_31 <= compressMaskVec_31;
        maskPipe <= in_1_bits_mask;
        source2Pipe <= in_1_bits_source2;
        lastCompressPipe <= in_1_bits_lastCompress;
        compressInitPipe <= compressInit;
        compressDeqValidPipe <= compressDeqValid;
        groupCounterPipe <= in_1_bits_groupCounter;
        validInputPipe <= in_1_bits_validInput;
        readFromScalarPipe <= in_1_bits_readFromScalar;
        ffoOutPipe <= completedLeftOr | {8{ffoValid}};
      end
      else if (newInstruction)
        compressInit <= 10'h0;
      if (_GEN_537) begin
        if (ffoValid) begin
          if (_GEN_536)
            ffoIndex <= 32'hFFFFFFFF;
        end
        else
          ffoIndex <=
            (firstLane[0] ? {in_1_bits_source2[28:5], firstLaneIndex, in_1_bits_source2[4:0]} : 32'h0) | (firstLane[1] ? {in_1_bits_source2[60:37], firstLaneIndex, in_1_bits_source2[36:32]} : 32'h0)
            | (firstLane[2] ? {in_1_bits_source2[92:69], firstLaneIndex, in_1_bits_source2[68:64]} : 32'h0) | (firstLane[3] ? {in_1_bits_source2[124:101], firstLaneIndex, in_1_bits_source2[100:96]} : 32'h0)
            | (firstLane[4] ? {in_1_bits_source2[156:133], firstLaneIndex, in_1_bits_source2[132:128]} : 32'h0) | (firstLane[5] ? {in_1_bits_source2[188:165], firstLaneIndex, in_1_bits_source2[164:160]} : 32'h0)
            | (firstLane[6] ? {in_1_bits_source2[220:197], firstLaneIndex, in_1_bits_source2[196:192]} : 32'h0) | (firstLane[7] ? {in_1_bits_source2[252:229], firstLaneIndex, in_1_bits_source2[228:224]} : 32'h0);
      end
      else if (mvRd)
        ffoIndex <= source1SigExtend;
      else if (_GEN_536)
        ffoIndex <= 32'hFFFFFFFF;
      ffoValid <= _GEN_537 | ~_GEN_536 & ffoValid;
      stage2Valid <= in_1_valid;
      newInstructionPipe <= newInstruction;
      if (stage2Valid)
        compressDataReg <= compressDeqValidPipe ? splitCompressResult_1 : splitCompressResult_0;
      if (newInstructionPipe | lastCompressEnq | outWire_compressValid)
        compressTailValid <= lastCompressEnq & compress;
      if (newInstructionPipe | outWire_compressValid)
        compressWriteGroupCount <= newInstructionPipe ? 6'h0 : compressWriteGroupCount + 6'h1;
      view__out_REG_data <= outWire_data;
      view__out_REG_mask <= outWire_mask;
      view__out_REG_groupCounter <= outWire_groupCounter;
      view__out_REG_ffoOutput <= outWire_ffoOutput;
      view__out_REG_compressValid <= outWire_compressValid;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:61];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [5:0] i = 6'h0; i < 6'h3E; i += 6'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        in_1_valid = _RANDOM[6'h0][0];
        in_1_bits_maskType = _RANDOM[6'h0][1];
        in_1_bits_eew = _RANDOM[6'h0][3:2];
        in_1_bits_uop = _RANDOM[6'h0][6:4];
        in_1_bits_readFromScalar = {_RANDOM[6'h0][31:7], _RANDOM[6'h1][6:0]};
        in_1_bits_source1 = {_RANDOM[6'h1][31:7], _RANDOM[6'h2][6:0]};
        in_1_bits_mask = {_RANDOM[6'h2][31:7], _RANDOM[6'h3][6:0]};
        in_1_bits_source2 = {_RANDOM[6'h3][31:7], _RANDOM[6'h4], _RANDOM[6'h5], _RANDOM[6'h6], _RANDOM[6'h7], _RANDOM[6'h8], _RANDOM[6'h9], _RANDOM[6'hA], _RANDOM[6'hB][6:0]};
        in_1_bits_pipeData = {_RANDOM[6'hB][31:7], _RANDOM[6'hC], _RANDOM[6'hD], _RANDOM[6'hE], _RANDOM[6'hF], _RANDOM[6'h10], _RANDOM[6'h11], _RANDOM[6'h12], _RANDOM[6'h13][6:0]};
        in_1_bits_groupCounter = _RANDOM[6'h13][12:7];
        in_1_bits_ffoInput = _RANDOM[6'h13][20:13];
        in_1_bits_validInput = _RANDOM[6'h13][28:21];
        in_1_bits_lastCompress = _RANDOM[6'h13][29];
        compressInit = {_RANDOM[6'h13][31:30], _RANDOM[6'h14][7:0]};
        ffoIndex = {_RANDOM[6'h14][31:8], _RANDOM[6'h15][7:0]};
        ffoValid = _RANDOM[6'h15][8];
        compressVecPipe_0 = _RANDOM[6'h15][18:9];
        compressVecPipe_1 = _RANDOM[6'h15][28:19];
        compressVecPipe_2 = {_RANDOM[6'h15][31:29], _RANDOM[6'h16][6:0]};
        compressVecPipe_3 = _RANDOM[6'h16][16:7];
        compressVecPipe_4 = _RANDOM[6'h16][26:17];
        compressVecPipe_5 = {_RANDOM[6'h16][31:27], _RANDOM[6'h17][4:0]};
        compressVecPipe_6 = _RANDOM[6'h17][14:5];
        compressVecPipe_7 = _RANDOM[6'h17][24:15];
        compressVecPipe_8 = {_RANDOM[6'h17][31:25], _RANDOM[6'h18][2:0]};
        compressVecPipe_9 = _RANDOM[6'h18][12:3];
        compressVecPipe_10 = _RANDOM[6'h18][22:13];
        compressVecPipe_11 = {_RANDOM[6'h18][31:23], _RANDOM[6'h19][0]};
        compressVecPipe_12 = _RANDOM[6'h19][10:1];
        compressVecPipe_13 = _RANDOM[6'h19][20:11];
        compressVecPipe_14 = _RANDOM[6'h19][30:21];
        compressVecPipe_15 = {_RANDOM[6'h19][31], _RANDOM[6'h1A][8:0]};
        compressVecPipe_16 = _RANDOM[6'h1A][18:9];
        compressVecPipe_17 = _RANDOM[6'h1A][28:19];
        compressVecPipe_18 = {_RANDOM[6'h1A][31:29], _RANDOM[6'h1B][6:0]};
        compressVecPipe_19 = _RANDOM[6'h1B][16:7];
        compressVecPipe_20 = _RANDOM[6'h1B][26:17];
        compressVecPipe_21 = {_RANDOM[6'h1B][31:27], _RANDOM[6'h1C][4:0]};
        compressVecPipe_22 = _RANDOM[6'h1C][14:5];
        compressVecPipe_23 = _RANDOM[6'h1C][24:15];
        compressVecPipe_24 = {_RANDOM[6'h1C][31:25], _RANDOM[6'h1D][2:0]};
        compressVecPipe_25 = _RANDOM[6'h1D][12:3];
        compressVecPipe_26 = _RANDOM[6'h1D][22:13];
        compressVecPipe_27 = {_RANDOM[6'h1D][31:23], _RANDOM[6'h1E][0]};
        compressVecPipe_28 = _RANDOM[6'h1E][10:1];
        compressVecPipe_29 = _RANDOM[6'h1E][20:11];
        compressVecPipe_30 = _RANDOM[6'h1E][30:21];
        compressVecPipe_31 = {_RANDOM[6'h1E][31], _RANDOM[6'h1F][8:0]};
        compressMaskVecPipe_0 = _RANDOM[6'h1F][9];
        compressMaskVecPipe_1 = _RANDOM[6'h1F][10];
        compressMaskVecPipe_2 = _RANDOM[6'h1F][11];
        compressMaskVecPipe_3 = _RANDOM[6'h1F][12];
        compressMaskVecPipe_4 = _RANDOM[6'h1F][13];
        compressMaskVecPipe_5 = _RANDOM[6'h1F][14];
        compressMaskVecPipe_6 = _RANDOM[6'h1F][15];
        compressMaskVecPipe_7 = _RANDOM[6'h1F][16];
        compressMaskVecPipe_8 = _RANDOM[6'h1F][17];
        compressMaskVecPipe_9 = _RANDOM[6'h1F][18];
        compressMaskVecPipe_10 = _RANDOM[6'h1F][19];
        compressMaskVecPipe_11 = _RANDOM[6'h1F][20];
        compressMaskVecPipe_12 = _RANDOM[6'h1F][21];
        compressMaskVecPipe_13 = _RANDOM[6'h1F][22];
        compressMaskVecPipe_14 = _RANDOM[6'h1F][23];
        compressMaskVecPipe_15 = _RANDOM[6'h1F][24];
        compressMaskVecPipe_16 = _RANDOM[6'h1F][25];
        compressMaskVecPipe_17 = _RANDOM[6'h1F][26];
        compressMaskVecPipe_18 = _RANDOM[6'h1F][27];
        compressMaskVecPipe_19 = _RANDOM[6'h1F][28];
        compressMaskVecPipe_20 = _RANDOM[6'h1F][29];
        compressMaskVecPipe_21 = _RANDOM[6'h1F][30];
        compressMaskVecPipe_22 = _RANDOM[6'h1F][31];
        compressMaskVecPipe_23 = _RANDOM[6'h20][0];
        compressMaskVecPipe_24 = _RANDOM[6'h20][1];
        compressMaskVecPipe_25 = _RANDOM[6'h20][2];
        compressMaskVecPipe_26 = _RANDOM[6'h20][3];
        compressMaskVecPipe_27 = _RANDOM[6'h20][4];
        compressMaskVecPipe_28 = _RANDOM[6'h20][5];
        compressMaskVecPipe_29 = _RANDOM[6'h20][6];
        compressMaskVecPipe_30 = _RANDOM[6'h20][7];
        compressMaskVecPipe_31 = _RANDOM[6'h20][8];
        maskPipe = {_RANDOM[6'h20][31:9], _RANDOM[6'h21][8:0]};
        source2Pipe = {_RANDOM[6'h21][31:9], _RANDOM[6'h22], _RANDOM[6'h23], _RANDOM[6'h24], _RANDOM[6'h25], _RANDOM[6'h26], _RANDOM[6'h27], _RANDOM[6'h28], _RANDOM[6'h29][8:0]};
        lastCompressPipe = _RANDOM[6'h29][9];
        stage2Valid = _RANDOM[6'h29][10];
        newInstructionPipe = _RANDOM[6'h29][11];
        compressInitPipe = _RANDOM[6'h29][21:12];
        compressDeqValidPipe = _RANDOM[6'h29][22];
        groupCounterPipe = _RANDOM[6'h29][28:23];
        compressDataReg = {_RANDOM[6'h29][31:29], _RANDOM[6'h2A], _RANDOM[6'h2B], _RANDOM[6'h2C], _RANDOM[6'h2D], _RANDOM[6'h2E], _RANDOM[6'h2F], _RANDOM[6'h30], _RANDOM[6'h31][28:0]};
        compressTailValid = _RANDOM[6'h31][29];
        compressWriteGroupCount = {_RANDOM[6'h31][31:30], _RANDOM[6'h32][3:0]};
        validInputPipe = _RANDOM[6'h32][11:4];
        readFromScalarPipe = {_RANDOM[6'h32][31:12], _RANDOM[6'h33][11:0]};
        ffoOutPipe = _RANDOM[6'h33][19:12];
        view__out_REG_data = {_RANDOM[6'h33][31:20], _RANDOM[6'h34], _RANDOM[6'h35], _RANDOM[6'h36], _RANDOM[6'h37], _RANDOM[6'h38], _RANDOM[6'h39], _RANDOM[6'h3A], _RANDOM[6'h3B][19:0]};
        view__out_REG_mask = {_RANDOM[6'h3B][31:20], _RANDOM[6'h3C][19:0]};
        view__out_REG_groupCounter = _RANDOM[6'h3C][25:20];
        view__out_REG_ffoOutput = {_RANDOM[6'h3C][31:26], _RANDOM[6'h3D][1:0]};
        view__out_REG_compressValid = _RANDOM[6'h3D][2];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign out_data = view__out_REG_data;
  assign out_mask = view__out_REG_mask;
  assign out_groupCounter = view__out_REG_groupCounter;
  assign out_ffoOutput = view__out_REG_ffoOutput;
  assign out_compressValid = view__out_REG_compressValid;
  assign writeData = ffoIndex;
  assign stageValid = stage2Valid | in_1_valid | compressTailValid;
endmodule

